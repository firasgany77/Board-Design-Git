-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 1 2022 18:02:02

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : in std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : in std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \PCH_PWRGD.count_rst_3\ : std_logic;
signal \PCH_PWRGD.count_rst_10\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.count_rst_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \RSMRST_PWRGD.count_rst_9\ : std_logic;
signal \RSMRST_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_3\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_4_4\ : std_logic;
signal \RSMRST_PWRGD.count_4_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_4_8\ : std_logic;
signal \RSMRST_PWRGD.count_rst_2_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_2\ : std_logic;
signal \RSMRST_PWRGD.count_rst_13\ : std_logic;
signal \RSMRST_PWRGD.count_4_6\ : std_logic;
signal \RSMRST_PWRGD.count_rst_6\ : std_logic;
signal \RSMRST_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_4_1\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_12\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_11_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_RNI166B31Z0Z_12_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_4_0\ : std_logic;
signal \RSMRST_PWRGD.count_4_14\ : std_logic;
signal \RSMRST_PWRGD.count_4_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_5\ : std_logic;
signal \RSMRST_PWRGD.count_4_11\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.count_clkZ0Z_5_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.count_clkZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.count_clk_1_13\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.count_clk_1_11\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.count_clk_1_12\ : std_logic;
signal \POWERLED.count_clk_0_12\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_off_1_13\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_off_1_5\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_1_14\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNINZ0Z4153\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.count_rst_14\ : std_logic;
signal \PCH_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_0\ : std_logic;
signal \PCH_PWRGD.count_rst_8\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_7\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_4\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_5_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_0\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_13_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_9\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.count_rst_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_5_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_8_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_6\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.count_i_0\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \RSMRST_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_14\ : std_logic;
signal \RSMRST_PWRGD.count_4_9\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_1\ : std_logic;
signal \RSMRST_PWRGD.count_rst_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_4_10\ : std_logic;
signal \RSMRST_PWRGD.count_4_13\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \RSMRST_PWRGD.count_rst_7\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_4\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_5\ : std_logic;
signal \RSMRST_PWRGD.count_rst_10\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.count_rst_11\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_9\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.count_rst_0\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.count_rst_3\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_12\ : std_logic;
signal \RSMRST_PWRGD.count_rst_4\ : std_logic;
signal \RSMRST_PWRGD.count_4_15\ : std_logic;
signal \RSMRST_PWRGD.N_240_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.count_4_12\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_1\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.N_178\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.count_clk_1_14\ : std_logic;
signal \POWERLED.count_clk_0_14\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_ns_1_1_0\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_1_0\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal \POWERLED.count_clkZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\ : std_logic;
signal \POWERLED.N_193\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.N_385\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.N_385_cascade_\ : std_logic;
signal \POWERLED.count_clk_en_0_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_4_i_a2_1\ : std_logic;
signal \POWERLED.count_clk_en_2_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_10\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.count_off_1_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI_3Z0Z_0\ : std_logic;
signal \POWERLED.func_state_RNI_3Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_1\ : std_logic;
signal \POWERLED.N_321_cascade_\ : std_logic;
signal \POWERLED.N_431\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_336_N\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_1\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_off_1_1_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.un34_clk_100khz_10\ : std_logic;
signal \POWERLED.un34_clk_100khz_8\ : std_logic;
signal \POWERLED.un34_clk_100khz_9_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.N_128\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \POWERLED.count_off_0_9\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_11\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_off_1_10\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.count_off_0_11\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \POWERLED.count_off_1_12\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \PCH_PWRGD.curr_state_7_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_1_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2857_i_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \PCH_PWRGD.curr_state_7_1_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa_cascade_\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.count_rst_7\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.count_rst_11\ : std_logic;
signal \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_3\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_0_1\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_0_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.N_277_0\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI1IPC1Z0Z_0\ : std_logic;
signal \PCH_PWRGD.N_277_0_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \PCH_PWRGD.N_2857_i\ : std_logic;
signal \PCH_PWRGD.N_413\ : std_logic;
signal \PCH_PWRGD.N_413_cascade_\ : std_logic;
signal \PCH_PWRGD.N_424\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_2859_i\ : std_logic;
signal \PCH_PWRGD.N_278_0\ : std_logic;
signal \RSMRST_PWRGD.count_rst_8\ : std_logic;
signal \RSMRST_PWRGD.count_4_3\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal \POWERLED.count_1_0_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_1_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_0_1\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \curr_state_RNIR5QD1_0_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_state_2_0\ : std_logic;
signal \RSMRST_PWRGD.m4_0_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_state_7_1\ : std_logic;
signal \RSMRST_PWRGD.count_RNI166B31Z0Z_12\ : std_logic;
signal \RSMRST_PWRGD.curr_state_1_1\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal \POWERLED.count_0_2\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.count_0_12\ : std_logic;
signal \POWERLED.curr_state_0_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.count_off_0_2\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_off_0_3\ : std_logic;
signal \POWERLED.count_off_1_3\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.count_off_1_4\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal vccst_en : std_logic;
signal \POWERLED.N_359_cascade_\ : std_logic;
signal \POWERLED.N_171_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_oZ0Z3\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_0_o3_out_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI3IN21Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_ns_1_1_1_cascade_\ : std_logic;
signal \POWERLED.N_2905_i_cascade_\ : std_logic;
signal \POWERLED.N_175_cascade_\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_a2Z0Z_3\ : std_logic;
signal \POWERLED.func_state_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI_4Z0Z_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_a2_1\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.N_301\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_\ : std_logic;
signal \POWERLED.N_238_cascade_\ : std_logic;
signal \POWERLED.N_118_f0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIS3763Z0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \POWERLED.N_171\ : std_logic;
signal \POWERLED.dutycycle_RNIS3763Z0Z_2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_2\ : std_logic;
signal \POWERLED.dutycycle_cascade_\ : std_logic;
signal \POWERLED.N_5_1\ : std_logic;
signal \POWERLED.g0_i_a6_0_1_cascade_\ : std_logic;
signal \POWERLED.g2_1_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_5_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_5_0_N_3_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.g0_i_1\ : std_logic;
signal \POWERLED.dutycycle_en_5_0_0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.count_off_0_6\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.count_off_0_7\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.count_off_1_8\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \HDA_STRAP.curr_state_2_1\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal \HDA_STRAP.curr_state_i_2_cascade_\ : std_logic;
signal \HDA_STRAP.i4_mux\ : std_logic;
signal \HDA_STRAP.N_208\ : std_logic;
signal \HDA_STRAP.curr_state_i_2\ : std_logic;
signal \HDA_STRAP.N_208_cascade_\ : std_logic;
signal \HDA_STRAP.HDA_SDO_ATP_0\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \POWERLED.func_state_enZ0\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \VPP_VDDQ.N_2897_i_cascade_\ : std_logic;
signal \POWERLED.count_0_4\ : std_logic;
signal \RSMRST_PWRGD.N_423\ : std_logic;
signal \RSMRST_PWRGD.count_0_sqmuxa\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \POWERLED.count_0_5\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \POWERLED.count_1_2\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.count_1_3\ : std_logic;
signal \POWERLED.un1_count_cry_2\ : std_logic;
signal \POWERLED.count_1_4\ : std_logic;
signal \POWERLED.un1_count_cry_3\ : std_logic;
signal \POWERLED.count_1_5\ : std_logic;
signal \POWERLED.un1_count_cry_4\ : std_logic;
signal \POWERLED.count_1_6\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \POWERLED.count_1_10\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.count_1_11\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.count_1_12\ : std_logic;
signal \POWERLED.un1_count_cry_11\ : std_logic;
signal \POWERLED.count_1_13\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.un1_count_cry_13\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.count_1_14\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.N_8_2_cascade_\ : std_logic;
signal \POWERLED.N_5_0_cascade_\ : std_logic;
signal \POWERLED.g0_5_0\ : std_logic;
signal \POWERLED.N_331_N_0_0_cascade_\ : std_logic;
signal \POWERLED.g3_1_0_1\ : std_logic;
signal \POWERLED.g3_1_0\ : std_logic;
signal \POWERLED.func_m1_0_a2Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o2_1\ : std_logic;
signal \POWERLED.N_433_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_ns_1_1\ : std_logic;
signal \POWERLED.func_state_1_m2_1\ : std_logic;
signal \POWERLED.N_345\ : std_logic;
signal \POWERLED.N_164\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_0\ : std_logic;
signal \POWERLED.N_344_cascade_\ : std_logic;
signal \POWERLED.N_343\ : std_logic;
signal \POWERLED.N_79\ : std_logic;
signal \POWERLED.func_state_RNI3IN21Z0Z_0\ : std_logic;
signal \POWERLED.N_433\ : std_logic;
signal \POWERLED.N_79_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_ns_1_0\ : std_logic;
signal \POWERLED.func_state_1_m2_0\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_2\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_a3_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIH0LB7Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \POWERLED.N_189_i\ : std_logic;
signal \POWERLED.N_189_i_cascade_\ : std_logic;
signal \POWERLED.N_122_f0_1_cascade_\ : std_logic;
signal \POWERLED.N_122_f0_1\ : std_logic;
signal \POWERLED.g0_i_a6_1_1_cascade_\ : std_logic;
signal \POWERLED.N_10_0\ : std_logic;
signal \tmp_1_rep1_RNI_cascade_\ : std_logic;
signal \POWERLED.N_358_cascade_\ : std_logic;
signal \POWERLED.N_12\ : std_logic;
signal \POWERLED.g0_i_a6_1\ : std_logic;
signal \POWERLED.N_358\ : std_logic;
signal \POWERLED.un1_clk_100khz_42_and_i_a2_3_0_cascade_\ : std_logic;
signal \POWERLED.N_434_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_0\ : std_logic;
signal \POWERLED.N_372_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_0\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_1\ : std_logic;
signal \POWERLED.dutycycle_eena_0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_1\ : std_logic;
signal \POWERLED.dutycycle_1_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_7\ : std_logic;
signal \POWERLED.dutycycleZ1Z_11\ : std_logic;
signal \POWERLED.dutycycle_eena_7_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_12_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_2\ : std_logic;
signal \N_414_cascade_\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.m6_i_0\ : std_logic;
signal \HDA_STRAP.m6_i_0_cascade_\ : std_logic;
signal \HDA_STRAP.curr_state_3_0\ : std_logic;
signal \HDA_STRAP.N_53_cascade_\ : std_logic;
signal \HDA_STRAP.N_285\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.N_285_cascade_\ : std_logic;
signal \HDA_STRAP.N_51\ : std_logic;
signal vccst_pwrgd : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0\ : std_logic;
signal \N_227\ : std_logic;
signal \N_227_cascade_\ : std_logic;
signal pch_pwrok : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \DSW_PWRGD.un4_count_11_cascade_\ : std_logic;
signal \DSW_PWRGD.un4_count_10\ : std_logic;
signal \DSW_PWRGD.un4_count_8\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER.un4_counter_7\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_0\ : std_logic;
signal vddq_ok : std_logic;
signal \VPP_VDDQ.N_2897_i\ : std_logic;
signal \VPP_VDDQ.N_297_0\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlt6_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_3\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \POWERLED.count_1_7\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.count_1_8\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \POWERLED.count_1_9\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.g0_8_sx\ : std_logic;
signal \SUSWARN_N_rep1\ : std_logic;
signal \N_414\ : std_logic;
signal \HDA_STRAP.count_enZ0\ : std_logic;
signal \COUNTER.un4_counter_7_THRU_CO\ : std_logic;
signal v1p8a_en : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRSTn_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.N_2989_i\ : std_logic;
signal \POWERLED_un1_clk_100khz_52_and_i_0\ : std_logic;
signal \COUNTER.N_96_mux_i_i_a8_1_cascade_\ : std_logic;
signal \tmp_1_rep1_RNIC08FV_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNII69M3Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_6_cascade_\ : std_logic;
signal \N_96_mux_i_i_3\ : std_logic;
signal \N_96_mux_i_i_3_cascade_\ : std_logic;
signal \COUNTER.N_96_mux_i_i_a8_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5\ : std_logic;
signal \POWERLED.N_31\ : std_logic;
signal \POWERLED.N_31_cascade_\ : std_logic;
signal \POWERLED.g0_i_a6_0\ : std_logic;
signal \POWERLED.N_237\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_0_1_1\ : std_logic;
signal \POWERLED.N_387_cascade_\ : std_logic;
signal slp_s3n : std_logic;
signal slp_s4n : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.N_372\ : std_logic;
signal \POWERLED.func_state_RNIDUQ02Z0Z_1\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_m2_0_1_cascade_\ : std_logic;
signal \POWERLED.N_233_N_cascade_\ : std_logic;
signal \POWERLED.N_311\ : std_logic;
signal \POWERLED.dutycycle_eena_13_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7TZ0Z3\ : std_logic;
signal \POWERLED.dutycycle_eena_13\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.N_388\ : std_logic;
signal \POWERLED_dutycycle_set_1\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\ : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_337_N\ : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3\ : std_logic;
signal \POWERLED.N_308\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_cZ0\ : std_logic;
signal \POWERLED.N_307\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \bfn_6_16_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9\ : std_logic;
signal \POWERLED.dutycycle_rst_6\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12\ : std_logic;
signal \POWERLED.N_175_i\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \VPP_VDDQ.count_3_2\ : std_logic;
signal \VPP_VDDQ.count_3_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6_cascade_\ : std_logic;
signal \VPP_VDDQ.count_3_10\ : std_logic;
signal \VPP_VDDQ.count_rst_5_cascade_\ : std_logic;
signal \VPP_VDDQ.N_3013_i_cascade_\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_8\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_RNI_1_10_cascade_\ : std_logic;
signal \VPP_VDDQ.count_3_11\ : std_logic;
signal \VPP_VDDQ.N_3013_i\ : std_logic;
signal \VPP_VDDQ.count_3_0\ : std_logic;
signal \VPP_VDDQ.count_en_cascade_\ : std_logic;
signal \VPP_VDDQ.count_3_1\ : std_logic;
signal \VPP_VDDQ.count_3_9\ : std_logic;
signal \VPP_VDDQ.count_3_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_11\ : std_logic;
signal \DSW_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_1\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_2\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \DSW_PWRGD.countZ0Z_3\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \DSW_PWRGD.countZ0Z_4\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \DSW_PWRGD.countZ0Z_5\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \DSW_PWRGD.countZ0Z_6\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \DSW_PWRGD.countZ0Z_7\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \DSW_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_9\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \DSW_PWRGD.countZ0Z_10\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \DSW_PWRGD.countZ0Z_11\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.m4_0_a2\ : std_logic;
signal \VPP_VDDQ.m4_0_cascade_\ : std_logic;
signal suswarn_n : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_2877_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\ : std_logic;
signal \VPP_VDDQ.N_2877_i_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \VPP_VDDQ.count_3_15\ : std_logic;
signal \POWERLED.N_203_i_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI0TA81_0Z0Z_0\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.g0_13_sx\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_a2_1_sx_cascade_\ : std_logic;
signal rsmrstn : std_logic;
signal \curr_state_RNIR5QD1_0_0\ : std_logic;
signal \POWERLED.g0_1\ : std_logic;
signal \SUSWARN_N_fast\ : std_logic;
signal \RSMRST_PWRGD_RSMRSTn_fast\ : std_logic;
signal \POWERLED.g1_2_0\ : std_logic;
signal \POWERLED.func_state_RNI3IN21_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI3IN21Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6\ : std_logic;
signal \POWERLED.N_312\ : std_logic;
signal \POWERLED.func_state\ : std_logic;
signal \POWERLED.N_389\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\ : std_logic;
signal \POWERLED.dutycycle_RNI554R1Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI778D2Z0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI778D2Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIKGV14Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIKGV14Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI554R1Z0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \POWERLED.N_332_N\ : std_logic;
signal \POWERLED.N_116_f0\ : std_logic;
signal \POWERLED.N_116_f0_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\ : std_logic;
signal \POWERLED.dutycycle_e_1_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.N_157_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\ : std_logic;
signal \POWERLED.dutycycle_en_4_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_10\ : std_logic;
signal \VPP_VDDQ.count_3_3\ : std_logic;
signal \VPP_VDDQ.count_3_4\ : std_logic;
signal \VPP_VDDQ.count_3_5\ : std_logic;
signal \VPP_VDDQ.un4_count_1_axb_0\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_rst_6\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.count_rst_7\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.count_rst_8\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_2_cZ0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.count_rst_9\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_3_cZ0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.count_rst_10\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_4_cZ0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.count_rst_11\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_6_cZ0\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_7_cZ0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.count_rst_13\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \VPP_VDDQ.count_RNI_1_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.count_rst_14\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_8_cZ0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.count_rst\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6CZ0\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_13\ : std_logic;
signal \DSW_PWRGD.countZ0Z_15\ : std_logic;
signal \DSW_PWRGD.countZ0Z_14\ : std_logic;
signal \DSW_PWRGD.countZ0Z_12\ : std_logic;
signal \DSW_PWRGD.un4_count_9\ : std_logic;
signal v33a_ok : std_logic;
signal v5a_ok : std_logic;
signal v1p8a_ok : std_logic;
signal slp_susn : std_logic;
signal \DSW_PWRGD.i3_mux_0_cascade_\ : std_logic;
signal \DSW_PWRGD.N_1_i\ : std_logic;
signal \DSW_PWRGD.N_6_cascade_\ : std_logic;
signal \DSW_PWRGD.un1_curr_state10_0\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2_c\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_c\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_c\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_c\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_c\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \DSW_PWRGD.N_22_0\ : std_logic;
signal \POWERLED.func_state_RNI1E8A4_0_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal \POWERLED.count_clk_en\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2898\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8\ : std_logic;
signal \POWERLED.curr_state_3_0\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_0\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.un1_count_cry_0_i\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.un85_clk_100khz_1\ : std_logic;
signal \POWERLED.N_6108_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.N_6109_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.un85_clk_100khz_3\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.N_6110_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.un85_clk_100khz_4\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.N_6111_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_8\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.N_6112_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_8\ : std_logic;
signal \POWERLED.N_6113_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_8\ : std_logic;
signal \POWERLED.N_6114_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.N_6115_i\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_8\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.N_6116_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_8\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.N_6117_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.N_6118_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.N_6119_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.N_6120_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.N_6121_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_6122_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_8\ : std_logic;
signal \POWERLED.N_96_mux_i_i_2_1\ : std_logic;
signal \N_96_mux_i_i_2\ : std_logic;
signal \N_13\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_8\ : std_logic;
signal \POWERLED.count_off_1_sqmuxa\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m4\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1\ : std_logic;
signal \POWERLED.N_2905_i\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\ : std_logic;
signal \POWERLED.N_19\ : std_logic;
signal \POWERLED.N_134_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m0\ : std_logic;
signal \POWERLED.g2_0_1_0\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m0_cascade_\ : std_logic;
signal \POWERLED.N_15\ : std_logic;
signal \POWERLED.N_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_6\ : std_logic;
signal \tmp_1_rep1_RNI\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_0\ : std_logic;
signal \POWERLED.N_361_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_9Z0Z_3\ : std_logic;
signal \POWERLED.N_361\ : std_logic;
signal \POWERLED.N_369\ : std_logic;
signal \POWERLED.d_i3_mux\ : std_logic;
signal \POWERLED.un1_i3_mux_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\ : std_logic;
signal \POWERLED.dutycycleZ1Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNIQU4T5Z0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_11\ : std_logic;
signal \POWERLED.N_156_N_cascade_\ : std_logic;
signal \POWERLED.N_158_N\ : std_logic;
signal \POWERLED.func_state_RNIHU7V2Z0Z_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.N_161_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_12\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\ : std_logic;
signal \POWERLED.dutycycle_en_12_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \VPP_VDDQ.count_rst_1\ : std_logic;
signal \VPP_VDDQ.count_3_12\ : std_logic;
signal \VPP_VDDQ.count_rst_12\ : std_logic;
signal \VPP_VDDQ.count_3_7\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \VPP_VDDQ.count_2_0_6\ : std_logic;
signal \VPP_VDDQ.count_3_13\ : std_logic;
signal \VPP_VDDQ.count_rst_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.count_en\ : std_logic;
signal \VPP_VDDQ.count_3_14\ : std_logic;
signal \VPP_VDDQ.count_rst_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_0_cascade_\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_2\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_3\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal v33dsw_ok : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \DSW_PWRGD.curr_state10\ : std_logic;
signal vccst_cpu_ok : std_logic;
signal v5s_ok : std_logic;
signal v33s_ok : std_logic;
signal dsw_pwrok : std_logic;
signal \N_392\ : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\ : std_logic;
signal v5s_enn : std_logic;
signal vccin_en : std_logic;
signal \DSW_PWRGD_un1_curr_state_0_sqmuxa_0\ : std_logic;
signal \un4_counter_7_c_RNIBJDJ\ : std_logic;
signal \un4_counter_7_c_RNI09TK5\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_2\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.g0_i_o3_0\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.N_8\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_5_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_4_7\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\ : std_logic;
signal \RSMRST_PWRGD.count_rst_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \POWERLED.mult1_un145_sum\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_2\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_2\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_7\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_8\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.N_428\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_13_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \POWERLED.dutycycle_en_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.g0_4_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_25_1_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_7_cascade_\ : std_logic;
signal \tmp_1_rep1_RNIC08FV_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_9\ : std_logic;
signal \POWERLED.func_m1_0_a2Z0Z_0\ : std_logic;
signal \POWERLED.N_235_N\ : std_logic;
signal \POWERLED.dutycycle_eena_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.dutycycle_eena_9_cascade_\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_pwrgd_en\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_12_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_14_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \VPP_VDDQ.count_2_rst_6\ : std_logic;
signal \VPP_VDDQ.count_2_rst_6_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.count_2_rst_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.count_2_rst_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.count_2_rst_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_10\ : std_logic;
signal \VPP_VDDQ.count_2_rst_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_12\ : std_logic;
signal \VPP_VDDQ.count_2_rst_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_14\ : std_logic;
signal \VPP_VDDQ.count_2_rst_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.count_2_rst_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \HDA_STRAP.count_1_0_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_0_cascade_\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_13_cascade_\ : std_logic;
signal \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_\ : std_logic;
signal \HDA_STRAP.count_1_0_0\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_7\ : std_logic;
signal \HDA_STRAP.count_1_0_8\ : std_logic;
signal \HDA_STRAP.count_1_0_6\ : std_logic;
signal \HDA_STRAP.count_1_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_6_cascade_\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_6\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_0\ : std_logic;
signal \HDA_STRAP.count_1_12\ : std_logic;
signal \HDA_STRAP.count_1_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_12_cascade_\ : std_logic;
signal \HDA_STRAP.count_1_5\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_2\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_3_cascade_\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_4\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_14\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_5\ : std_logic;
signal \HDA_STRAP.count_1_13\ : std_logic;
signal \HDA_STRAP.count_1_3\ : std_logic;
signal \VCCST_EN_i_0_o3_0\ : std_logic;
signal vpp_en : std_logic;
signal \VPP_VDDQ.N_194\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_pwrgd_en_g\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8_cascade_\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_4_sf\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \POWERLED.un1_clk_100khz_43_and_i_0_d_0\ : std_logic;
signal \POWERLED.m21_e_1_cascade_\ : std_logic;
signal \POWERLED.N_5\ : std_logic;
signal \POWERLED.mult1_un47_sum\ : std_logic;
signal \POWERLED.mult1_un47_sum_i\ : std_logic;
signal \POWERLED.g2_0_0_0\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_6\ : std_logic;
signal \POWERLED.g2_0_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_a1_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_8\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_11\ : std_logic;
signal \POWERLED.g0_0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_a3_0\ : std_logic;
signal \POWERLED.N_371\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.g2\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_11\ : std_logic;
signal \POWERLED.g0_1_0\ : std_logic;
signal \POWERLED.func_state_RNI_6Z0Z_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_40_and_i_0_d_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.func_m1_0_a2_0_isoZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_14_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_1_4\ : std_logic;
signal \POWERLED.dutycycle_en_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_13\ : std_logic;
signal \POWERLED.func_state_RNI3IN21_0Z0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_1_0_tz\ : std_logic;
signal \POWERLED.un1_dutycycle_53_3_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.count_2_rst_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_4\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_12\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_5_cascade_\ : std_logic;
signal \VPP_VDDQ.N_1_i_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_rst_3\ : std_logic;
signal \VPP_VDDQ.count_2_rst_3_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_11\ : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.count_2_rst_8_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_rst_7_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.count_2_0_sqmuxa\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2_0_4\ : std_logic;
signal \VPP_VDDQ.count_2_rst_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_2_cascade_\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_1\ : std_logic;
signal \HDA_STRAP.count_RNIZ0Z_1\ : std_logic;
signal \HDA_STRAP.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_1_cascade_\ : std_logic;
signal \HDA_STRAP.count_1_1\ : std_logic;
signal \HDA_STRAP.count_1_2\ : std_logic;
signal \HDA_STRAP.count_1_0_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_1\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_3\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_5\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.count_1_6\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_5_cZ0\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_8\ : std_logic;
signal \HDA_STRAP.count_1_8\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_7\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_9\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.count_1_11\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_13\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_15\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_16\ : std_logic;
signal \HDA_STRAP.count_1_16\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_15\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_16\ : std_logic;
signal \HDA_STRAP.count_RNI6OA47Z0Z_8\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\ : std_logic;
signal \HDA_STRAP.count_0_17\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\ : std_logic;
signal \HDA_STRAP.count_1_4\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\ : std_logic;
signal \HDA_STRAP.count_1_7\ : std_logic;
signal \HDA_STRAP.count_1_10\ : std_logic;
signal \HDA_STRAP.count_1_0_10\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3\ : std_logic;
signal \HDA_STRAP.count_1_14\ : std_logic;
signal fpga_osc : std_logic;
signal \HDA_STRAP.count_en_g\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.g0_7_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.g3_1_3_0_cascade_\ : std_logic;
signal \POWERLED.g0_10_0_0_0\ : std_logic;
signal \POWERLED.N_3034_0_0_0\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \POWERLED.N_203_i\ : std_logic;
signal \POWERLED.g0_10_0_0_1\ : std_logic;
signal \POWERLED.N_175\ : std_logic;
signal \POWERLED.g3_1_3_0\ : std_logic;
signal \POWERLED.N_3034_0_0_2\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_4_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_10_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_a0_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_a1_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_5_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_31_a7_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_a0_1\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_6\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_39_c_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_49_0_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_49_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_39_c_1_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_53_34_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_36_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_34_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_12\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    \VCCINAUX_VR_PE_wire\ <= VCCINAUX_VR_PE;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    \VCCIN_VR_PE_wire\ <= VCCIN_VR_PE;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38057\,
            DIN => \N__38056\,
            DOUT => \N__38055\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38057\,
            PADOUT => \N__38056\,
            PADIN => \N__38055\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38048\,
            DIN => \N__38047\,
            DOUT => \N__38046\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38048\,
            PADOUT => \N__38047\,
            PADIN => \N__38046\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38039\,
            DIN => \N__38038\,
            DOUT => \N__38037\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38039\,
            PADOUT => \N__38038\,
            PADIN => \N__38037\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21973\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38030\,
            DIN => \N__38029\,
            DOUT => \N__38028\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38030\,
            PADOUT => \N__38029\,
            PADIN => \N__38028\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19084\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38021\,
            DIN => \N__38020\,
            DOUT => \N__38019\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38021\,
            PADOUT => \N__38020\,
            PADIN => \N__38019\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38012\,
            DIN => \N__38011\,
            DOUT => \N__38010\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38012\,
            PADOUT => \N__38011\,
            PADIN => \N__38010\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38003\,
            DIN => \N__38002\,
            DOUT => \N__38001\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38003\,
            PADOUT => \N__38002\,
            PADIN => \N__38001\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37994\,
            DIN => \N__37993\,
            DOUT => \N__37992\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37994\,
            PADOUT => \N__37993\,
            PADIN => \N__37992\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37985\,
            DIN => \N__37984\,
            DOUT => \N__37983\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37985\,
            PADOUT => \N__37984\,
            PADIN => \N__37983\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27989\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__37976\,
            DIN => \N__37975\,
            DOUT => \N__37974\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37976\,
            PADOUT => \N__37975\,
            PADIN => \N__37974\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37967\,
            DIN => \N__37966\,
            DOUT => \N__37965\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37967\,
            PADOUT => \N__37966\,
            PADIN => \N__37965\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37958\,
            DIN => \N__37957\,
            DOUT => \N__37956\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37958\,
            PADOUT => \N__37957\,
            PADIN => \N__37956\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17143\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37949\,
            DIN => \N__37948\,
            DOUT => \N__37947\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37949\,
            PADOUT => \N__37948\,
            PADIN => \N__37947\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37940\,
            DIN => \N__37939\,
            DOUT => \N__37938\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37940\,
            PADOUT => \N__37939\,
            PADIN => \N__37938\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37931\,
            DIN => \N__37930\,
            DOUT => \N__37929\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37931\,
            PADOUT => \N__37930\,
            PADIN => \N__37929\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37922\,
            DIN => \N__37921\,
            DOUT => \N__37920\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37922\,
            PADOUT => \N__37921\,
            PADIN => \N__37920\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37913\,
            DIN => \N__37912\,
            DOUT => \N__37911\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37913\,
            PADOUT => \N__37912\,
            PADIN => \N__37911\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18793\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__37904\,
            DIN => \N__37903\,
            DOUT => \N__37902\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37904\,
            PADOUT => \N__37903\,
            PADIN => \N__37902\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37895\,
            DIN => \N__37894\,
            DOUT => \N__37893\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37895\,
            PADOUT => \N__37894\,
            PADIN => \N__37893\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37886\,
            DIN => \N__37885\,
            DOUT => \N__37884\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37886\,
            PADOUT => \N__37885\,
            PADIN => \N__37884\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23746\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37877\,
            DIN => \N__37876\,
            DOUT => \N__37875\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37877\,
            PADOUT => \N__37876\,
            PADIN => \N__37875\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37868\,
            DIN => \N__37867\,
            DOUT => \N__37866\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37868\,
            PADOUT => \N__37867\,
            PADIN => \N__37866\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37859\,
            DIN => \N__37858\,
            DOUT => \N__37857\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37859\,
            PADOUT => \N__37858\,
            PADIN => \N__37857\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__37850\,
            DIN => \N__37849\,
            DOUT => \N__37848\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37850\,
            PADOUT => \N__37849\,
            PADIN => \N__37848\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37841\,
            DIN => \N__37840\,
            DOUT => \N__37839\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37841\,
            PADOUT => \N__37840\,
            PADIN => \N__37839\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24331\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37832\,
            DIN => \N__37831\,
            DOUT => \N__37830\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37832\,
            PADOUT => \N__37831\,
            PADIN => \N__37830\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37823\,
            DIN => \N__37822\,
            DOUT => \N__37821\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37823\,
            PADOUT => \N__37822\,
            PADIN => \N__37821\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21142\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37814\,
            DIN => \N__37813\,
            DOUT => \N__37812\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37814\,
            PADOUT => \N__37813\,
            PADIN => \N__37812\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21091\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37805\,
            DIN => \N__37804\,
            DOUT => \N__37803\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37805\,
            PADOUT => \N__37804\,
            PADIN => \N__37803\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37796\,
            DIN => \N__37795\,
            DOUT => \N__37794\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37796\,
            PADOUT => \N__37795\,
            PADIN => \N__37794\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37787\,
            DIN => \N__37786\,
            DOUT => \N__37785\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37787\,
            PADOUT => \N__37786\,
            PADIN => \N__37785\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37778\,
            DIN => \N__37777\,
            DOUT => \N__37776\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37778\,
            PADOUT => \N__37777\,
            PADIN => \N__37776\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37769\,
            DIN => \N__37768\,
            DOUT => \N__37767\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37769\,
            PADOUT => \N__37768\,
            PADIN => \N__37767\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37760\,
            DIN => \N__37759\,
            DOUT => \N__37758\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37760\,
            PADOUT => \N__37759\,
            PADIN => \N__37758\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19483\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37751\,
            DIN => \N__37750\,
            DOUT => \N__37749\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37751\,
            PADOUT => \N__37750\,
            PADIN => \N__37749\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37742\,
            DIN => \N__37741\,
            DOUT => \N__37740\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37742\,
            PADOUT => \N__37741\,
            PADIN => \N__37740\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31093\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__37733\,
            DIN => \N__37732\,
            DOUT => \N__37731\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37733\,
            PADOUT => \N__37732\,
            PADIN => \N__37731\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37724\,
            DIN => \N__37723\,
            DOUT => \N__37722\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37724\,
            PADOUT => \N__37723\,
            PADIN => \N__37722\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37715\,
            DIN => \N__37714\,
            DOUT => \N__37713\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37715\,
            PADOUT => \N__37714\,
            PADIN => \N__37713\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37706\,
            DIN => \N__37705\,
            DOUT => \N__37704\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37706\,
            PADOUT => \N__37705\,
            PADIN => \N__37704\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37697\,
            DIN => \N__37696\,
            DOUT => \N__37695\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37697\,
            PADOUT => \N__37696\,
            PADIN => \N__37695\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25194\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37688\,
            DIN => \N__37687\,
            DOUT => \N__37686\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37688\,
            PADOUT => \N__37687\,
            PADIN => \N__37686\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37679\,
            DIN => \N__37678\,
            DOUT => \N__37677\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37679\,
            PADOUT => \N__37678\,
            PADIN => \N__37677\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27990\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37670\,
            DIN => \N__37669\,
            DOUT => \N__37668\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37670\,
            PADOUT => \N__37669\,
            PADIN => \N__37668\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37661\,
            DIN => \N__37660\,
            DOUT => \N__37659\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37661\,
            PADOUT => \N__37660\,
            PADIN => \N__37659\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28081\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37652\,
            DIN => \N__37651\,
            DOUT => \N__37650\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37652\,
            PADOUT => \N__37651\,
            PADIN => \N__37650\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25249\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37643\,
            DIN => \N__37642\,
            DOUT => \N__37641\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37643\,
            PADOUT => \N__37642\,
            PADIN => \N__37641\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37634\,
            DIN => \N__37633\,
            DOUT => \N__37632\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37634\,
            PADOUT => \N__37633\,
            PADIN => \N__37632\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__37625\,
            DIN => \N__37624\,
            DOUT => \N__37623\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37625\,
            PADOUT => \N__37624\,
            PADIN => \N__37623\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37616\,
            DIN => \N__37615\,
            DOUT => \N__37614\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37616\,
            PADOUT => \N__37615\,
            PADIN => \N__37614\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37607\,
            DIN => \N__37606\,
            DOUT => \N__37605\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37607\,
            PADOUT => \N__37606\,
            PADIN => \N__37605\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27868\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37598\,
            DIN => \N__37597\,
            DOUT => \N__37596\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37598\,
            PADOUT => \N__37597\,
            PADIN => \N__37596\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37589\,
            DIN => \N__37588\,
            DOUT => \N__37587\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37589\,
            PADOUT => \N__37588\,
            PADIN => \N__37587\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37580\,
            DIN => \N__37579\,
            DOUT => \N__37578\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37580\,
            PADOUT => \N__37579\,
            PADIN => \N__37578\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37571\,
            DIN => \N__37570\,
            DOUT => \N__37569\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37571\,
            PADOUT => \N__37570\,
            PADIN => \N__37569\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37562\,
            DIN => \N__37561\,
            DOUT => \N__37560\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37562\,
            PADOUT => \N__37561\,
            PADIN => \N__37560\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37553\,
            DIN => \N__37552\,
            DOUT => \N__37551\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37553\,
            PADOUT => \N__37552\,
            PADIN => \N__37551\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37544\,
            DIN => \N__37543\,
            DOUT => \N__37542\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37544\,
            PADOUT => \N__37543\,
            PADIN => \N__37542\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21078\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37535\,
            DIN => \N__37534\,
            DOUT => \N__37533\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37535\,
            PADOUT => \N__37534\,
            PADIN => \N__37533\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__8718\ : CascadeMux
    port map (
            O => \N__37516\,
            I => \N__37505\
        );

    \I__8717\ : CascadeMux
    port map (
            O => \N__37515\,
            I => \N__37502\
        );

    \I__8716\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37498\
        );

    \I__8715\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37493\
        );

    \I__8714\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37493\
        );

    \I__8713\ : CascadeMux
    port map (
            O => \N__37511\,
            I => \N__37489\
        );

    \I__8712\ : InMux
    port map (
            O => \N__37510\,
            I => \N__37486\
        );

    \I__8711\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37479\
        );

    \I__8710\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37479\
        );

    \I__8709\ : InMux
    port map (
            O => \N__37505\,
            I => \N__37479\
        );

    \I__8708\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37474\
        );

    \I__8707\ : InMux
    port map (
            O => \N__37501\,
            I => \N__37474\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__37498\,
            I => \N__37471\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__37493\,
            I => \N__37468\
        );

    \I__8704\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37463\
        );

    \I__8703\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37463\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__37486\,
            I => \N__37460\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37457\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__37474\,
            I => \N__37454\
        );

    \I__8699\ : Span4Mux_s0_h
    port map (
            O => \N__37471\,
            I => \N__37447\
        );

    \I__8698\ : Span4Mux_s2_v
    port map (
            O => \N__37468\,
            I => \N__37447\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__37463\,
            I => \N__37447\
        );

    \I__8696\ : Span4Mux_s2_v
    port map (
            O => \N__37460\,
            I => \N__37443\
        );

    \I__8695\ : Span12Mux_s2_v
    port map (
            O => \N__37457\,
            I => \N__37440\
        );

    \I__8694\ : Span4Mux_s2_v
    port map (
            O => \N__37454\,
            I => \N__37435\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__37447\,
            I => \N__37435\
        );

    \I__8692\ : InMux
    port map (
            O => \N__37446\,
            I => \N__37432\
        );

    \I__8691\ : Odrv4
    port map (
            O => \N__37443\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__8690\ : Odrv12
    port map (
            O => \N__37440\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__8689\ : Odrv4
    port map (
            O => \N__37435\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__37432\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__8687\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37420\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__37420\,
            I => \POWERLED.un1_dutycycle_53_39_c_1_0\
        );

    \I__8685\ : CascadeMux
    port map (
            O => \N__37417\,
            I => \N__37409\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__37416\,
            I => \N__37406\
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__37415\,
            I => \N__37402\
        );

    \I__8682\ : InMux
    port map (
            O => \N__37414\,
            I => \N__37389\
        );

    \I__8681\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37389\
        );

    \I__8680\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37389\
        );

    \I__8679\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37382\
        );

    \I__8678\ : InMux
    port map (
            O => \N__37406\,
            I => \N__37382\
        );

    \I__8677\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37382\
        );

    \I__8676\ : InMux
    port map (
            O => \N__37402\,
            I => \N__37377\
        );

    \I__8675\ : InMux
    port map (
            O => \N__37401\,
            I => \N__37377\
        );

    \I__8674\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37370\
        );

    \I__8673\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37370\
        );

    \I__8672\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37370\
        );

    \I__8671\ : CascadeMux
    port map (
            O => \N__37397\,
            I => \N__37366\
        );

    \I__8670\ : CascadeMux
    port map (
            O => \N__37396\,
            I => \N__37362\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__37389\,
            I => \N__37355\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__37382\,
            I => \N__37348\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37348\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__37370\,
            I => \N__37348\
        );

    \I__8665\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37337\
        );

    \I__8664\ : InMux
    port map (
            O => \N__37366\,
            I => \N__37337\
        );

    \I__8663\ : InMux
    port map (
            O => \N__37365\,
            I => \N__37337\
        );

    \I__8662\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37337\
        );

    \I__8661\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37337\
        );

    \I__8660\ : InMux
    port map (
            O => \N__37360\,
            I => \N__37327\
        );

    \I__8659\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37327\
        );

    \I__8658\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37327\
        );

    \I__8657\ : Span4Mux_s0_h
    port map (
            O => \N__37355\,
            I => \N__37320\
        );

    \I__8656\ : Span4Mux_s2_v
    port map (
            O => \N__37348\,
            I => \N__37320\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37320\
        );

    \I__8654\ : InMux
    port map (
            O => \N__37336\,
            I => \N__37317\
        );

    \I__8653\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37314\
        );

    \I__8652\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37311\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__37327\,
            I => \N__37308\
        );

    \I__8650\ : Span4Mux_h
    port map (
            O => \N__37320\,
            I => \N__37305\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__37317\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__37314\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__37311\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__8646\ : Odrv4
    port map (
            O => \N__37308\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__8645\ : Odrv4
    port map (
            O => \N__37305\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__37294\,
            I => \N__37287\
        );

    \I__8643\ : CascadeMux
    port map (
            O => \N__37293\,
            I => \N__37284\
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__37292\,
            I => \N__37272\
        );

    \I__8641\ : InMux
    port map (
            O => \N__37291\,
            I => \N__37262\
        );

    \I__8640\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37262\
        );

    \I__8639\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37262\
        );

    \I__8638\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37262\
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__37283\,
            I => \N__37256\
        );

    \I__8636\ : CascadeMux
    port map (
            O => \N__37282\,
            I => \N__37252\
        );

    \I__8635\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37242\
        );

    \I__8634\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37242\
        );

    \I__8633\ : InMux
    port map (
            O => \N__37279\,
            I => \N__37242\
        );

    \I__8632\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37242\
        );

    \I__8631\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37231\
        );

    \I__8630\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37231\
        );

    \I__8629\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37231\
        );

    \I__8628\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37231\
        );

    \I__8627\ : InMux
    port map (
            O => \N__37271\,
            I => \N__37231\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__37262\,
            I => \N__37228\
        );

    \I__8625\ : CascadeMux
    port map (
            O => \N__37261\,
            I => \N__37224\
        );

    \I__8624\ : InMux
    port map (
            O => \N__37260\,
            I => \N__37219\
        );

    \I__8623\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37214\
        );

    \I__8622\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37214\
        );

    \I__8621\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37211\
        );

    \I__8620\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37208\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__37251\,
            I => \N__37204\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__37242\,
            I => \N__37197\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__37231\,
            I => \N__37197\
        );

    \I__8616\ : Span4Mux_s0_h
    port map (
            O => \N__37228\,
            I => \N__37197\
        );

    \I__8615\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37192\
        );

    \I__8614\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37192\
        );

    \I__8613\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37187\
        );

    \I__8612\ : InMux
    port map (
            O => \N__37222\,
            I => \N__37187\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__37219\,
            I => \N__37178\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37178\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__37211\,
            I => \N__37178\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__37208\,
            I => \N__37178\
        );

    \I__8607\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37175\
        );

    \I__8606\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37172\
        );

    \I__8605\ : Span4Mux_h
    port map (
            O => \N__37197\,
            I => \N__37169\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37164\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__37187\,
            I => \N__37164\
        );

    \I__8602\ : Span12Mux_s5_h
    port map (
            O => \N__37178\,
            I => \N__37161\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__37175\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__37172\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__37169\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__8598\ : Odrv12
    port map (
            O => \N__37164\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__8597\ : Odrv12
    port map (
            O => \N__37161\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__37150\,
            I => \N__37138\
        );

    \I__8595\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37135\
        );

    \I__8594\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37132\
        );

    \I__8593\ : InMux
    port map (
            O => \N__37147\,
            I => \N__37129\
        );

    \I__8592\ : InMux
    port map (
            O => \N__37146\,
            I => \N__37126\
        );

    \I__8591\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37122\
        );

    \I__8590\ : InMux
    port map (
            O => \N__37144\,
            I => \N__37116\
        );

    \I__8589\ : InMux
    port map (
            O => \N__37143\,
            I => \N__37116\
        );

    \I__8588\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37111\
        );

    \I__8587\ : InMux
    port map (
            O => \N__37141\,
            I => \N__37111\
        );

    \I__8586\ : InMux
    port map (
            O => \N__37138\,
            I => \N__37107\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__37135\,
            I => \N__37100\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__37132\,
            I => \N__37100\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__37129\,
            I => \N__37100\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__37126\,
            I => \N__37097\
        );

    \I__8581\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37094\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37091\
        );

    \I__8579\ : InMux
    port map (
            O => \N__37121\,
            I => \N__37088\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37083\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__37111\,
            I => \N__37083\
        );

    \I__8576\ : InMux
    port map (
            O => \N__37110\,
            I => \N__37080\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__37107\,
            I => \N__37077\
        );

    \I__8574\ : Span4Mux_v
    port map (
            O => \N__37100\,
            I => \N__37070\
        );

    \I__8573\ : Span4Mux_h
    port map (
            O => \N__37097\,
            I => \N__37070\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__37094\,
            I => \N__37070\
        );

    \I__8571\ : Span4Mux_v
    port map (
            O => \N__37091\,
            I => \N__37063\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__37088\,
            I => \N__37063\
        );

    \I__8569\ : Span4Mux_v
    port map (
            O => \N__37083\,
            I => \N__37063\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__37080\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__37077\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__37070\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__37063\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__8564\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37051\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__37051\,
            I => \POWERLED.un1_dutycycle_53_34_1\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__37048\,
            I => \POWERLED.un1_dutycycle_53_36_0_cascade_\
        );

    \I__8561\ : InMux
    port map (
            O => \N__37045\,
            I => \N__37042\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__37042\,
            I => \POWERLED.un1_dutycycle_53_34_0\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__37039\,
            I => \N__37036\
        );

    \I__8558\ : InMux
    port map (
            O => \N__37036\,
            I => \N__37033\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__37030\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__37030\,
            I => \N__37027\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__37027\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_12\
        );

    \I__8554\ : CascadeMux
    port map (
            O => \N__37024\,
            I => \POWERLED.un1_dutycycle_53_4_a0_1_cascade_\
        );

    \I__8553\ : InMux
    port map (
            O => \N__37021\,
            I => \N__37018\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__37018\,
            I => \POWERLED.un1_dutycycle_53_9_3\
        );

    \I__8551\ : CascadeMux
    port map (
            O => \N__37015\,
            I => \N__37012\
        );

    \I__8550\ : InMux
    port map (
            O => \N__37012\,
            I => \N__37009\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__37009\,
            I => \N__36999\
        );

    \I__8548\ : InMux
    port map (
            O => \N__37008\,
            I => \N__36996\
        );

    \I__8547\ : InMux
    port map (
            O => \N__37007\,
            I => \N__36993\
        );

    \I__8546\ : InMux
    port map (
            O => \N__37006\,
            I => \N__36990\
        );

    \I__8545\ : InMux
    port map (
            O => \N__37005\,
            I => \N__36987\
        );

    \I__8544\ : CascadeMux
    port map (
            O => \N__37004\,
            I => \N__36984\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__37003\,
            I => \N__36979\
        );

    \I__8542\ : CascadeMux
    port map (
            O => \N__37002\,
            I => \N__36974\
        );

    \I__8541\ : Span4Mux_v
    port map (
            O => \N__36999\,
            I => \N__36968\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__36996\,
            I => \N__36968\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36965\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__36990\,
            I => \N__36960\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__36987\,
            I => \N__36960\
        );

    \I__8536\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36957\
        );

    \I__8535\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36952\
        );

    \I__8534\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36952\
        );

    \I__8533\ : InMux
    port map (
            O => \N__36979\,
            I => \N__36947\
        );

    \I__8532\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36947\
        );

    \I__8531\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36940\
        );

    \I__8530\ : InMux
    port map (
            O => \N__36974\,
            I => \N__36940\
        );

    \I__8529\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36940\
        );

    \I__8528\ : Span4Mux_s3_h
    port map (
            O => \N__36968\,
            I => \N__36935\
        );

    \I__8527\ : Span4Mux_s3_h
    port map (
            O => \N__36965\,
            I => \N__36935\
        );

    \I__8526\ : Span4Mux_s3_h
    port map (
            O => \N__36960\,
            I => \N__36932\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__36957\,
            I => \N__36929\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__36952\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__36947\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__36940\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__36935\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__36932\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__36929\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__8518\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36913\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__36913\,
            I => \POWERLED.un1_dutycycle_53_31_a1_2\
        );

    \I__8516\ : CascadeMux
    port map (
            O => \N__36910\,
            I => \POWERLED.un1_dutycycle_53_9_5_1_cascade_\
        );

    \I__8515\ : InMux
    port map (
            O => \N__36907\,
            I => \N__36904\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__36904\,
            I => \POWERLED.un1_dutycycle_53_9_5\
        );

    \I__8513\ : CascadeMux
    port map (
            O => \N__36901\,
            I => \POWERLED.un1_dutycycle_53_31_a7_0_cascade_\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__36898\,
            I => \N__36895\
        );

    \I__8511\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36889\
        );

    \I__8510\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36889\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__36889\,
            I => \POWERLED.un1_dutycycle_53_4_a0_1\
        );

    \I__8508\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36883\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__36883\,
            I => \POWERLED.dutycycle_RNIZ0Z_6\
        );

    \I__8506\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36856\
        );

    \I__8505\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36856\
        );

    \I__8504\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36856\
        );

    \I__8503\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36856\
        );

    \I__8502\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36849\
        );

    \I__8501\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36849\
        );

    \I__8500\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36839\
        );

    \I__8499\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36839\
        );

    \I__8498\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36839\
        );

    \I__8497\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36832\
        );

    \I__8496\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36832\
        );

    \I__8495\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36832\
        );

    \I__8494\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36827\
        );

    \I__8493\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36827\
        );

    \I__8492\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36824\
        );

    \I__8491\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36819\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__36856\,
            I => \N__36816\
        );

    \I__8489\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36811\
        );

    \I__8488\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36811\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__36849\,
            I => \N__36808\
        );

    \I__8486\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36801\
        );

    \I__8485\ : InMux
    port map (
            O => \N__36847\,
            I => \N__36801\
        );

    \I__8484\ : InMux
    port map (
            O => \N__36846\,
            I => \N__36801\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__36839\,
            I => \N__36798\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__36832\,
            I => \N__36793\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__36827\,
            I => \N__36793\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__36824\,
            I => \N__36790\
        );

    \I__8479\ : InMux
    port map (
            O => \N__36823\,
            I => \N__36781\
        );

    \I__8478\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36781\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__36819\,
            I => \N__36776\
        );

    \I__8476\ : Span4Mux_s2_v
    port map (
            O => \N__36816\,
            I => \N__36776\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__36811\,
            I => \N__36773\
        );

    \I__8474\ : Span4Mux_s0_h
    port map (
            O => \N__36808\,
            I => \N__36766\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__36801\,
            I => \N__36766\
        );

    \I__8472\ : Span4Mux_s2_v
    port map (
            O => \N__36798\,
            I => \N__36766\
        );

    \I__8471\ : Span4Mux_v
    port map (
            O => \N__36793\,
            I => \N__36761\
        );

    \I__8470\ : Span4Mux_s1_h
    port map (
            O => \N__36790\,
            I => \N__36761\
        );

    \I__8469\ : CascadeMux
    port map (
            O => \N__36789\,
            I => \N__36758\
        );

    \I__8468\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36750\
        );

    \I__8467\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36750\
        );

    \I__8466\ : InMux
    port map (
            O => \N__36786\,
            I => \N__36747\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__36781\,
            I => \N__36742\
        );

    \I__8464\ : Span4Mux_s2_h
    port map (
            O => \N__36776\,
            I => \N__36742\
        );

    \I__8463\ : Span4Mux_s2_v
    port map (
            O => \N__36773\,
            I => \N__36737\
        );

    \I__8462\ : Span4Mux_h
    port map (
            O => \N__36766\,
            I => \N__36737\
        );

    \I__8461\ : Span4Mux_h
    port map (
            O => \N__36761\,
            I => \N__36734\
        );

    \I__8460\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36729\
        );

    \I__8459\ : InMux
    port map (
            O => \N__36757\,
            I => \N__36729\
        );

    \I__8458\ : InMux
    port map (
            O => \N__36756\,
            I => \N__36726\
        );

    \I__8457\ : InMux
    port map (
            O => \N__36755\,
            I => \N__36723\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__36750\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__36747\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__36742\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8453\ : Odrv4
    port map (
            O => \N__36737\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8452\ : Odrv4
    port map (
            O => \N__36734\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__36729\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__36726\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__36723\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__8448\ : CascadeMux
    port map (
            O => \N__36706\,
            I => \N__36703\
        );

    \I__8447\ : InMux
    port map (
            O => \N__36703\,
            I => \N__36694\
        );

    \I__8446\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36687\
        );

    \I__8445\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36684\
        );

    \I__8444\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36675\
        );

    \I__8443\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36675\
        );

    \I__8442\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36675\
        );

    \I__8441\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36672\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__36694\,
            I => \N__36669\
        );

    \I__8439\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36666\
        );

    \I__8438\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36661\
        );

    \I__8437\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36661\
        );

    \I__8436\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36656\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__36687\,
            I => \N__36644\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__36684\,
            I => \N__36641\
        );

    \I__8433\ : InMux
    port map (
            O => \N__36683\,
            I => \N__36636\
        );

    \I__8432\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36636\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__36675\,
            I => \N__36633\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__36672\,
            I => \N__36628\
        );

    \I__8429\ : Span4Mux_s1_v
    port map (
            O => \N__36669\,
            I => \N__36628\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__36666\,
            I => \N__36623\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__36661\,
            I => \N__36623\
        );

    \I__8426\ : InMux
    port map (
            O => \N__36660\,
            I => \N__36618\
        );

    \I__8425\ : InMux
    port map (
            O => \N__36659\,
            I => \N__36618\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36615\
        );

    \I__8423\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36612\
        );

    \I__8422\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36603\
        );

    \I__8421\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36603\
        );

    \I__8420\ : InMux
    port map (
            O => \N__36652\,
            I => \N__36603\
        );

    \I__8419\ : InMux
    port map (
            O => \N__36651\,
            I => \N__36603\
        );

    \I__8418\ : InMux
    port map (
            O => \N__36650\,
            I => \N__36598\
        );

    \I__8417\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36598\
        );

    \I__8416\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36593\
        );

    \I__8415\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36593\
        );

    \I__8414\ : Span12Mux_s8_h
    port map (
            O => \N__36644\,
            I => \N__36590\
        );

    \I__8413\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36577\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__36636\,
            I => \N__36577\
        );

    \I__8411\ : Span4Mux_v
    port map (
            O => \N__36633\,
            I => \N__36577\
        );

    \I__8410\ : Span4Mux_s0_h
    port map (
            O => \N__36628\,
            I => \N__36577\
        );

    \I__8409\ : Span4Mux_v
    port map (
            O => \N__36623\,
            I => \N__36577\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__36618\,
            I => \N__36577\
        );

    \I__8407\ : Odrv12
    port map (
            O => \N__36615\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__36612\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__36603\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__36598\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__36593\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8402\ : Odrv12
    port map (
            O => \N__36590\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__36577\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__8400\ : CascadeMux
    port map (
            O => \N__36562\,
            I => \N__36552\
        );

    \I__8399\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36548\
        );

    \I__8398\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36543\
        );

    \I__8397\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36543\
        );

    \I__8396\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36538\
        );

    \I__8395\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36538\
        );

    \I__8394\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36531\
        );

    \I__8393\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36531\
        );

    \I__8392\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36531\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__36551\,
            I => \N__36527\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__36548\,
            I => \N__36524\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__36543\,
            I => \N__36519\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__36538\,
            I => \N__36514\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__36531\,
            I => \N__36514\
        );

    \I__8386\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36511\
        );

    \I__8385\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36508\
        );

    \I__8384\ : Span4Mux_s2_v
    port map (
            O => \N__36524\,
            I => \N__36505\
        );

    \I__8383\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36500\
        );

    \I__8382\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36500\
        );

    \I__8381\ : Span4Mux_s2_v
    port map (
            O => \N__36519\,
            I => \N__36495\
        );

    \I__8380\ : Span4Mux_s2_v
    port map (
            O => \N__36514\,
            I => \N__36495\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36486\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__36508\,
            I => \N__36486\
        );

    \I__8377\ : Sp12to4
    port map (
            O => \N__36505\,
            I => \N__36486\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__36500\,
            I => \N__36486\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__36495\,
            I => \N__36483\
        );

    \I__8374\ : Odrv12
    port map (
            O => \N__36486\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_7\
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__36483\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_7\
        );

    \I__8372\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36475\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__36475\,
            I => \POWERLED.un1_dutycycle_53_39_c_1\
        );

    \I__8370\ : CascadeMux
    port map (
            O => \N__36472\,
            I => \N__36466\
        );

    \I__8369\ : InMux
    port map (
            O => \N__36471\,
            I => \N__36457\
        );

    \I__8368\ : InMux
    port map (
            O => \N__36470\,
            I => \N__36453\
        );

    \I__8367\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36450\
        );

    \I__8366\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36447\
        );

    \I__8365\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36444\
        );

    \I__8364\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36439\
        );

    \I__8363\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36439\
        );

    \I__8362\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36434\
        );

    \I__8361\ : InMux
    port map (
            O => \N__36461\,
            I => \N__36429\
        );

    \I__8360\ : InMux
    port map (
            O => \N__36460\,
            I => \N__36429\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__36457\,
            I => \N__36426\
        );

    \I__8358\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36423\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__36453\,
            I => \N__36420\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__36450\,
            I => \N__36416\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36413\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__36444\,
            I => \N__36410\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__36439\,
            I => \N__36407\
        );

    \I__8352\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36402\
        );

    \I__8351\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36402\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36391\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__36429\,
            I => \N__36391\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__36426\,
            I => \N__36391\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__36423\,
            I => \N__36391\
        );

    \I__8346\ : Span4Mux_s0_h
    port map (
            O => \N__36420\,
            I => \N__36391\
        );

    \I__8345\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36388\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__36416\,
            I => \N__36385\
        );

    \I__8343\ : Span4Mux_v
    port map (
            O => \N__36413\,
            I => \N__36378\
        );

    \I__8342\ : Span4Mux_v
    port map (
            O => \N__36410\,
            I => \N__36378\
        );

    \I__8341\ : Span4Mux_s1_h
    port map (
            O => \N__36407\,
            I => \N__36378\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__36402\,
            I => \N__36375\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__36391\,
            I => \N__36372\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__36388\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__8337\ : Odrv4
    port map (
            O => \N__36385\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__8336\ : Odrv4
    port map (
            O => \N__36378\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__36375\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__8334\ : Odrv4
    port map (
            O => \N__36372\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__36361\,
            I => \N__36358\
        );

    \I__8332\ : InMux
    port map (
            O => \N__36358\,
            I => \N__36355\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__36355\,
            I => \POWERLED.un1_dutycycle_53_49_0_0\
        );

    \I__8330\ : InMux
    port map (
            O => \N__36352\,
            I => \N__36348\
        );

    \I__8329\ : InMux
    port map (
            O => \N__36351\,
            I => \N__36345\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__36348\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_9\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__36345\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_9\
        );

    \I__8326\ : InMux
    port map (
            O => \N__36340\,
            I => \N__36334\
        );

    \I__8325\ : InMux
    port map (
            O => \N__36339\,
            I => \N__36334\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__36334\,
            I => \N__36331\
        );

    \I__8323\ : Span4Mux_s1_v
    port map (
            O => \N__36331\,
            I => \N__36328\
        );

    \I__8322\ : Odrv4
    port map (
            O => \N__36328\,
            I => \POWERLED.un1_dutycycle_53_49_0\
        );

    \I__8321\ : CascadeMux
    port map (
            O => \N__36325\,
            I => \POWERLED.g3_1_3_0_cascade_\
        );

    \I__8320\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36319\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__36319\,
            I => \POWERLED.g0_10_0_0_0\
        );

    \I__8318\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36313\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__36313\,
            I => \N__36310\
        );

    \I__8316\ : Odrv12
    port map (
            O => \N__36310\,
            I => \POWERLED.N_3034_0_0_0\
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__36307\,
            I => \N__36304\
        );

    \I__8314\ : InMux
    port map (
            O => \N__36304\,
            I => \N__36300\
        );

    \I__8313\ : InMux
    port map (
            O => \N__36303\,
            I => \N__36297\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__36300\,
            I => \N__36294\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__36297\,
            I => \N__36291\
        );

    \I__8310\ : Span4Mux_s2_h
    port map (
            O => \N__36294\,
            I => \N__36288\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__36291\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__8308\ : Odrv4
    port map (
            O => \N__36288\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__8307\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36280\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__36280\,
            I => \N__36277\
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__36277\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__8304\ : InMux
    port map (
            O => \N__36274\,
            I => \N__36270\
        );

    \I__8303\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36267\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__36270\,
            I => \N__36264\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__36267\,
            I => \N__36261\
        );

    \I__8300\ : Span4Mux_s2_h
    port map (
            O => \N__36264\,
            I => \N__36258\
        );

    \I__8299\ : Odrv12
    port map (
            O => \N__36261\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__36258\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__36253\,
            I => \N__36250\
        );

    \I__8296\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36247\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__36247\,
            I => \N__36244\
        );

    \I__8294\ : Odrv4
    port map (
            O => \N__36244\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__8293\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36238\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__36238\,
            I => \N__36232\
        );

    \I__8291\ : CascadeMux
    port map (
            O => \N__36237\,
            I => \N__36229\
        );

    \I__8290\ : CascadeMux
    port map (
            O => \N__36236\,
            I => \N__36226\
        );

    \I__8289\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36222\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__36232\,
            I => \N__36219\
        );

    \I__8287\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36216\
        );

    \I__8286\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36213\
        );

    \I__8285\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36210\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__36222\,
            I => \N__36207\
        );

    \I__8283\ : Odrv4
    port map (
            O => \N__36219\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__36216\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__36213\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__36210\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__36207\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__8278\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36193\
        );

    \I__8277\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36190\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__36190\,
            I => \N__36187\
        );

    \I__8275\ : Span4Mux_h
    port map (
            O => \N__36187\,
            I => \N__36184\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__36184\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__36181\,
            I => \N__36173\
        );

    \I__8272\ : CascadeMux
    port map (
            O => \N__36180\,
            I => \N__36170\
        );

    \I__8271\ : InMux
    port map (
            O => \N__36179\,
            I => \N__36167\
        );

    \I__8270\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36162\
        );

    \I__8269\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36162\
        );

    \I__8268\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36157\
        );

    \I__8267\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36152\
        );

    \I__8266\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36152\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__36167\,
            I => \N__36141\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__36162\,
            I => \N__36141\
        );

    \I__8263\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36138\
        );

    \I__8262\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36135\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__36157\,
            I => \N__36126\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__36152\,
            I => \N__36126\
        );

    \I__8259\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36121\
        );

    \I__8258\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36121\
        );

    \I__8257\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36116\
        );

    \I__8256\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36116\
        );

    \I__8255\ : CascadeMux
    port map (
            O => \N__36147\,
            I => \N__36113\
        );

    \I__8254\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36109\
        );

    \I__8253\ : Span4Mux_s1_h
    port map (
            O => \N__36141\,
            I => \N__36106\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__36138\,
            I => \N__36101\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36101\
        );

    \I__8250\ : InMux
    port map (
            O => \N__36134\,
            I => \N__36094\
        );

    \I__8249\ : InMux
    port map (
            O => \N__36133\,
            I => \N__36094\
        );

    \I__8248\ : InMux
    port map (
            O => \N__36132\,
            I => \N__36094\
        );

    \I__8247\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36091\
        );

    \I__8246\ : Span4Mux_s2_v
    port map (
            O => \N__36126\,
            I => \N__36086\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__36121\,
            I => \N__36086\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__36116\,
            I => \N__36083\
        );

    \I__8243\ : InMux
    port map (
            O => \N__36113\,
            I => \N__36078\
        );

    \I__8242\ : InMux
    port map (
            O => \N__36112\,
            I => \N__36078\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__36109\,
            I => \N__36075\
        );

    \I__8240\ : Span4Mux_h
    port map (
            O => \N__36106\,
            I => \N__36066\
        );

    \I__8239\ : Span4Mux_s3_v
    port map (
            O => \N__36101\,
            I => \N__36066\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__36094\,
            I => \N__36066\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__36091\,
            I => \N__36066\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__36086\,
            I => \N__36059\
        );

    \I__8235\ : Span4Mux_v
    port map (
            O => \N__36083\,
            I => \N__36059\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__36078\,
            I => \N__36059\
        );

    \I__8233\ : Odrv12
    port map (
            O => \N__36075\,
            I => \POWERLED.N_203_i\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__36066\,
            I => \POWERLED.N_203_i\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__36059\,
            I => \POWERLED.N_203_i\
        );

    \I__8230\ : InMux
    port map (
            O => \N__36052\,
            I => \N__36049\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__36049\,
            I => \POWERLED.g0_10_0_0_1\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__36046\,
            I => \N__36041\
        );

    \I__8227\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36038\
        );

    \I__8226\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36032\
        );

    \I__8225\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36032\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__36038\,
            I => \N__36024\
        );

    \I__8223\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36021\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__36032\,
            I => \N__36018\
        );

    \I__8221\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36015\
        );

    \I__8220\ : InMux
    port map (
            O => \N__36030\,
            I => \N__36006\
        );

    \I__8219\ : InMux
    port map (
            O => \N__36029\,
            I => \N__36006\
        );

    \I__8218\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36006\
        );

    \I__8217\ : InMux
    port map (
            O => \N__36027\,
            I => \N__36006\
        );

    \I__8216\ : Span4Mux_s1_v
    port map (
            O => \N__36024\,
            I => \N__36001\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__35996\
        );

    \I__8214\ : Span4Mux_s3_h
    port map (
            O => \N__36018\,
            I => \N__35996\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__36015\,
            I => \N__35991\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__36006\,
            I => \N__35988\
        );

    \I__8211\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35983\
        );

    \I__8210\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35983\
        );

    \I__8209\ : Span4Mux_v
    port map (
            O => \N__36001\,
            I => \N__35980\
        );

    \I__8208\ : Span4Mux_h
    port map (
            O => \N__35996\,
            I => \N__35977\
        );

    \I__8207\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35972\
        );

    \I__8206\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35972\
        );

    \I__8205\ : Span4Mux_h
    port map (
            O => \N__35991\,
            I => \N__35967\
        );

    \I__8204\ : Span4Mux_h
    port map (
            O => \N__35988\,
            I => \N__35967\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__35983\,
            I => \N__35964\
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__35980\,
            I => \POWERLED.N_175\
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__35977\,
            I => \POWERLED.N_175\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__35972\,
            I => \POWERLED.N_175\
        );

    \I__8199\ : Odrv4
    port map (
            O => \N__35967\,
            I => \POWERLED.N_175\
        );

    \I__8198\ : Odrv12
    port map (
            O => \N__35964\,
            I => \POWERLED.N_175\
        );

    \I__8197\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__35950\,
            I => \POWERLED.g3_1_3_0\
        );

    \I__8195\ : InMux
    port map (
            O => \N__35947\,
            I => \N__35944\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__35944\,
            I => \POWERLED.N_3034_0_0_2\
        );

    \I__8193\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35934\
        );

    \I__8191\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35931\
        );

    \I__8190\ : Span4Mux_s2_h
    port map (
            O => \N__35934\,
            I => \N__35928\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__35931\,
            I => \N__35925\
        );

    \I__8188\ : Odrv4
    port map (
            O => \N__35928\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__8187\ : Odrv4
    port map (
            O => \N__35925\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__35920\,
            I => \N__35917\
        );

    \I__8185\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35914\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__35914\,
            I => \N__35911\
        );

    \I__8183\ : Odrv12
    port map (
            O => \N__35911\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__35908\,
            I => \N__35905\
        );

    \I__8181\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35902\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__35902\,
            I => \POWERLED.un1_dutycycle_53_10_4_1\
        );

    \I__8179\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35896\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35893\
        );

    \I__8177\ : Odrv12
    port map (
            O => \N__35893\,
            I => \POWERLED.un1_dutycycle_53_10_4\
        );

    \I__8176\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35887\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__35887\,
            I => \N__35884\
        );

    \I__8174\ : Odrv4
    port map (
            O => \N__35884\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__8173\ : InMux
    port map (
            O => \N__35881\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__8172\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35875\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__35875\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__8170\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35869\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__35869\,
            I => \N__35866\
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__35866\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__8167\ : InMux
    port map (
            O => \N__35863\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__8166\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35857\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__35857\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__35854\,
            I => \N__35851\
        );

    \I__8163\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35848\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__35848\,
            I => \N__35845\
        );

    \I__8161\ : Span4Mux_v
    port map (
            O => \N__35845\,
            I => \N__35842\
        );

    \I__8160\ : Odrv4
    port map (
            O => \N__35842\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__8159\ : InMux
    port map (
            O => \N__35839\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__8158\ : InMux
    port map (
            O => \N__35836\,
            I => \N__35833\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__35833\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__8156\ : CascadeMux
    port map (
            O => \N__35830\,
            I => \N__35827\
        );

    \I__8155\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35824\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__35824\,
            I => \N__35821\
        );

    \I__8153\ : Span4Mux_v
    port map (
            O => \N__35821\,
            I => \N__35818\
        );

    \I__8152\ : Odrv4
    port map (
            O => \N__35818\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__8151\ : InMux
    port map (
            O => \N__35815\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__35812\,
            I => \N__35808\
        );

    \I__8149\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35800\
        );

    \I__8148\ : InMux
    port map (
            O => \N__35808\,
            I => \N__35800\
        );

    \I__8147\ : InMux
    port map (
            O => \N__35807\,
            I => \N__35800\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__35800\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__8145\ : CascadeMux
    port map (
            O => \N__35797\,
            I => \N__35794\
        );

    \I__8144\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35791\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__35791\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__8142\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35785\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__35785\,
            I => \N__35782\
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__35782\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__8139\ : InMux
    port map (
            O => \N__35779\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__8138\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35773\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__35773\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__8136\ : InMux
    port map (
            O => \N__35770\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__8135\ : CascadeMux
    port map (
            O => \N__35767\,
            I => \N__35763\
        );

    \I__8134\ : InMux
    port map (
            O => \N__35766\,
            I => \N__35758\
        );

    \I__8133\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35758\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35753\
        );

    \I__8131\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35750\
        );

    \I__8130\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35747\
        );

    \I__8129\ : Odrv4
    port map (
            O => \N__35753\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__35750\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__35747\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__8126\ : CascadeMux
    port map (
            O => \N__35740\,
            I => \POWERLED.mult1_un68_sum_s_8_cascade_\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__35737\,
            I => \N__35733\
        );

    \I__8124\ : InMux
    port map (
            O => \N__35736\,
            I => \N__35725\
        );

    \I__8123\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35725\
        );

    \I__8122\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35725\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35722\
        );

    \I__8120\ : Odrv4
    port map (
            O => \N__35722\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__8119\ : CascadeMux
    port map (
            O => \N__35719\,
            I => \N__35716\
        );

    \I__8118\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35713\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35710\
        );

    \I__8116\ : Span4Mux_s2_h
    port map (
            O => \N__35710\,
            I => \N__35707\
        );

    \I__8115\ : Span4Mux_v
    port map (
            O => \N__35707\,
            I => \N__35704\
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__35704\,
            I => \POWERLED.g0_7_1\
        );

    \I__8113\ : CascadeMux
    port map (
            O => \N__35701\,
            I => \N__35694\
        );

    \I__8112\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35689\
        );

    \I__8111\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35686\
        );

    \I__8110\ : InMux
    port map (
            O => \N__35698\,
            I => \N__35680\
        );

    \I__8109\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35677\
        );

    \I__8108\ : InMux
    port map (
            O => \N__35694\,
            I => \N__35670\
        );

    \I__8107\ : InMux
    port map (
            O => \N__35693\,
            I => \N__35670\
        );

    \I__8106\ : InMux
    port map (
            O => \N__35692\,
            I => \N__35670\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35667\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__35686\,
            I => \N__35664\
        );

    \I__8103\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35661\
        );

    \I__8102\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35658\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__35683\,
            I => \N__35651\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35648\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__35677\,
            I => \N__35643\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__35670\,
            I => \N__35643\
        );

    \I__8097\ : Span4Mux_h
    port map (
            O => \N__35667\,
            I => \N__35640\
        );

    \I__8096\ : Span4Mux_v
    port map (
            O => \N__35664\,
            I => \N__35633\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__35661\,
            I => \N__35633\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__35658\,
            I => \N__35633\
        );

    \I__8093\ : InMux
    port map (
            O => \N__35657\,
            I => \N__35630\
        );

    \I__8092\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35627\
        );

    \I__8091\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35624\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__35654\,
            I => \N__35621\
        );

    \I__8089\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35618\
        );

    \I__8088\ : Span12Mux_v
    port map (
            O => \N__35648\,
            I => \N__35615\
        );

    \I__8087\ : Span12Mux_s7_h
    port map (
            O => \N__35643\,
            I => \N__35612\
        );

    \I__8086\ : Span4Mux_v
    port map (
            O => \N__35640\,
            I => \N__35607\
        );

    \I__8085\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35607\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35600\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__35627\,
            I => \N__35600\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__35624\,
            I => \N__35600\
        );

    \I__8081\ : InMux
    port map (
            O => \N__35621\,
            I => \N__35597\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__35618\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__8079\ : Odrv12
    port map (
            O => \N__35615\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__8078\ : Odrv12
    port map (
            O => \N__35612\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__8077\ : Odrv4
    port map (
            O => \N__35607\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__8076\ : Odrv4
    port map (
            O => \N__35600\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__35597\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__8074\ : InMux
    port map (
            O => \N__35584\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__35581\,
            I => \N__35578\
        );

    \I__8072\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35575\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__35575\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__8070\ : InMux
    port map (
            O => \N__35572\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__8069\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35566\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__35566\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__8067\ : InMux
    port map (
            O => \N__35563\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__35560\,
            I => \N__35556\
        );

    \I__8065\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35550\
        );

    \I__8064\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35550\
        );

    \I__8063\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35547\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__35550\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__35547\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__35542\,
            I => \N__35539\
        );

    \I__8059\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35536\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__35536\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__8057\ : InMux
    port map (
            O => \N__35533\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__8056\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35527\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__35527\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__35524\,
            I => \N__35520\
        );

    \I__8053\ : CascadeMux
    port map (
            O => \N__35523\,
            I => \N__35516\
        );

    \I__8052\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35509\
        );

    \I__8051\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35509\
        );

    \I__8050\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35509\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__35509\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__8048\ : InMux
    port map (
            O => \N__35506\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__35503\,
            I => \N__35500\
        );

    \I__8046\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35497\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__35497\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__8044\ : InMux
    port map (
            O => \N__35494\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__35491\,
            I => \N__35488\
        );

    \I__8042\ : InMux
    port map (
            O => \N__35488\,
            I => \N__35485\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__35485\,
            I => \N__35482\
        );

    \I__8040\ : Span4Mux_h
    port map (
            O => \N__35482\,
            I => \N__35479\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__35479\,
            I => \POWERLED.mult1_un68_sum_i_8\
        );

    \I__8038\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35472\
        );

    \I__8037\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35469\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__35472\,
            I => \N__35464\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35464\
        );

    \I__8034\ : Span4Mux_v
    port map (
            O => \N__35464\,
            I => \N__35461\
        );

    \I__8033\ : Odrv4
    port map (
            O => \N__35461\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__8032\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35455\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__35455\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__8030\ : InMux
    port map (
            O => \N__35452\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__8029\ : CascadeMux
    port map (
            O => \N__35449\,
            I => \N__35446\
        );

    \I__8028\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35443\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__35443\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__8026\ : InMux
    port map (
            O => \N__35440\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__8025\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35434\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__35434\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__8023\ : InMux
    port map (
            O => \N__35431\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__8022\ : CascadeMux
    port map (
            O => \N__35428\,
            I => \N__35425\
        );

    \I__8021\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35422\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__35422\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__8019\ : InMux
    port map (
            O => \N__35419\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__8018\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35413\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__35413\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__8016\ : InMux
    port map (
            O => \N__35410\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__8015\ : InMux
    port map (
            O => \N__35407\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__8014\ : InMux
    port map (
            O => \N__35404\,
            I => \N__35401\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__35401\,
            I => \N__35397\
        );

    \I__8012\ : CascadeMux
    port map (
            O => \N__35400\,
            I => \N__35394\
        );

    \I__8011\ : Span4Mux_h
    port map (
            O => \N__35397\,
            I => \N__35388\
        );

    \I__8010\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35381\
        );

    \I__8009\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35381\
        );

    \I__8008\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35381\
        );

    \I__8007\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35378\
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__35388\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__35381\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__35378\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__35371\,
            I => \N__35368\
        );

    \I__8002\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35365\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__35365\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__8000\ : InMux
    port map (
            O => \N__35362\,
            I => \N__35358\
        );

    \I__7999\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35355\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35350\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__35355\,
            I => \N__35350\
        );

    \I__7996\ : Odrv4
    port map (
            O => \N__35350\,
            I => \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3\
        );

    \I__7995\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35344\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__35344\,
            I => \HDA_STRAP.count_1_14\
        );

    \I__7993\ : ClkMux
    port map (
            O => \N__35341\,
            I => \N__35333\
        );

    \I__7992\ : ClkMux
    port map (
            O => \N__35340\,
            I => \N__35329\
        );

    \I__7991\ : ClkMux
    port map (
            O => \N__35339\,
            I => \N__35326\
        );

    \I__7990\ : ClkMux
    port map (
            O => \N__35338\,
            I => \N__35323\
        );

    \I__7989\ : ClkMux
    port map (
            O => \N__35337\,
            I => \N__35308\
        );

    \I__7988\ : ClkMux
    port map (
            O => \N__35336\,
            I => \N__35304\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__35333\,
            I => \N__35300\
        );

    \I__7986\ : ClkMux
    port map (
            O => \N__35332\,
            I => \N__35297\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__35329\,
            I => \N__35292\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35292\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__35323\,
            I => \N__35289\
        );

    \I__7982\ : ClkMux
    port map (
            O => \N__35322\,
            I => \N__35286\
        );

    \I__7981\ : ClkMux
    port map (
            O => \N__35321\,
            I => \N__35283\
        );

    \I__7980\ : ClkMux
    port map (
            O => \N__35320\,
            I => \N__35278\
        );

    \I__7979\ : ClkMux
    port map (
            O => \N__35319\,
            I => \N__35273\
        );

    \I__7978\ : ClkMux
    port map (
            O => \N__35318\,
            I => \N__35270\
        );

    \I__7977\ : ClkMux
    port map (
            O => \N__35317\,
            I => \N__35267\
        );

    \I__7976\ : ClkMux
    port map (
            O => \N__35316\,
            I => \N__35264\
        );

    \I__7975\ : ClkMux
    port map (
            O => \N__35315\,
            I => \N__35261\
        );

    \I__7974\ : ClkMux
    port map (
            O => \N__35314\,
            I => \N__35255\
        );

    \I__7973\ : ClkMux
    port map (
            O => \N__35313\,
            I => \N__35251\
        );

    \I__7972\ : ClkMux
    port map (
            O => \N__35312\,
            I => \N__35247\
        );

    \I__7971\ : ClkMux
    port map (
            O => \N__35311\,
            I => \N__35244\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__35308\,
            I => \N__35239\
        );

    \I__7969\ : ClkMux
    port map (
            O => \N__35307\,
            I => \N__35236\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__35304\,
            I => \N__35232\
        );

    \I__7967\ : ClkMux
    port map (
            O => \N__35303\,
            I => \N__35229\
        );

    \I__7966\ : Span4Mux_s3_v
    port map (
            O => \N__35300\,
            I => \N__35224\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35221\
        );

    \I__7964\ : Span4Mux_s3_v
    port map (
            O => \N__35292\,
            I => \N__35206\
        );

    \I__7963\ : Span4Mux_s1_h
    port map (
            O => \N__35289\,
            I => \N__35206\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__35286\,
            I => \N__35206\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__35283\,
            I => \N__35206\
        );

    \I__7960\ : ClkMux
    port map (
            O => \N__35282\,
            I => \N__35203\
        );

    \I__7959\ : ClkMux
    port map (
            O => \N__35281\,
            I => \N__35200\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__35278\,
            I => \N__35194\
        );

    \I__7957\ : ClkMux
    port map (
            O => \N__35277\,
            I => \N__35191\
        );

    \I__7956\ : ClkMux
    port map (
            O => \N__35276\,
            I => \N__35188\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35184\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35181\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35178\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__35264\,
            I => \N__35170\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35170\
        );

    \I__7950\ : ClkMux
    port map (
            O => \N__35260\,
            I => \N__35167\
        );

    \I__7949\ : ClkMux
    port map (
            O => \N__35259\,
            I => \N__35164\
        );

    \I__7948\ : ClkMux
    port map (
            O => \N__35258\,
            I => \N__35161\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__35255\,
            I => \N__35156\
        );

    \I__7946\ : ClkMux
    port map (
            O => \N__35254\,
            I => \N__35153\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35148\
        );

    \I__7944\ : ClkMux
    port map (
            O => \N__35250\,
            I => \N__35145\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__35247\,
            I => \N__35142\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__35244\,
            I => \N__35139\
        );

    \I__7941\ : ClkMux
    port map (
            O => \N__35243\,
            I => \N__35136\
        );

    \I__7940\ : ClkMux
    port map (
            O => \N__35242\,
            I => \N__35133\
        );

    \I__7939\ : Span4Mux_s2_v
    port map (
            O => \N__35239\,
            I => \N__35126\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__35236\,
            I => \N__35126\
        );

    \I__7937\ : ClkMux
    port map (
            O => \N__35235\,
            I => \N__35123\
        );

    \I__7936\ : Span4Mux_s1_v
    port map (
            O => \N__35232\,
            I => \N__35115\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__35229\,
            I => \N__35115\
        );

    \I__7934\ : ClkMux
    port map (
            O => \N__35228\,
            I => \N__35112\
        );

    \I__7933\ : ClkMux
    port map (
            O => \N__35227\,
            I => \N__35109\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__35224\,
            I => \N__35103\
        );

    \I__7931\ : Span4Mux_s3_v
    port map (
            O => \N__35221\,
            I => \N__35103\
        );

    \I__7930\ : ClkMux
    port map (
            O => \N__35220\,
            I => \N__35100\
        );

    \I__7929\ : ClkMux
    port map (
            O => \N__35219\,
            I => \N__35097\
        );

    \I__7928\ : ClkMux
    port map (
            O => \N__35218\,
            I => \N__35094\
        );

    \I__7927\ : ClkMux
    port map (
            O => \N__35217\,
            I => \N__35089\
        );

    \I__7926\ : ClkMux
    port map (
            O => \N__35216\,
            I => \N__35085\
        );

    \I__7925\ : ClkMux
    port map (
            O => \N__35215\,
            I => \N__35076\
        );

    \I__7924\ : Span4Mux_v
    port map (
            O => \N__35206\,
            I => \N__35068\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35068\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__35200\,
            I => \N__35068\
        );

    \I__7921\ : ClkMux
    port map (
            O => \N__35199\,
            I => \N__35065\
        );

    \I__7920\ : ClkMux
    port map (
            O => \N__35198\,
            I => \N__35062\
        );

    \I__7919\ : ClkMux
    port map (
            O => \N__35197\,
            I => \N__35059\
        );

    \I__7918\ : Span4Mux_h
    port map (
            O => \N__35194\,
            I => \N__35053\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__35191\,
            I => \N__35053\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__35188\,
            I => \N__35050\
        );

    \I__7915\ : ClkMux
    port map (
            O => \N__35187\,
            I => \N__35047\
        );

    \I__7914\ : Span4Mux_s3_v
    port map (
            O => \N__35184\,
            I => \N__35038\
        );

    \I__7913\ : Span4Mux_s3_v
    port map (
            O => \N__35181\,
            I => \N__35038\
        );

    \I__7912\ : Span4Mux_h
    port map (
            O => \N__35178\,
            I => \N__35038\
        );

    \I__7911\ : ClkMux
    port map (
            O => \N__35177\,
            I => \N__35035\
        );

    \I__7910\ : ClkMux
    port map (
            O => \N__35176\,
            I => \N__35032\
        );

    \I__7909\ : ClkMux
    port map (
            O => \N__35175\,
            I => \N__35029\
        );

    \I__7908\ : Span4Mux_v
    port map (
            O => \N__35170\,
            I => \N__35020\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__35167\,
            I => \N__35020\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__35164\,
            I => \N__35020\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__35161\,
            I => \N__35020\
        );

    \I__7904\ : ClkMux
    port map (
            O => \N__35160\,
            I => \N__35014\
        );

    \I__7903\ : ClkMux
    port map (
            O => \N__35159\,
            I => \N__35011\
        );

    \I__7902\ : Span4Mux_s1_h
    port map (
            O => \N__35156\,
            I => \N__35005\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__35153\,
            I => \N__35005\
        );

    \I__7900\ : ClkMux
    port map (
            O => \N__35152\,
            I => \N__35002\
        );

    \I__7899\ : ClkMux
    port map (
            O => \N__35151\,
            I => \N__34998\
        );

    \I__7898\ : Span4Mux_s2_h
    port map (
            O => \N__35148\,
            I => \N__34993\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__35145\,
            I => \N__34993\
        );

    \I__7896\ : Span4Mux_h
    port map (
            O => \N__35142\,
            I => \N__34987\
        );

    \I__7895\ : Span4Mux_s2_v
    port map (
            O => \N__35139\,
            I => \N__34982\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__35136\,
            I => \N__34982\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__35133\,
            I => \N__34979\
        );

    \I__7892\ : ClkMux
    port map (
            O => \N__35132\,
            I => \N__34976\
        );

    \I__7891\ : ClkMux
    port map (
            O => \N__35131\,
            I => \N__34973\
        );

    \I__7890\ : Span4Mux_v
    port map (
            O => \N__35126\,
            I => \N__34970\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__35123\,
            I => \N__34967\
        );

    \I__7888\ : ClkMux
    port map (
            O => \N__35122\,
            I => \N__34964\
        );

    \I__7887\ : ClkMux
    port map (
            O => \N__35121\,
            I => \N__34961\
        );

    \I__7886\ : ClkMux
    port map (
            O => \N__35120\,
            I => \N__34958\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__35115\,
            I => \N__34955\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__35112\,
            I => \N__34952\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__35109\,
            I => \N__34949\
        );

    \I__7882\ : ClkMux
    port map (
            O => \N__35108\,
            I => \N__34946\
        );

    \I__7881\ : Span4Mux_v
    port map (
            O => \N__35103\,
            I => \N__34940\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__35100\,
            I => \N__34940\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__35097\,
            I => \N__34935\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__35094\,
            I => \N__34935\
        );

    \I__7877\ : ClkMux
    port map (
            O => \N__35093\,
            I => \N__34932\
        );

    \I__7876\ : ClkMux
    port map (
            O => \N__35092\,
            I => \N__34929\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__35089\,
            I => \N__34926\
        );

    \I__7874\ : ClkMux
    port map (
            O => \N__35088\,
            I => \N__34923\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__35085\,
            I => \N__34920\
        );

    \I__7872\ : ClkMux
    port map (
            O => \N__35084\,
            I => \N__34917\
        );

    \I__7871\ : ClkMux
    port map (
            O => \N__35083\,
            I => \N__34914\
        );

    \I__7870\ : ClkMux
    port map (
            O => \N__35082\,
            I => \N__34911\
        );

    \I__7869\ : ClkMux
    port map (
            O => \N__35081\,
            I => \N__34908\
        );

    \I__7868\ : ClkMux
    port map (
            O => \N__35080\,
            I => \N__34905\
        );

    \I__7867\ : ClkMux
    port map (
            O => \N__35079\,
            I => \N__34902\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__34899\
        );

    \I__7865\ : ClkMux
    port map (
            O => \N__35075\,
            I => \N__34896\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__35068\,
            I => \N__34886\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__35065\,
            I => \N__34886\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__34886\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__35059\,
            I => \N__34886\
        );

    \I__7860\ : ClkMux
    port map (
            O => \N__35058\,
            I => \N__34883\
        );

    \I__7859\ : Span4Mux_v
    port map (
            O => \N__35053\,
            I => \N__34876\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__35050\,
            I => \N__34876\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__35047\,
            I => \N__34876\
        );

    \I__7856\ : ClkMux
    port map (
            O => \N__35046\,
            I => \N__34873\
        );

    \I__7855\ : ClkMux
    port map (
            O => \N__35045\,
            I => \N__34870\
        );

    \I__7854\ : Span4Mux_v
    port map (
            O => \N__35038\,
            I => \N__34863\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__34863\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__35032\,
            I => \N__34863\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__35029\,
            I => \N__34860\
        );

    \I__7850\ : Span4Mux_v
    port map (
            O => \N__35020\,
            I => \N__34857\
        );

    \I__7849\ : ClkMux
    port map (
            O => \N__35019\,
            I => \N__34854\
        );

    \I__7848\ : ClkMux
    port map (
            O => \N__35018\,
            I => \N__34851\
        );

    \I__7847\ : ClkMux
    port map (
            O => \N__35017\,
            I => \N__34847\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34842\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__35011\,
            I => \N__34842\
        );

    \I__7844\ : ClkMux
    port map (
            O => \N__35010\,
            I => \N__34839\
        );

    \I__7843\ : Span4Mux_h
    port map (
            O => \N__35005\,
            I => \N__34834\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__35002\,
            I => \N__34834\
        );

    \I__7841\ : ClkMux
    port map (
            O => \N__35001\,
            I => \N__34831\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__34998\,
            I => \N__34828\
        );

    \I__7839\ : Span4Mux_h
    port map (
            O => \N__34993\,
            I => \N__34825\
        );

    \I__7838\ : ClkMux
    port map (
            O => \N__34992\,
            I => \N__34822\
        );

    \I__7837\ : ClkMux
    port map (
            O => \N__34991\,
            I => \N__34816\
        );

    \I__7836\ : ClkMux
    port map (
            O => \N__34990\,
            I => \N__34813\
        );

    \I__7835\ : Span4Mux_v
    port map (
            O => \N__34987\,
            I => \N__34805\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__34982\,
            I => \N__34805\
        );

    \I__7833\ : Span4Mux_v
    port map (
            O => \N__34979\,
            I => \N__34805\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34976\,
            I => \N__34800\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__34973\,
            I => \N__34800\
        );

    \I__7830\ : Span4Mux_v
    port map (
            O => \N__34970\,
            I => \N__34793\
        );

    \I__7829\ : Span4Mux_s2_h
    port map (
            O => \N__34967\,
            I => \N__34793\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__34964\,
            I => \N__34793\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34790\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__34958\,
            I => \N__34787\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__34955\,
            I => \N__34778\
        );

    \I__7824\ : Span4Mux_v
    port map (
            O => \N__34952\,
            I => \N__34778\
        );

    \I__7823\ : Span4Mux_s3_h
    port map (
            O => \N__34949\,
            I => \N__34778\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__34946\,
            I => \N__34778\
        );

    \I__7821\ : ClkMux
    port map (
            O => \N__34945\,
            I => \N__34775\
        );

    \I__7820\ : Span4Mux_v
    port map (
            O => \N__34940\,
            I => \N__34772\
        );

    \I__7819\ : Span4Mux_v
    port map (
            O => \N__34935\,
            I => \N__34767\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__34932\,
            I => \N__34767\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__34929\,
            I => \N__34764\
        );

    \I__7816\ : Span4Mux_v
    port map (
            O => \N__34926\,
            I => \N__34761\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__34923\,
            I => \N__34752\
        );

    \I__7814\ : Span4Mux_h
    port map (
            O => \N__34920\,
            I => \N__34752\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__34917\,
            I => \N__34752\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__34914\,
            I => \N__34752\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__34911\,
            I => \N__34749\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34746\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__34905\,
            I => \N__34743\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__34902\,
            I => \N__34736\
        );

    \I__7807\ : Span4Mux_s2_h
    port map (
            O => \N__34899\,
            I => \N__34736\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__34896\,
            I => \N__34736\
        );

    \I__7805\ : ClkMux
    port map (
            O => \N__34895\,
            I => \N__34733\
        );

    \I__7804\ : Span4Mux_v
    port map (
            O => \N__34886\,
            I => \N__34728\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__34883\,
            I => \N__34728\
        );

    \I__7802\ : Span4Mux_v
    port map (
            O => \N__34876\,
            I => \N__34721\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__34873\,
            I => \N__34721\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__34870\,
            I => \N__34721\
        );

    \I__7799\ : Span4Mux_v
    port map (
            O => \N__34863\,
            I => \N__34710\
        );

    \I__7798\ : Span4Mux_h
    port map (
            O => \N__34860\,
            I => \N__34710\
        );

    \I__7797\ : Span4Mux_h
    port map (
            O => \N__34857\,
            I => \N__34710\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__34854\,
            I => \N__34710\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__34851\,
            I => \N__34710\
        );

    \I__7794\ : ClkMux
    port map (
            O => \N__34850\,
            I => \N__34707\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__34847\,
            I => \N__34704\
        );

    \I__7792\ : Span4Mux_v
    port map (
            O => \N__34842\,
            I => \N__34699\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34699\
        );

    \I__7790\ : Span4Mux_v
    port map (
            O => \N__34834\,
            I => \N__34694\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__34831\,
            I => \N__34694\
        );

    \I__7788\ : Span4Mux_s1_h
    port map (
            O => \N__34828\,
            I => \N__34691\
        );

    \I__7787\ : Span4Mux_v
    port map (
            O => \N__34825\,
            I => \N__34686\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__34822\,
            I => \N__34686\
        );

    \I__7785\ : ClkMux
    port map (
            O => \N__34821\,
            I => \N__34683\
        );

    \I__7784\ : ClkMux
    port map (
            O => \N__34820\,
            I => \N__34680\
        );

    \I__7783\ : ClkMux
    port map (
            O => \N__34819\,
            I => \N__34675\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34670\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__34813\,
            I => \N__34670\
        );

    \I__7780\ : ClkMux
    port map (
            O => \N__34812\,
            I => \N__34667\
        );

    \I__7779\ : Span4Mux_v
    port map (
            O => \N__34805\,
            I => \N__34660\
        );

    \I__7778\ : Span4Mux_v
    port map (
            O => \N__34800\,
            I => \N__34660\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__34793\,
            I => \N__34660\
        );

    \I__7776\ : Span4Mux_v
    port map (
            O => \N__34790\,
            I => \N__34655\
        );

    \I__7775\ : Span4Mux_s1_h
    port map (
            O => \N__34787\,
            I => \N__34655\
        );

    \I__7774\ : Span4Mux_v
    port map (
            O => \N__34778\,
            I => \N__34650\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__34775\,
            I => \N__34650\
        );

    \I__7772\ : Span4Mux_v
    port map (
            O => \N__34772\,
            I => \N__34639\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__34767\,
            I => \N__34639\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__34764\,
            I => \N__34639\
        );

    \I__7769\ : Span4Mux_h
    port map (
            O => \N__34761\,
            I => \N__34639\
        );

    \I__7768\ : Span4Mux_v
    port map (
            O => \N__34752\,
            I => \N__34639\
        );

    \I__7767\ : IoSpan4Mux
    port map (
            O => \N__34749\,
            I => \N__34636\
        );

    \I__7766\ : Span4Mux_v
    port map (
            O => \N__34746\,
            I => \N__34627\
        );

    \I__7765\ : Span4Mux_s2_h
    port map (
            O => \N__34743\,
            I => \N__34627\
        );

    \I__7764\ : Span4Mux_v
    port map (
            O => \N__34736\,
            I => \N__34627\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34627\
        );

    \I__7762\ : Span4Mux_h
    port map (
            O => \N__34728\,
            I => \N__34618\
        );

    \I__7761\ : IoSpan4Mux
    port map (
            O => \N__34721\,
            I => \N__34618\
        );

    \I__7760\ : Span4Mux_v
    port map (
            O => \N__34710\,
            I => \N__34618\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__34707\,
            I => \N__34618\
        );

    \I__7758\ : Span4Mux_s1_h
    port map (
            O => \N__34704\,
            I => \N__34613\
        );

    \I__7757\ : Span4Mux_s1_h
    port map (
            O => \N__34699\,
            I => \N__34613\
        );

    \I__7756\ : Span4Mux_v
    port map (
            O => \N__34694\,
            I => \N__34604\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__34691\,
            I => \N__34604\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__34686\,
            I => \N__34604\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__34683\,
            I => \N__34604\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34601\
        );

    \I__7751\ : ClkMux
    port map (
            O => \N__34679\,
            I => \N__34598\
        );

    \I__7750\ : ClkMux
    port map (
            O => \N__34678\,
            I => \N__34594\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__34675\,
            I => \N__34587\
        );

    \I__7748\ : Span4Mux_h
    port map (
            O => \N__34670\,
            I => \N__34587\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34587\
        );

    \I__7746\ : Span4Mux_v
    port map (
            O => \N__34660\,
            I => \N__34581\
        );

    \I__7745\ : Span4Mux_h
    port map (
            O => \N__34655\,
            I => \N__34581\
        );

    \I__7744\ : IoSpan4Mux
    port map (
            O => \N__34650\,
            I => \N__34576\
        );

    \I__7743\ : IoSpan4Mux
    port map (
            O => \N__34639\,
            I => \N__34576\
        );

    \I__7742\ : IoSpan4Mux
    port map (
            O => \N__34636\,
            I => \N__34569\
        );

    \I__7741\ : IoSpan4Mux
    port map (
            O => \N__34627\,
            I => \N__34569\
        );

    \I__7740\ : IoSpan4Mux
    port map (
            O => \N__34618\,
            I => \N__34569\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__34613\,
            I => \N__34560\
        );

    \I__7738\ : Span4Mux_v
    port map (
            O => \N__34604\,
            I => \N__34560\
        );

    \I__7737\ : Span4Mux_v
    port map (
            O => \N__34601\,
            I => \N__34560\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__34598\,
            I => \N__34560\
        );

    \I__7735\ : ClkMux
    port map (
            O => \N__34597\,
            I => \N__34557\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__34594\,
            I => \N__34552\
        );

    \I__7733\ : Sp12to4
    port map (
            O => \N__34587\,
            I => \N__34552\
        );

    \I__7732\ : ClkMux
    port map (
            O => \N__34586\,
            I => \N__34549\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__34581\,
            I => fpga_osc
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__34576\,
            I => fpga_osc
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__34569\,
            I => fpga_osc
        );

    \I__7728\ : Odrv4
    port map (
            O => \N__34560\,
            I => fpga_osc
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__34557\,
            I => fpga_osc
        );

    \I__7726\ : Odrv12
    port map (
            O => \N__34552\,
            I => fpga_osc
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__34549\,
            I => fpga_osc
        );

    \I__7724\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34498\
        );

    \I__7723\ : InMux
    port map (
            O => \N__34533\,
            I => \N__34498\
        );

    \I__7722\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34498\
        );

    \I__7721\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34498\
        );

    \I__7720\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34498\
        );

    \I__7719\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34491\
        );

    \I__7718\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34491\
        );

    \I__7717\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34491\
        );

    \I__7716\ : InMux
    port map (
            O => \N__34526\,
            I => \N__34480\
        );

    \I__7715\ : InMux
    port map (
            O => \N__34525\,
            I => \N__34480\
        );

    \I__7714\ : InMux
    port map (
            O => \N__34524\,
            I => \N__34480\
        );

    \I__7713\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34480\
        );

    \I__7712\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34480\
        );

    \I__7711\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34471\
        );

    \I__7710\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34471\
        );

    \I__7709\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34471\
        );

    \I__7708\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34471\
        );

    \I__7707\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34464\
        );

    \I__7706\ : InMux
    port map (
            O => \N__34516\,
            I => \N__34464\
        );

    \I__7705\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34464\
        );

    \I__7704\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34453\
        );

    \I__7703\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34453\
        );

    \I__7702\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34453\
        );

    \I__7701\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34453\
        );

    \I__7700\ : InMux
    port map (
            O => \N__34510\,
            I => \N__34453\
        );

    \I__7699\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34450\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__34498\,
            I => \N__34440\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__34491\,
            I => \N__34437\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__34480\,
            I => \N__34434\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__34471\,
            I => \N__34431\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__34464\,
            I => \N__34428\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__34453\,
            I => \N__34425\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__34450\,
            I => \N__34422\
        );

    \I__7691\ : CEMux
    port map (
            O => \N__34449\,
            I => \N__34393\
        );

    \I__7690\ : CEMux
    port map (
            O => \N__34448\,
            I => \N__34393\
        );

    \I__7689\ : CEMux
    port map (
            O => \N__34447\,
            I => \N__34393\
        );

    \I__7688\ : CEMux
    port map (
            O => \N__34446\,
            I => \N__34393\
        );

    \I__7687\ : CEMux
    port map (
            O => \N__34445\,
            I => \N__34393\
        );

    \I__7686\ : CEMux
    port map (
            O => \N__34444\,
            I => \N__34393\
        );

    \I__7685\ : CEMux
    port map (
            O => \N__34443\,
            I => \N__34393\
        );

    \I__7684\ : Glb2LocalMux
    port map (
            O => \N__34440\,
            I => \N__34393\
        );

    \I__7683\ : Glb2LocalMux
    port map (
            O => \N__34437\,
            I => \N__34393\
        );

    \I__7682\ : Glb2LocalMux
    port map (
            O => \N__34434\,
            I => \N__34393\
        );

    \I__7681\ : Glb2LocalMux
    port map (
            O => \N__34431\,
            I => \N__34393\
        );

    \I__7680\ : Glb2LocalMux
    port map (
            O => \N__34428\,
            I => \N__34393\
        );

    \I__7679\ : Glb2LocalMux
    port map (
            O => \N__34425\,
            I => \N__34393\
        );

    \I__7678\ : Glb2LocalMux
    port map (
            O => \N__34422\,
            I => \N__34393\
        );

    \I__7677\ : GlobalMux
    port map (
            O => \N__34393\,
            I => \N__34390\
        );

    \I__7676\ : gio2CtrlBuf
    port map (
            O => \N__34390\,
            I => \HDA_STRAP.count_en_g\
        );

    \I__7675\ : InMux
    port map (
            O => \N__34387\,
            I => \N__34384\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__34384\,
            I => \N__34380\
        );

    \I__7673\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34377\
        );

    \I__7672\ : Span4Mux_s3_h
    port map (
            O => \N__34380\,
            I => \N__34374\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__34377\,
            I => \N__34371\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__34374\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__7669\ : Odrv12
    port map (
            O => \N__34371\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__7668\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34363\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__34363\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__7666\ : InMux
    port map (
            O => \N__34360\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__7665\ : CascadeMux
    port map (
            O => \N__34357\,
            I => \N__34354\
        );

    \I__7664\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34351\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__34351\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__7662\ : InMux
    port map (
            O => \N__34348\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__7661\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34342\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__34342\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__7659\ : InMux
    port map (
            O => \N__34339\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__34336\,
            I => \N__34333\
        );

    \I__7657\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34330\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__34330\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__7655\ : InMux
    port map (
            O => \N__34327\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__7654\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34321\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__34321\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__7652\ : InMux
    port map (
            O => \N__34318\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__7651\ : InMux
    port map (
            O => \N__34315\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__7650\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34308\
        );

    \I__7649\ : CascadeMux
    port map (
            O => \N__34311\,
            I => \N__34305\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34299\
        );

    \I__7647\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34292\
        );

    \I__7646\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34292\
        );

    \I__7645\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34292\
        );

    \I__7644\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34289\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__34299\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__34292\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__34289\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__34282\,
            I => \N__34278\
        );

    \I__7639\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34270\
        );

    \I__7638\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34270\
        );

    \I__7637\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34270\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__34270\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__7635\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34263\
        );

    \I__7634\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34260\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__34263\,
            I => \N__34257\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__34260\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__7631\ : Odrv4
    port map (
            O => \N__34257\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__7630\ : InMux
    port map (
            O => \N__34252\,
            I => \HDA_STRAP.un2_count_1_cry_13\
        );

    \I__7629\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__34246\,
            I => \HDA_STRAP.un2_count_1_axb_15\
        );

    \I__7627\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34234\
        );

    \I__7626\ : InMux
    port map (
            O => \N__34242\,
            I => \N__34234\
        );

    \I__7625\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34234\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__34234\,
            I => \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0\
        );

    \I__7623\ : InMux
    port map (
            O => \N__34231\,
            I => \HDA_STRAP.un2_count_1_cry_14\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__34228\,
            I => \N__34225\
        );

    \I__7621\ : InMux
    port map (
            O => \N__34225\,
            I => \N__34222\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__34222\,
            I => \HDA_STRAP.un2_count_1_axb_16\
        );

    \I__7619\ : CascadeMux
    port map (
            O => \N__34219\,
            I => \N__34216\
        );

    \I__7618\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34211\
        );

    \I__7617\ : InMux
    port map (
            O => \N__34215\,
            I => \N__34206\
        );

    \I__7616\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34206\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__34211\,
            I => \HDA_STRAP.count_1_16\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__34206\,
            I => \HDA_STRAP.count_1_16\
        );

    \I__7613\ : InMux
    port map (
            O => \N__34201\,
            I => \HDA_STRAP.un2_count_1_cry_15\
        );

    \I__7612\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34189\
        );

    \I__7611\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34189\
        );

    \I__7610\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34189\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34182\
        );

    \I__7608\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34179\
        );

    \I__7607\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34176\
        );

    \I__7606\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34171\
        );

    \I__7605\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34171\
        );

    \I__7604\ : Span4Mux_s0_v
    port map (
            O => \N__34182\,
            I => \N__34168\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__34179\,
            I => \N__34161\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__34176\,
            I => \N__34161\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34161\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__34168\,
            I => \N__34155\
        );

    \I__7599\ : Span4Mux_v
    port map (
            O => \N__34161\,
            I => \N__34152\
        );

    \I__7598\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34147\
        );

    \I__7597\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34147\
        );

    \I__7596\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34144\
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__34155\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__7594\ : Odrv4
    port map (
            O => \N__34152\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__34147\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__34144\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__7591\ : InMux
    port map (
            O => \N__34135\,
            I => \bfn_12_7_0_\
        );

    \I__7590\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34129\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__34129\,
            I => \N__34125\
        );

    \I__7588\ : InMux
    port map (
            O => \N__34128\,
            I => \N__34122\
        );

    \I__7587\ : Span12Mux_s7_h
    port map (
            O => \N__34125\,
            I => \N__34119\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__34122\,
            I => \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\
        );

    \I__7585\ : Odrv12
    port map (
            O => \N__34119\,
            I => \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\
        );

    \I__7584\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__34111\,
            I => \N__34108\
        );

    \I__7582\ : Span4Mux_s3_h
    port map (
            O => \N__34108\,
            I => \N__34105\
        );

    \I__7581\ : Odrv4
    port map (
            O => \N__34105\,
            I => \HDA_STRAP.count_0_17\
        );

    \I__7580\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34098\
        );

    \I__7579\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34095\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__34098\,
            I => \N__34092\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__34095\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__34092\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__7575\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34083\
        );

    \I__7574\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34080\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__34075\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34075\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__34075\,
            I => \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\
        );

    \I__7570\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34069\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__34069\,
            I => \HDA_STRAP.count_1_4\
        );

    \I__7568\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34062\
        );

    \I__7567\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34059\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__34062\,
            I => \N__34054\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__34059\,
            I => \N__34054\
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__34054\,
            I => \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\
        );

    \I__7563\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34048\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__34048\,
            I => \HDA_STRAP.count_1_7\
        );

    \I__7561\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34042\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__34042\,
            I => \N__34038\
        );

    \I__7559\ : InMux
    port map (
            O => \N__34041\,
            I => \N__34035\
        );

    \I__7558\ : Odrv4
    port map (
            O => \N__34038\,
            I => \HDA_STRAP.count_1_10\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__34035\,
            I => \HDA_STRAP.count_1_10\
        );

    \I__7556\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34027\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__34024\
        );

    \I__7554\ : Odrv4
    port map (
            O => \N__34024\,
            I => \HDA_STRAP.count_1_0_10\
        );

    \I__7553\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34018\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__34018\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__7551\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34009\
        );

    \I__7550\ : InMux
    port map (
            O => \N__34014\,
            I => \N__34009\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__34009\,
            I => \HDA_STRAP.count_1_6\
        );

    \I__7548\ : InMux
    port map (
            O => \N__34006\,
            I => \HDA_STRAP.un2_count_1_cry_5_cZ0\
        );

    \I__7547\ : InMux
    port map (
            O => \N__34003\,
            I => \N__34000\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__34000\,
            I => \N__33996\
        );

    \I__7545\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33993\
        );

    \I__7544\ : Span4Mux_s0_h
    port map (
            O => \N__33996\,
            I => \N__33990\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__33993\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__33990\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__7541\ : InMux
    port map (
            O => \N__33985\,
            I => \HDA_STRAP.un2_count_1_cry_6\
        );

    \I__7540\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33979\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__33979\,
            I => \HDA_STRAP.un2_count_1_axb_8\
        );

    \I__7538\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33967\
        );

    \I__7537\ : InMux
    port map (
            O => \N__33975\,
            I => \N__33967\
        );

    \I__7536\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33967\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__33967\,
            I => \HDA_STRAP.count_1_8\
        );

    \I__7534\ : InMux
    port map (
            O => \N__33964\,
            I => \HDA_STRAP.un2_count_1_cry_7\
        );

    \I__7533\ : InMux
    port map (
            O => \N__33961\,
            I => \N__33958\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__33958\,
            I => \HDA_STRAP.un2_count_1_axb_9\
        );

    \I__7531\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33946\
        );

    \I__7530\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33946\
        );

    \I__7529\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33946\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__33946\,
            I => \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84\
        );

    \I__7527\ : InMux
    port map (
            O => \N__33943\,
            I => \bfn_12_6_0_\
        );

    \I__7526\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33936\
        );

    \I__7525\ : CascadeMux
    port map (
            O => \N__33939\,
            I => \N__33933\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__33936\,
            I => \N__33930\
        );

    \I__7523\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33927\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__33930\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__33927\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__7520\ : InMux
    port map (
            O => \N__33922\,
            I => \HDA_STRAP.un2_count_1_cry_9\
        );

    \I__7519\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33915\
        );

    \I__7518\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33912\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__33915\,
            I => \N__33907\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__33912\,
            I => \N__33907\
        );

    \I__7515\ : Odrv4
    port map (
            O => \N__33907\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__7514\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33898\
        );

    \I__7513\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33898\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33895\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__33895\,
            I => \HDA_STRAP.count_1_11\
        );

    \I__7510\ : InMux
    port map (
            O => \N__33892\,
            I => \HDA_STRAP.un2_count_1_cry_10\
        );

    \I__7509\ : InMux
    port map (
            O => \N__33889\,
            I => \N__33886\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__33886\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__7507\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__7506\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33877\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__33877\,
            I => \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3\
        );

    \I__7504\ : InMux
    port map (
            O => \N__33874\,
            I => \HDA_STRAP.un2_count_1_cry_11\
        );

    \I__7503\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33868\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__33868\,
            I => \HDA_STRAP.un2_count_1_axb_13\
        );

    \I__7501\ : InMux
    port map (
            O => \N__33865\,
            I => \N__33856\
        );

    \I__7500\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33856\
        );

    \I__7499\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33856\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__33856\,
            I => \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\
        );

    \I__7497\ : InMux
    port map (
            O => \N__33853\,
            I => \HDA_STRAP.un2_count_1_cry_12\
        );

    \I__7496\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33847\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__33847\,
            I => \HDA_STRAP.count_1_2\
        );

    \I__7494\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33841\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__33841\,
            I => \HDA_STRAP.count_1_0_11\
        );

    \I__7492\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33829\
        );

    \I__7491\ : InMux
    port map (
            O => \N__33837\,
            I => \N__33829\
        );

    \I__7490\ : InMux
    port map (
            O => \N__33836\,
            I => \N__33826\
        );

    \I__7489\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33821\
        );

    \I__7488\ : InMux
    port map (
            O => \N__33834\,
            I => \N__33821\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__33829\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__33826\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__33821\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__7484\ : CascadeMux
    port map (
            O => \N__33814\,
            I => \N__33811\
        );

    \I__7483\ : InMux
    port map (
            O => \N__33811\,
            I => \N__33807\
        );

    \I__7482\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33804\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__33807\,
            I => \N__33801\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__33804\,
            I => \HDA_STRAP.un2_count_1_axb_1\
        );

    \I__7479\ : Odrv4
    port map (
            O => \N__33801\,
            I => \HDA_STRAP.un2_count_1_axb_1\
        );

    \I__7478\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33793\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__33793\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__33790\,
            I => \N__33786\
        );

    \I__7475\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33781\
        );

    \I__7474\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33781\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__33781\,
            I => \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614\
        );

    \I__7472\ : InMux
    port map (
            O => \N__33778\,
            I => \HDA_STRAP.un2_count_1_cry_1\
        );

    \I__7471\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33772\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__33772\,
            I => \N__33769\
        );

    \I__7469\ : Odrv4
    port map (
            O => \N__33769\,
            I => \HDA_STRAP.un2_count_1_axb_3\
        );

    \I__7468\ : CascadeMux
    port map (
            O => \N__33766\,
            I => \N__33762\
        );

    \I__7467\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33754\
        );

    \I__7466\ : InMux
    port map (
            O => \N__33762\,
            I => \N__33754\
        );

    \I__7465\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33754\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__33754\,
            I => \N__33751\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__33751\,
            I => \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824\
        );

    \I__7462\ : InMux
    port map (
            O => \N__33748\,
            I => \HDA_STRAP.un2_count_1_cry_2\
        );

    \I__7461\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33741\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33738\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33735\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__33738\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__33735\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__7456\ : InMux
    port map (
            O => \N__33730\,
            I => \HDA_STRAP.un2_count_1_cry_3\
        );

    \I__7455\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33724\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__33724\,
            I => \HDA_STRAP.un2_count_1_axb_5\
        );

    \I__7453\ : InMux
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__33718\,
            I => \N__33713\
        );

    \I__7451\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33708\
        );

    \I__7450\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33708\
        );

    \I__7449\ : Odrv4
    port map (
            O => \N__33713\,
            I => \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__33708\,
            I => \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\
        );

    \I__7447\ : InMux
    port map (
            O => \N__33703\,
            I => \HDA_STRAP.un2_count_1_cry_4\
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__33700\,
            I => \VPP_VDDQ.count_2_rst_7_cascade_\
        );

    \I__7445\ : InMux
    port map (
            O => \N__33697\,
            I => \N__33692\
        );

    \I__7444\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33687\
        );

    \I__7443\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33687\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__33692\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__33687\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__7440\ : CascadeMux
    port map (
            O => \N__33682\,
            I => \N__33676\
        );

    \I__7439\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33672\
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__33680\,
            I => \N__33669\
        );

    \I__7437\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33666\
        );

    \I__7436\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33661\
        );

    \I__7435\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33661\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33658\
        );

    \I__7433\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33655\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__33666\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__33661\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__33658\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__33655\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7428\ : CascadeMux
    port map (
            O => \N__33646\,
            I => \VPP_VDDQ.count_2Z0Z_1_cascade_\
        );

    \I__7427\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33640\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__33640\,
            I => \VPP_VDDQ.count_2_0_1\
        );

    \I__7425\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33633\
        );

    \I__7424\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33630\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__33633\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__33630\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__7421\ : CascadeMux
    port map (
            O => \N__33625\,
            I => \N__33622\
        );

    \I__7420\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33619\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__33619\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__7418\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33610\
        );

    \I__7417\ : SRMux
    port map (
            O => \N__33615\,
            I => \N__33610\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__7415\ : Span4Mux_s1_v
    port map (
            O => \N__33607\,
            I => \N__33596\
        );

    \I__7414\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33593\
        );

    \I__7413\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33586\
        );

    \I__7412\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33586\
        );

    \I__7411\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33586\
        );

    \I__7410\ : SRMux
    port map (
            O => \N__33602\,
            I => \N__33583\
        );

    \I__7409\ : SRMux
    port map (
            O => \N__33601\,
            I => \N__33580\
        );

    \I__7408\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33564\
        );

    \I__7407\ : SRMux
    port map (
            O => \N__33599\,
            I => \N__33564\
        );

    \I__7406\ : IoSpan4Mux
    port map (
            O => \N__33596\,
            I => \N__33552\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__33593\,
            I => \N__33552\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33552\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__33583\,
            I => \N__33544\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33541\
        );

    \I__7401\ : SRMux
    port map (
            O => \N__33579\,
            I => \N__33538\
        );

    \I__7400\ : InMux
    port map (
            O => \N__33578\,
            I => \N__33531\
        );

    \I__7399\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33531\
        );

    \I__7398\ : SRMux
    port map (
            O => \N__33576\,
            I => \N__33531\
        );

    \I__7397\ : InMux
    port map (
            O => \N__33575\,
            I => \N__33528\
        );

    \I__7396\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33517\
        );

    \I__7395\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33517\
        );

    \I__7394\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33517\
        );

    \I__7393\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33517\
        );

    \I__7392\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33512\
        );

    \I__7391\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33512\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__33564\,
            I => \N__33509\
        );

    \I__7389\ : InMux
    port map (
            O => \N__33563\,
            I => \N__33498\
        );

    \I__7388\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33498\
        );

    \I__7387\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33498\
        );

    \I__7386\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33498\
        );

    \I__7385\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33498\
        );

    \I__7384\ : IoSpan4Mux
    port map (
            O => \N__33552\,
            I => \N__33495\
        );

    \I__7383\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33492\
        );

    \I__7382\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33485\
        );

    \I__7381\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33485\
        );

    \I__7380\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33485\
        );

    \I__7379\ : SRMux
    port map (
            O => \N__33547\,
            I => \N__33482\
        );

    \I__7378\ : Span4Mux_v
    port map (
            O => \N__33544\,
            I => \N__33477\
        );

    \I__7377\ : Span4Mux_s2_h
    port map (
            O => \N__33541\,
            I => \N__33477\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__33538\,
            I => \N__33472\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__33531\,
            I => \N__33472\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33469\
        );

    \I__7373\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33464\
        );

    \I__7372\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33464\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__33517\,
            I => \N__33459\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__33512\,
            I => \N__33459\
        );

    \I__7369\ : Span4Mux_s1_h
    port map (
            O => \N__33509\,
            I => \N__33452\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__33498\,
            I => \N__33452\
        );

    \I__7367\ : IoSpan4Mux
    port map (
            O => \N__33495\,
            I => \N__33452\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__33492\,
            I => \N__33447\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33447\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__33482\,
            I => \N__33444\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__33477\,
            I => \N__33441\
        );

    \I__7362\ : Span4Mux_s3_v
    port map (
            O => \N__33472\,
            I => \N__33434\
        );

    \I__7361\ : Span4Mux_v
    port map (
            O => \N__33469\,
            I => \N__33434\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__33464\,
            I => \N__33434\
        );

    \I__7359\ : Span4Mux_s2_v
    port map (
            O => \N__33459\,
            I => \N__33427\
        );

    \I__7358\ : Span4Mux_s2_v
    port map (
            O => \N__33452\,
            I => \N__33427\
        );

    \I__7357\ : Span4Mux_s1_h
    port map (
            O => \N__33447\,
            I => \N__33427\
        );

    \I__7356\ : Span12Mux_s6_v
    port map (
            O => \N__33444\,
            I => \N__33424\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__33441\,
            I => \N__33421\
        );

    \I__7354\ : Span4Mux_h
    port map (
            O => \N__33434\,
            I => \N__33418\
        );

    \I__7353\ : Span4Mux_h
    port map (
            O => \N__33427\,
            I => \N__33415\
        );

    \I__7352\ : Odrv12
    port map (
            O => \N__33424\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__33421\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__7350\ : Odrv4
    port map (
            O => \N__33418\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__7349\ : Odrv4
    port map (
            O => \N__33415\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__7348\ : CEMux
    port map (
            O => \N__33406\,
            I => \N__33400\
        );

    \I__7347\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33395\
        );

    \I__7346\ : CEMux
    port map (
            O => \N__33404\,
            I => \N__33395\
        );

    \I__7345\ : CEMux
    port map (
            O => \N__33403\,
            I => \N__33392\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__33400\,
            I => \N__33373\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__33395\,
            I => \N__33373\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__33392\,
            I => \N__33373\
        );

    \I__7341\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33368\
        );

    \I__7340\ : CEMux
    port map (
            O => \N__33390\,
            I => \N__33368\
        );

    \I__7339\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33363\
        );

    \I__7338\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33363\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__33387\,
            I => \N__33356\
        );

    \I__7336\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33350\
        );

    \I__7335\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33350\
        );

    \I__7334\ : CEMux
    port map (
            O => \N__33384\,
            I => \N__33347\
        );

    \I__7333\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33344\
        );

    \I__7332\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33337\
        );

    \I__7331\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33337\
        );

    \I__7330\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33337\
        );

    \I__7329\ : Sp12to4
    port map (
            O => \N__33373\,
            I => \N__33334\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33322\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__33363\,
            I => \N__33322\
        );

    \I__7326\ : CEMux
    port map (
            O => \N__33362\,
            I => \N__33319\
        );

    \I__7325\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33312\
        );

    \I__7324\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33312\
        );

    \I__7323\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33312\
        );

    \I__7322\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33307\
        );

    \I__7321\ : CEMux
    port map (
            O => \N__33355\,
            I => \N__33307\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33304\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__33347\,
            I => \N__33301\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__33344\,
            I => \N__33296\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__33337\,
            I => \N__33296\
        );

    \I__7316\ : Span12Mux_s3_v
    port map (
            O => \N__33334\,
            I => \N__33293\
        );

    \I__7315\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33282\
        );

    \I__7314\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33282\
        );

    \I__7313\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33282\
        );

    \I__7312\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33282\
        );

    \I__7311\ : InMux
    port map (
            O => \N__33329\,
            I => \N__33282\
        );

    \I__7310\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33279\
        );

    \I__7309\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33276\
        );

    \I__7308\ : Span4Mux_s2_h
    port map (
            O => \N__33322\,
            I => \N__33273\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33268\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__33312\,
            I => \N__33268\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__33307\,
            I => \N__33263\
        );

    \I__7304\ : Span4Mux_s3_v
    port map (
            O => \N__33304\,
            I => \N__33263\
        );

    \I__7303\ : Span4Mux_h
    port map (
            O => \N__33301\,
            I => \N__33258\
        );

    \I__7302\ : Span4Mux_s2_h
    port map (
            O => \N__33296\,
            I => \N__33258\
        );

    \I__7301\ : Odrv12
    port map (
            O => \N__33293\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__33282\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__33279\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__33276\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__33273\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__33268\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__33263\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7294\ : Odrv4
    port map (
            O => \N__33258\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__7293\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33238\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__7291\ : Odrv4
    port map (
            O => \N__33235\,
            I => \VPP_VDDQ.count_2_0_4\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__33232\,
            I => \N__33228\
        );

    \I__7289\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33225\
        );

    \I__7288\ : InMux
    port map (
            O => \N__33228\,
            I => \N__33222\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__33225\,
            I => \VPP_VDDQ.count_2_rst_4\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__33222\,
            I => \VPP_VDDQ.count_2_rst_4\
        );

    \I__7285\ : InMux
    port map (
            O => \N__33217\,
            I => \N__33213\
        );

    \I__7284\ : InMux
    port map (
            O => \N__33216\,
            I => \N__33210\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__33213\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__33210\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__33205\,
            I => \HDA_STRAP.countZ0Z_2_cascade_\
        );

    \I__7280\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33199\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__33199\,
            I => \HDA_STRAP.un25_clk_100khz_1\
        );

    \I__7278\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33193\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__33193\,
            I => \HDA_STRAP.count_RNIZ0Z_1\
        );

    \I__7276\ : CascadeMux
    port map (
            O => \N__33190\,
            I => \HDA_STRAP.count_RNIZ0Z_1_cascade_\
        );

    \I__7275\ : CascadeMux
    port map (
            O => \N__33187\,
            I => \HDA_STRAP.un2_count_1_axb_1_cascade_\
        );

    \I__7274\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33178\
        );

    \I__7273\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33178\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__33178\,
            I => \HDA_STRAP.count_1_1\
        );

    \I__7271\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33172\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__33172\,
            I => \VPP_VDDQ.un29_clk_100khz_4\
        );

    \I__7269\ : InMux
    port map (
            O => \N__33169\,
            I => \N__33166\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__33166\,
            I => \N__33163\
        );

    \I__7267\ : Span4Mux_s2_v
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__33160\,
            I => \VPP_VDDQ.un29_clk_100khz_12\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__33157\,
            I => \VPP_VDDQ.un29_clk_100khz_5_cascade_\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__33154\,
            I => \VPP_VDDQ.N_1_i_cascade_\
        );

    \I__7263\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__33148\,
            I => \VPP_VDDQ.count_2_rst_3\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__33145\,
            I => \VPP_VDDQ.count_2_rst_3_cascade_\
        );

    \I__7260\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33138\
        );

    \I__7259\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33135\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__33138\,
            I => \VPP_VDDQ.un1_count_2_1_axb_5\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__33135\,
            I => \VPP_VDDQ.un1_count_2_1_axb_5\
        );

    \I__7256\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__7255\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33124\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__33124\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__33121\,
            I => \VPP_VDDQ.un1_count_2_1_axb_5_cascade_\
        );

    \I__7252\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33112\
        );

    \I__7251\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33112\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__33112\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__7249\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33106\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__33106\,
            I => \N__33103\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__33103\,
            I => \N__33099\
        );

    \I__7246\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33096\
        );

    \I__7245\ : Sp12to4
    port map (
            O => \N__33099\,
            I => \N__33093\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__33096\,
            I => \N__33090\
        );

    \I__7243\ : Odrv12
    port map (
            O => \N__33093\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__33090\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__7241\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33082\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__33082\,
            I => \VPP_VDDQ.un29_clk_100khz_11\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__33079\,
            I => \N__33076\
        );

    \I__7238\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33067\
        );

    \I__7237\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33067\
        );

    \I__7236\ : InMux
    port map (
            O => \N__33074\,
            I => \N__33067\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__33067\,
            I => \N__33061\
        );

    \I__7234\ : CascadeMux
    port map (
            O => \N__33066\,
            I => \N__33057\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__33065\,
            I => \N__33050\
        );

    \I__7232\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33046\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__33061\,
            I => \N__33043\
        );

    \I__7230\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33040\
        );

    \I__7229\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33037\
        );

    \I__7228\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33032\
        );

    \I__7227\ : InMux
    port map (
            O => \N__33055\,
            I => \N__33032\
        );

    \I__7226\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33023\
        );

    \I__7225\ : InMux
    port map (
            O => \N__33053\,
            I => \N__33023\
        );

    \I__7224\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33023\
        );

    \I__7223\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33023\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__33046\,
            I => \N__33018\
        );

    \I__7221\ : Span4Mux_h
    port map (
            O => \N__33043\,
            I => \N__33018\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__33040\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__33037\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__33032\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__33023\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__33018\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7215\ : InMux
    port map (
            O => \N__33007\,
            I => \N__33004\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__33004\,
            I => \N__33001\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__33001\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__32998\,
            I => \VPP_VDDQ.count_2_rst_8_cascade_\
        );

    \I__7211\ : CascadeMux
    port map (
            O => \N__32995\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__7210\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32986\
        );

    \I__7209\ : InMux
    port map (
            O => \N__32991\,
            I => \N__32986\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__32986\,
            I => \N__32983\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__32983\,
            I => \POWERLED.dutycycle_en_10\
        );

    \I__7206\ : InMux
    port map (
            O => \N__32980\,
            I => \N__32974\
        );

    \I__7205\ : InMux
    port map (
            O => \N__32979\,
            I => \N__32974\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__7203\ : Odrv12
    port map (
            O => \N__32971\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__32968\,
            I => \N__32964\
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \N__32961\
        );

    \I__7200\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32956\
        );

    \I__7199\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32956\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__32956\,
            I => \POWERLED.dutycycleZ1Z_13\
        );

    \I__7197\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32948\
        );

    \I__7196\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32945\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__32951\,
            I => \N__32934\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32948\,
            I => \N__32927\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32927\
        );

    \I__7192\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32920\
        );

    \I__7191\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32920\
        );

    \I__7190\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32920\
        );

    \I__7189\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32915\
        );

    \I__7188\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32912\
        );

    \I__7187\ : CascadeMux
    port map (
            O => \N__32939\,
            I => \N__32905\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__32938\,
            I => \N__32902\
        );

    \I__7185\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32898\
        );

    \I__7184\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32886\
        );

    \I__7183\ : InMux
    port map (
            O => \N__32933\,
            I => \N__32881\
        );

    \I__7182\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32881\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__32927\,
            I => \N__32876\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32876\
        );

    \I__7179\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32873\
        );

    \I__7178\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32868\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__32915\,
            I => \N__32865\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32862\
        );

    \I__7175\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32855\
        );

    \I__7174\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32855\
        );

    \I__7173\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32855\
        );

    \I__7172\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32850\
        );

    \I__7171\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32843\
        );

    \I__7170\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32843\
        );

    \I__7169\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32843\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__32898\,
            I => \N__32840\
        );

    \I__7167\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32837\
        );

    \I__7166\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32828\
        );

    \I__7165\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32828\
        );

    \I__7164\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32828\
        );

    \I__7163\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32828\
        );

    \I__7162\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32819\
        );

    \I__7161\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32819\
        );

    \I__7160\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32819\
        );

    \I__7159\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32819\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32814\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32814\
        );

    \I__7156\ : Span4Mux_v
    port map (
            O => \N__32876\,
            I => \N__32809\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__32873\,
            I => \N__32809\
        );

    \I__7154\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32804\
        );

    \I__7153\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32804\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__32868\,
            I => \N__32801\
        );

    \I__7151\ : Span4Mux_s3_v
    port map (
            O => \N__32865\,
            I => \N__32798\
        );

    \I__7150\ : Span4Mux_s3_v
    port map (
            O => \N__32862\,
            I => \N__32793\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__32855\,
            I => \N__32793\
        );

    \I__7148\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32788\
        );

    \I__7147\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32788\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__32850\,
            I => \N__32783\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32783\
        );

    \I__7144\ : Span4Mux_h
    port map (
            O => \N__32840\,
            I => \N__32780\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32767\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32767\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32767\
        );

    \I__7140\ : Span4Mux_h
    port map (
            O => \N__32814\,
            I => \N__32767\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__32809\,
            I => \N__32767\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32767\
        );

    \I__7137\ : Odrv12
    port map (
            O => \N__32801\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__32798\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__32793\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__32788\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__32783\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__32780\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__32767\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1\
        );

    \I__7130\ : CascadeMux
    port map (
            O => \N__32752\,
            I => \N__32745\
        );

    \I__7129\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32742\
        );

    \I__7128\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32739\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__32749\,
            I => \N__32736\
        );

    \I__7126\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32733\
        );

    \I__7125\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32730\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__32742\,
            I => \N__32725\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__32739\,
            I => \N__32725\
        );

    \I__7122\ : InMux
    port map (
            O => \N__32736\,
            I => \N__32721\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__32733\,
            I => \N__32718\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__32730\,
            I => \N__32713\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__32725\,
            I => \N__32713\
        );

    \I__7118\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32708\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__32721\,
            I => \N__32705\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__32718\,
            I => \N__32702\
        );

    \I__7115\ : IoSpan4Mux
    port map (
            O => \N__32713\,
            I => \N__32699\
        );

    \I__7114\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32694\
        );

    \I__7113\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32694\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32689\
        );

    \I__7111\ : Span4Mux_h
    port map (
            O => \N__32705\,
            I => \N__32689\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__32702\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__32699\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__32694\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__32689\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__32680\,
            I => \N__32674\
        );

    \I__7105\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32668\
        );

    \I__7104\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32665\
        );

    \I__7103\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32660\
        );

    \I__7102\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32660\
        );

    \I__7101\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32657\
        );

    \I__7100\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32652\
        );

    \I__7099\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32652\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32644\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__32665\,
            I => \N__32644\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32644\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__32657\,
            I => \N__32641\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__32652\,
            I => \N__32638\
        );

    \I__7093\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32635\
        );

    \I__7092\ : Span4Mux_s3_h
    port map (
            O => \N__32644\,
            I => \N__32632\
        );

    \I__7091\ : Span12Mux_s7_h
    port map (
            O => \N__32641\,
            I => \N__32629\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__32638\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__32635\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__32632\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__7087\ : Odrv12
    port map (
            O => \N__32629\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__32620\,
            I => \POWERLED.dutycycleZ0Z_10_cascade_\
        );

    \I__7085\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32614\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__32614\,
            I => \POWERLED.un1_dutycycle_53_2_1_0_tz\
        );

    \I__7083\ : CascadeMux
    port map (
            O => \N__32611\,
            I => \POWERLED.un1_dutycycle_53_3_1_cascade_\
        );

    \I__7082\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32604\
        );

    \I__7081\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32601\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32596\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__32601\,
            I => \N__32596\
        );

    \I__7078\ : Span4Mux_h
    port map (
            O => \N__32596\,
            I => \N__32593\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__32593\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_9\
        );

    \I__7076\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32586\
        );

    \I__7075\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32583\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__32586\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__32583\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\
        );

    \I__7072\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32575\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__32575\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__32572\,
            I => \VPP_VDDQ.count_2_rst_0_cascade_\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__32569\,
            I => \N__32565\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \N__32561\
        );

    \I__7067\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32558\
        );

    \I__7066\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32555\
        );

    \I__7065\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32552\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__32558\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__32555\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__32552\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__32545\,
            I => \VPP_VDDQ.count_2Z0Z_8_cascade_\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__32542\,
            I => \N__32538\
        );

    \I__7059\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32532\
        );

    \I__7058\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32532\
        );

    \I__7057\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32528\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32525\
        );

    \I__7055\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32522\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__32528\,
            I => \N__32519\
        );

    \I__7053\ : Span4Mux_h
    port map (
            O => \N__32525\,
            I => \N__32514\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__32522\,
            I => \N__32514\
        );

    \I__7051\ : Span4Mux_s2_h
    port map (
            O => \N__32519\,
            I => \N__32511\
        );

    \I__7050\ : Span4Mux_s2_h
    port map (
            O => \N__32514\,
            I => \N__32508\
        );

    \I__7049\ : Odrv4
    port map (
            O => \N__32511\,
            I => \POWERLED.func_state_RNI_6Z0Z_0\
        );

    \I__7048\ : Odrv4
    port map (
            O => \N__32508\,
            I => \POWERLED.func_state_RNI_6Z0Z_0\
        );

    \I__7047\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32500\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__32500\,
            I => \N__32497\
        );

    \I__7045\ : Odrv12
    port map (
            O => \N__32497\,
            I => \POWERLED.un1_clk_100khz_40_and_i_0_d_0\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__32494\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_9_cascade_\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__32491\,
            I => \N__32488\
        );

    \I__7042\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32485\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__32485\,
            I => \N__32482\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__32482\,
            I => \N__32479\
        );

    \I__7039\ : Odrv4
    port map (
            O => \N__32479\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__7038\ : SRMux
    port map (
            O => \N__32476\,
            I => \N__32473\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32463\
        );

    \I__7036\ : SRMux
    port map (
            O => \N__32472\,
            I => \N__32460\
        );

    \I__7035\ : SRMux
    port map (
            O => \N__32471\,
            I => \N__32456\
        );

    \I__7034\ : SRMux
    port map (
            O => \N__32470\,
            I => \N__32453\
        );

    \I__7033\ : SRMux
    port map (
            O => \N__32469\,
            I => \N__32450\
        );

    \I__7032\ : SRMux
    port map (
            O => \N__32468\,
            I => \N__32447\
        );

    \I__7031\ : SRMux
    port map (
            O => \N__32467\,
            I => \N__32444\
        );

    \I__7030\ : SRMux
    port map (
            O => \N__32466\,
            I => \N__32441\
        );

    \I__7029\ : Span4Mux_s2_v
    port map (
            O => \N__32463\,
            I => \N__32435\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__32460\,
            I => \N__32435\
        );

    \I__7027\ : SRMux
    port map (
            O => \N__32459\,
            I => \N__32432\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__32456\,
            I => \N__32428\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__32453\,
            I => \N__32425\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__32450\,
            I => \N__32422\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32418\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__32444\,
            I => \N__32413\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__32441\,
            I => \N__32413\
        );

    \I__7020\ : SRMux
    port map (
            O => \N__32440\,
            I => \N__32410\
        );

    \I__7019\ : Span4Mux_v
    port map (
            O => \N__32435\,
            I => \N__32405\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__32432\,
            I => \N__32405\
        );

    \I__7017\ : SRMux
    port map (
            O => \N__32431\,
            I => \N__32402\
        );

    \I__7016\ : Span4Mux_s1_v
    port map (
            O => \N__32428\,
            I => \N__32397\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__32425\,
            I => \N__32397\
        );

    \I__7014\ : Span4Mux_s1_v
    port map (
            O => \N__32422\,
            I => \N__32394\
        );

    \I__7013\ : SRMux
    port map (
            O => \N__32421\,
            I => \N__32391\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__32418\,
            I => \N__32387\
        );

    \I__7011\ : Span4Mux_s1_v
    port map (
            O => \N__32413\,
            I => \N__32384\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__32410\,
            I => \N__32381\
        );

    \I__7009\ : Span4Mux_h
    port map (
            O => \N__32405\,
            I => \N__32378\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__32402\,
            I => \N__32375\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__32397\,
            I => \N__32370\
        );

    \I__7006\ : Span4Mux_v
    port map (
            O => \N__32394\,
            I => \N__32370\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__32391\,
            I => \N__32367\
        );

    \I__7004\ : SRMux
    port map (
            O => \N__32390\,
            I => \N__32364\
        );

    \I__7003\ : Span4Mux_h
    port map (
            O => \N__32387\,
            I => \N__32361\
        );

    \I__7002\ : Span4Mux_v
    port map (
            O => \N__32384\,
            I => \N__32358\
        );

    \I__7001\ : Span4Mux_s2_v
    port map (
            O => \N__32381\,
            I => \N__32353\
        );

    \I__7000\ : Span4Mux_s2_v
    port map (
            O => \N__32378\,
            I => \N__32353\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__32375\,
            I => \N__32348\
        );

    \I__6998\ : Span4Mux_h
    port map (
            O => \N__32370\,
            I => \N__32348\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__32367\,
            I => \POWERLED.func_m1_0_a2_0_isoZ0\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__32364\,
            I => \POWERLED.func_m1_0_a2_0_isoZ0\
        );

    \I__6995\ : Odrv4
    port map (
            O => \N__32361\,
            I => \POWERLED.func_m1_0_a2_0_isoZ0\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__32358\,
            I => \POWERLED.func_m1_0_a2_0_isoZ0\
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__32353\,
            I => \POWERLED.func_m1_0_a2_0_isoZ0\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__32348\,
            I => \POWERLED.func_m1_0_a2_0_isoZ0\
        );

    \I__6991\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32332\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__32332\,
            I => \N__32329\
        );

    \I__6989\ : Odrv12
    port map (
            O => \N__32329\,
            I => \POWERLED.un1_dutycycle_53_axb_14_1\
        );

    \I__6988\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32316\
        );

    \I__6987\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32313\
        );

    \I__6986\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32309\
        );

    \I__6985\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32306\
        );

    \I__6984\ : InMux
    port map (
            O => \N__32322\,
            I => \N__32303\
        );

    \I__6983\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32298\
        );

    \I__6982\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32298\
        );

    \I__6981\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32295\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__32316\,
            I => \N__32290\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__32313\,
            I => \N__32290\
        );

    \I__6978\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32287\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32284\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32281\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__32303\,
            I => \N__32278\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__32298\,
            I => \N__32275\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__32295\,
            I => \N__32270\
        );

    \I__6972\ : Span4Mux_h
    port map (
            O => \N__32290\,
            I => \N__32270\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__32287\,
            I => \N__32265\
        );

    \I__6970\ : Span4Mux_s2_v
    port map (
            O => \N__32284\,
            I => \N__32265\
        );

    \I__6969\ : Span4Mux_s1_v
    port map (
            O => \N__32281\,
            I => \N__32262\
        );

    \I__6968\ : Span4Mux_s2_v
    port map (
            O => \N__32278\,
            I => \N__32257\
        );

    \I__6967\ : Span4Mux_s2_v
    port map (
            O => \N__32275\,
            I => \N__32257\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__32270\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__32265\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__6964\ : Odrv4
    port map (
            O => \N__32262\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__32257\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__6962\ : CascadeMux
    port map (
            O => \N__32248\,
            I => \N__32245\
        );

    \I__6961\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32242\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32239\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__32239\,
            I => \N__32236\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__32236\,
            I => \POWERLED.un2_count_clk_17_0_a2_1_4\
        );

    \I__6957\ : CascadeMux
    port map (
            O => \N__32233\,
            I => \POWERLED.un1_dutycycle_53_4_a1_0_cascade_\
        );

    \I__6956\ : CascadeMux
    port map (
            O => \N__32230\,
            I => \N__32227\
        );

    \I__6955\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32224\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32221\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__32221\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__32218\,
            I => \POWERLED.un1_dutycycle_53_9_4_cascade_\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__32215\,
            I => \N__32212\
        );

    \I__6950\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32209\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32206\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__32206\,
            I => \N__32203\
        );

    \I__6947\ : Odrv4
    port map (
            O => \N__32203\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_11\
        );

    \I__6946\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32197\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__32197\,
            I => \POWERLED.g0_0_1\
        );

    \I__6944\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32191\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32188\
        );

    \I__6942\ : Span4Mux_s2_v
    port map (
            O => \N__32188\,
            I => \N__32185\
        );

    \I__6941\ : Span4Mux_h
    port map (
            O => \N__32185\,
            I => \N__32182\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__32182\,
            I => \POWERLED.un1_dutycycle_53_4_a3_0\
        );

    \I__6939\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32173\
        );

    \I__6938\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32169\
        );

    \I__6937\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32164\
        );

    \I__6936\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32164\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__32173\,
            I => \N__32160\
        );

    \I__6934\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32157\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__32169\,
            I => \N__32152\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32152\
        );

    \I__6931\ : CascadeMux
    port map (
            O => \N__32163\,
            I => \N__32149\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__32160\,
            I => \N__32146\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__32157\,
            I => \N__32141\
        );

    \I__6928\ : Span12Mux_v
    port map (
            O => \N__32152\,
            I => \N__32141\
        );

    \I__6927\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32138\
        );

    \I__6926\ : Odrv4
    port map (
            O => \N__32146\,
            I => \POWERLED.N_371\
        );

    \I__6925\ : Odrv12
    port map (
            O => \N__32141\,
            I => \POWERLED.N_371\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__32138\,
            I => \POWERLED.N_371\
        );

    \I__6923\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32127\
        );

    \I__6922\ : CascadeMux
    port map (
            O => \N__32130\,
            I => \N__32124\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__32127\,
            I => \N__32116\
        );

    \I__6920\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32113\
        );

    \I__6919\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32110\
        );

    \I__6918\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32106\
        );

    \I__6917\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32101\
        );

    \I__6916\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32101\
        );

    \I__6915\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32098\
        );

    \I__6914\ : Span4Mux_v
    port map (
            O => \N__32116\,
            I => \N__32094\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32089\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32089\
        );

    \I__6911\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32086\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__32083\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__32101\,
            I => \N__32080\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__32098\,
            I => \N__32075\
        );

    \I__6907\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32069\
        );

    \I__6906\ : Span4Mux_v
    port map (
            O => \N__32094\,
            I => \N__32060\
        );

    \I__6905\ : Span4Mux_s3_h
    port map (
            O => \N__32089\,
            I => \N__32060\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32060\
        );

    \I__6903\ : Span4Mux_v
    port map (
            O => \N__32083\,
            I => \N__32055\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__32080\,
            I => \N__32055\
        );

    \I__6901\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32050\
        );

    \I__6900\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32050\
        );

    \I__6899\ : Span4Mux_h
    port map (
            O => \N__32075\,
            I => \N__32047\
        );

    \I__6898\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32040\
        );

    \I__6897\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32040\
        );

    \I__6896\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32040\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32037\
        );

    \I__6894\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32034\
        );

    \I__6893\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32031\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__32060\,
            I => \N__32028\
        );

    \I__6891\ : Sp12to4
    port map (
            O => \N__32055\,
            I => \N__32023\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__32023\
        );

    \I__6889\ : Span4Mux_v
    port map (
            O => \N__32047\,
            I => \N__32018\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32018\
        );

    \I__6887\ : Odrv12
    port map (
            O => \N__32037\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__32034\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__32031\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__32028\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6883\ : Odrv12
    port map (
            O => \N__32023\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__32018\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__32005\,
            I => \N__32002\
        );

    \I__6880\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31999\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__31999\,
            I => \N__31996\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__31996\,
            I => \N__31993\
        );

    \I__6877\ : Span4Mux_h
    port map (
            O => \N__31993\,
            I => \N__31990\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__31990\,
            I => \POWERLED.g2\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__31987\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_10_cascade_\
        );

    \I__6874\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31981\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__31981\,
            I => \N__31977\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__31980\,
            I => \N__31971\
        );

    \I__6871\ : Span4Mux_v
    port map (
            O => \N__31977\,
            I => \N__31968\
        );

    \I__6870\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31965\
        );

    \I__6869\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31962\
        );

    \I__6868\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31959\
        );

    \I__6867\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31956\
        );

    \I__6866\ : Span4Mux_s0_v
    port map (
            O => \N__31968\,
            I => \N__31951\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__31965\,
            I => \N__31951\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__31962\,
            I => \N__31946\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__31959\,
            I => \N__31946\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__31956\,
            I => \N__31938\
        );

    \I__6861\ : Sp12to4
    port map (
            O => \N__31951\,
            I => \N__31938\
        );

    \I__6860\ : Span12Mux_v
    port map (
            O => \N__31946\,
            I => \N__31938\
        );

    \I__6859\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31935\
        );

    \I__6858\ : Odrv12
    port map (
            O => \N__31938\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__31935\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6856\ : CascadeMux
    port map (
            O => \N__31930\,
            I => \N__31927\
        );

    \I__6855\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31924\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__31924\,
            I => \N__31921\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__31921\,
            I => \N__31918\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__31918\,
            I => \POWERLED.dutycycle_RNIZ0Z_11\
        );

    \I__6851\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31912\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__31912\,
            I => \POWERLED.g0_1_0\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__31909\,
            I => \POWERLED.m21_e_1_cascade_\
        );

    \I__6848\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31898\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31898\
        );

    \I__6846\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31893\
        );

    \I__6845\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31893\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31890\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31885\
        );

    \I__6842\ : Span4Mux_h
    port map (
            O => \N__31890\,
            I => \N__31885\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__31885\,
            I => \N__31882\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__31882\,
            I => \POWERLED.N_5\
        );

    \I__6839\ : CascadeMux
    port map (
            O => \N__31879\,
            I => \N__31876\
        );

    \I__6838\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31872\
        );

    \I__6837\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31869\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__31872\,
            I => \N__31866\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__31869\,
            I => \N__31863\
        );

    \I__6834\ : Span4Mux_s2_h
    port map (
            O => \N__31866\,
            I => \N__31860\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__31863\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__31860\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__31855\,
            I => \N__31852\
        );

    \I__6830\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31849\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31846\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__31846\,
            I => \POWERLED.mult1_un47_sum_i\
        );

    \I__6827\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31840\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31837\
        );

    \I__6825\ : Span4Mux_h
    port map (
            O => \N__31837\,
            I => \N__31834\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__31834\,
            I => \POWERLED.g2_0_0_0\
        );

    \I__6823\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31820\
        );

    \I__6822\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31820\
        );

    \I__6821\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31820\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__31828\,
            I => \N__31815\
        );

    \I__6819\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31812\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31809\
        );

    \I__6817\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31806\
        );

    \I__6816\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31803\
        );

    \I__6815\ : InMux
    port map (
            O => \N__31815\,
            I => \N__31800\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__31812\,
            I => \N__31797\
        );

    \I__6813\ : Span4Mux_v
    port map (
            O => \N__31809\,
            I => \N__31794\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__31806\,
            I => \N__31791\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31788\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__31800\,
            I => \N__31785\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__31797\,
            I => \N__31778\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__31794\,
            I => \N__31778\
        );

    \I__6807\ : Span4Mux_v
    port map (
            O => \N__31791\,
            I => \N__31778\
        );

    \I__6806\ : Span4Mux_v
    port map (
            O => \N__31788\,
            I => \N__31773\
        );

    \I__6805\ : Span4Mux_h
    port map (
            O => \N__31785\,
            I => \N__31773\
        );

    \I__6804\ : Span4Mux_h
    port map (
            O => \N__31778\,
            I => \N__31770\
        );

    \I__6803\ : Odrv4
    port map (
            O => \N__31773\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__6802\ : Odrv4
    port map (
            O => \N__31770\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__6801\ : CascadeMux
    port map (
            O => \N__31765\,
            I => \POWERLED.g2_0_0_cascade_\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__31762\,
            I => \POWERLED.mult1_un54_sum_s_8_cascade_\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__31759\,
            I => \N__31756\
        );

    \I__6798\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31753\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__31753\,
            I => \N__31750\
        );

    \I__6796\ : Span4Mux_s2_h
    port map (
            O => \N__31750\,
            I => \N__31747\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__31747\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__6794\ : InMux
    port map (
            O => \N__31744\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__31741\,
            I => \N__31738\
        );

    \I__6792\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31735\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__31735\,
            I => \N__31732\
        );

    \I__6790\ : Span4Mux_s2_h
    port map (
            O => \N__31732\,
            I => \N__31729\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__31729\,
            I => \POWERLED.mult1_un47_sum_s_4_sf\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__31726\,
            I => \N__31723\
        );

    \I__6787\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31720\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__31720\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__6785\ : InMux
    port map (
            O => \N__31717\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__6784\ : CascadeMux
    port map (
            O => \N__31714\,
            I => \N__31711\
        );

    \I__6783\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31708\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__31708\,
            I => \N__31705\
        );

    \I__6781\ : Span4Mux_s2_h
    port map (
            O => \N__31705\,
            I => \N__31702\
        );

    \I__6780\ : Odrv4
    port map (
            O => \N__31702\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__31699\,
            I => \N__31696\
        );

    \I__6778\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31693\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__31693\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__6776\ : InMux
    port map (
            O => \N__31690\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__6775\ : InMux
    port map (
            O => \N__31687\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__6774\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31681\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__31681\,
            I => \N__31677\
        );

    \I__6772\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31674\
        );

    \I__6771\ : Span4Mux_h
    port map (
            O => \N__31677\,
            I => \N__31671\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__31674\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__6769\ : Odrv4
    port map (
            O => \N__31671\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__6768\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31663\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__31663\,
            I => \N__31659\
        );

    \I__6766\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31655\
        );

    \I__6765\ : Span12Mux_s10_h
    port map (
            O => \N__31659\,
            I => \N__31651\
        );

    \I__6764\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31648\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31645\
        );

    \I__6762\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31642\
        );

    \I__6761\ : Odrv12
    port map (
            O => \N__31651\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__31648\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__31645\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__31642\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6757\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31628\
        );

    \I__6756\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31625\
        );

    \I__6755\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31622\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__31628\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__31625\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__31622\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__6750\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__31609\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__6748\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__6746\ : Span12Mux_s3_v
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__6745\ : Odrv12
    port map (
            O => \N__31597\,
            I => \POWERLED.un1_clk_100khz_43_and_i_0_d_0\
        );

    \I__6744\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31590\
        );

    \I__6743\ : CascadeMux
    port map (
            O => \N__31593\,
            I => \N__31585\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__31590\,
            I => \N__31582\
        );

    \I__6741\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31575\
        );

    \I__6740\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31575\
        );

    \I__6739\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31575\
        );

    \I__6738\ : Span4Mux_h
    port map (
            O => \N__31582\,
            I => \N__31571\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__31575\,
            I => \N__31568\
        );

    \I__6736\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31565\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__31571\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__6734\ : Odrv12
    port map (
            O => \N__31568\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__31565\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__6732\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31554\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__31557\,
            I => \N__31551\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31545\
        );

    \I__6729\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31538\
        );

    \I__6728\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31538\
        );

    \I__6727\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31538\
        );

    \I__6726\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31535\
        );

    \I__6725\ : Odrv12
    port map (
            O => \N__31545\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__31538\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__31535\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__31528\,
            I => \N__31525\
        );

    \I__6721\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31516\
        );

    \I__6720\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31516\
        );

    \I__6719\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31516\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__31516\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__6717\ : InMux
    port map (
            O => \N__31513\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__6716\ : InMux
    port map (
            O => \N__31510\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__6715\ : InMux
    port map (
            O => \N__31507\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__6714\ : InMux
    port map (
            O => \N__31504\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__6713\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31498\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__31498\,
            I => \N__31493\
        );

    \I__6711\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31490\
        );

    \I__6710\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31487\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__31493\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__31490\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__31487\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__31480\,
            I => \N__31477\
        );

    \I__6705\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31474\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31471\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__31471\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__6702\ : InMux
    port map (
            O => \N__31468\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__31465\,
            I => \N__31462\
        );

    \I__6700\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__31459\,
            I => \N__31456\
        );

    \I__6698\ : Odrv4
    port map (
            O => \N__31456\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__6697\ : InMux
    port map (
            O => \N__31453\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__6696\ : InMux
    port map (
            O => \N__31450\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__6695\ : CascadeMux
    port map (
            O => \N__31447\,
            I => \N__31443\
        );

    \I__6694\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31435\
        );

    \I__6693\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31435\
        );

    \I__6692\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31435\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__31435\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__6690\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31429\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31425\
        );

    \I__6688\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__6687\ : Span4Mux_v
    port map (
            O => \N__31425\,
            I => \N__31419\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__31422\,
            I => \N__31416\
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__31419\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__6684\ : Odrv12
    port map (
            O => \N__31416\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__31411\,
            I => \N__31408\
        );

    \I__6682\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31405\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31402\
        );

    \I__6680\ : Span4Mux_v
    port map (
            O => \N__31402\,
            I => \N__31399\
        );

    \I__6679\ : Odrv4
    port map (
            O => \N__31399\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__6678\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31393\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__31393\,
            I => \N__31390\
        );

    \I__6676\ : Odrv4
    port map (
            O => \N__31390\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__6675\ : InMux
    port map (
            O => \N__31387\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__6674\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31381\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__31381\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__6672\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31375\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__6670\ : Odrv4
    port map (
            O => \N__31372\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__6669\ : InMux
    port map (
            O => \N__31369\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__6668\ : CascadeMux
    port map (
            O => \N__31366\,
            I => \N__31363\
        );

    \I__6667\ : InMux
    port map (
            O => \N__31363\,
            I => \N__31360\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__31360\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__31357\,
            I => \N__31354\
        );

    \I__6664\ : InMux
    port map (
            O => \N__31354\,
            I => \N__31351\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__31351\,
            I => \N__31348\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__31348\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__6661\ : InMux
    port map (
            O => \N__31345\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__6660\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31339\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__31339\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__6658\ : CascadeMux
    port map (
            O => \N__31336\,
            I => \N__31333\
        );

    \I__6657\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31330\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__31330\,
            I => \N__31327\
        );

    \I__6655\ : Odrv12
    port map (
            O => \N__31327\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__6654\ : InMux
    port map (
            O => \N__31324\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__31321\,
            I => \N__31318\
        );

    \I__6652\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31315\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__31315\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__6650\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31309\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__31309\,
            I => \N__31306\
        );

    \I__6648\ : Odrv4
    port map (
            O => \N__31306\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__6647\ : InMux
    port map (
            O => \N__31303\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__6646\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31297\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__31297\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__6644\ : InMux
    port map (
            O => \N__31294\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__6643\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31288\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31284\
        );

    \I__6641\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31281\
        );

    \I__6640\ : Span4Mux_s3_h
    port map (
            O => \N__31284\,
            I => \N__31278\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31275\
        );

    \I__6638\ : Odrv4
    port map (
            O => \N__31278\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__6637\ : Odrv12
    port map (
            O => \N__31275\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__6636\ : CascadeMux
    port map (
            O => \N__31270\,
            I => \N__31267\
        );

    \I__6635\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31261\
        );

    \I__6633\ : Span4Mux_s1_h
    port map (
            O => \N__31261\,
            I => \N__31258\
        );

    \I__6632\ : Odrv4
    port map (
            O => \N__31258\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__6631\ : InMux
    port map (
            O => \N__31255\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__6630\ : InMux
    port map (
            O => \N__31252\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__6629\ : InMux
    port map (
            O => \N__31249\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__6628\ : InMux
    port map (
            O => \N__31246\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__6627\ : InMux
    port map (
            O => \N__31243\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__31240\,
            I => \N__31237\
        );

    \I__6625\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31233\
        );

    \I__6624\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31230\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__31233\,
            I => \HDA_STRAP.count_1_5\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__31230\,
            I => \HDA_STRAP.count_1_5\
        );

    \I__6621\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31222\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__31222\,
            I => \HDA_STRAP.un25_clk_100khz_2\
        );

    \I__6619\ : CascadeMux
    port map (
            O => \N__31219\,
            I => \HDA_STRAP.un25_clk_100khz_3_cascade_\
        );

    \I__6618\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31213\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__31213\,
            I => \N__31210\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__31210\,
            I => \HDA_STRAP.un25_clk_100khz_4\
        );

    \I__6615\ : InMux
    port map (
            O => \N__31207\,
            I => \N__31204\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__31204\,
            I => \N__31201\
        );

    \I__6613\ : Odrv4
    port map (
            O => \N__31201\,
            I => \HDA_STRAP.un25_clk_100khz_14\
        );

    \I__6612\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31195\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__31195\,
            I => \HDA_STRAP.un25_clk_100khz_5\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__31192\,
            I => \N__31189\
        );

    \I__6609\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31185\
        );

    \I__6608\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31182\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__31185\,
            I => \HDA_STRAP.count_1_13\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__31182\,
            I => \HDA_STRAP.count_1_13\
        );

    \I__6605\ : InMux
    port map (
            O => \N__31177\,
            I => \N__31171\
        );

    \I__6604\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31171\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__31171\,
            I => \HDA_STRAP.count_1_3\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__31168\,
            I => \N__31163\
        );

    \I__6601\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31160\
        );

    \I__6600\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31157\
        );

    \I__6599\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31148\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__31160\,
            I => \N__31145\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31142\
        );

    \I__6596\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31133\
        );

    \I__6595\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31133\
        );

    \I__6594\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31133\
        );

    \I__6593\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31133\
        );

    \I__6592\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31128\
        );

    \I__6591\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31128\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__31148\,
            I => \N__31125\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__31145\,
            I => \N__31122\
        );

    \I__6588\ : Span4Mux_s2_h
    port map (
            O => \N__31142\,
            I => \N__31119\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__31133\,
            I => \N__31116\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31113\
        );

    \I__6585\ : Span4Mux_v
    port map (
            O => \N__31125\,
            I => \N__31108\
        );

    \I__6584\ : Span4Mux_v
    port map (
            O => \N__31122\,
            I => \N__31108\
        );

    \I__6583\ : Span4Mux_h
    port map (
            O => \N__31119\,
            I => \N__31103\
        );

    \I__6582\ : Span4Mux_h
    port map (
            O => \N__31116\,
            I => \N__31103\
        );

    \I__6581\ : Span4Mux_h
    port map (
            O => \N__31113\,
            I => \N__31100\
        );

    \I__6580\ : Odrv4
    port map (
            O => \N__31108\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__6579\ : Odrv4
    port map (
            O => \N__31103\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__6578\ : Odrv4
    port map (
            O => \N__31100\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__6577\ : IoInMux
    port map (
            O => \N__31093\,
            I => \N__31090\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31087\
        );

    \I__6575\ : IoSpan4Mux
    port map (
            O => \N__31087\,
            I => \N__31084\
        );

    \I__6574\ : IoSpan4Mux
    port map (
            O => \N__31084\,
            I => \N__31081\
        );

    \I__6573\ : Odrv4
    port map (
            O => \N__31081\,
            I => vpp_en
        );

    \I__6572\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31075\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__31075\,
            I => \N__31072\
        );

    \I__6570\ : Span4Mux_s3_h
    port map (
            O => \N__31072\,
            I => \N__31069\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__31069\,
            I => \N__31066\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__31066\,
            I => \N__31061\
        );

    \I__6567\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31056\
        );

    \I__6566\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31056\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__31061\,
            I => \VPP_VDDQ.N_194\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__31056\,
            I => \VPP_VDDQ.N_194\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__31051\,
            I => \N__31048\
        );

    \I__6562\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31041\
        );

    \I__6561\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31041\
        );

    \I__6560\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31038\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__31041\,
            I => \N__31033\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__31038\,
            I => \N__31030\
        );

    \I__6557\ : InMux
    port map (
            O => \N__31037\,
            I => \N__31025\
        );

    \I__6556\ : InMux
    port map (
            O => \N__31036\,
            I => \N__31025\
        );

    \I__6555\ : Span12Mux_s8_h
    port map (
            O => \N__31033\,
            I => \N__31022\
        );

    \I__6554\ : Span4Mux_h
    port map (
            O => \N__31030\,
            I => \N__31019\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__31025\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6552\ : Odrv12
    port map (
            O => \N__31022\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__31019\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6550\ : InMux
    port map (
            O => \N__31012\,
            I => \N__31009\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__31009\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__31006\,
            I => \N__30993\
        );

    \I__6547\ : InMux
    port map (
            O => \N__31005\,
            I => \N__30989\
        );

    \I__6546\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30984\
        );

    \I__6545\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30984\
        );

    \I__6544\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30981\
        );

    \I__6543\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30978\
        );

    \I__6542\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30975\
        );

    \I__6541\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30972\
        );

    \I__6540\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30969\
        );

    \I__6539\ : InMux
    port map (
            O => \N__30997\,
            I => \N__30964\
        );

    \I__6538\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30964\
        );

    \I__6537\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30959\
        );

    \I__6536\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30959\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__30989\,
            I => \N__30956\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30939\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__30981\,
            I => \N__30936\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__30978\,
            I => \N__30933\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30930\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30927\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__30969\,
            I => \N__30924\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__30964\,
            I => \N__30921\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__30959\,
            I => \N__30918\
        );

    \I__6526\ : Glb2LocalMux
    port map (
            O => \N__30956\,
            I => \N__30871\
        );

    \I__6525\ : CEMux
    port map (
            O => \N__30955\,
            I => \N__30871\
        );

    \I__6524\ : CEMux
    port map (
            O => \N__30954\,
            I => \N__30871\
        );

    \I__6523\ : CEMux
    port map (
            O => \N__30953\,
            I => \N__30871\
        );

    \I__6522\ : CEMux
    port map (
            O => \N__30952\,
            I => \N__30871\
        );

    \I__6521\ : CEMux
    port map (
            O => \N__30951\,
            I => \N__30871\
        );

    \I__6520\ : CEMux
    port map (
            O => \N__30950\,
            I => \N__30871\
        );

    \I__6519\ : CEMux
    port map (
            O => \N__30949\,
            I => \N__30871\
        );

    \I__6518\ : CEMux
    port map (
            O => \N__30948\,
            I => \N__30871\
        );

    \I__6517\ : CEMux
    port map (
            O => \N__30947\,
            I => \N__30871\
        );

    \I__6516\ : CEMux
    port map (
            O => \N__30946\,
            I => \N__30871\
        );

    \I__6515\ : CEMux
    port map (
            O => \N__30945\,
            I => \N__30871\
        );

    \I__6514\ : CEMux
    port map (
            O => \N__30944\,
            I => \N__30871\
        );

    \I__6513\ : CEMux
    port map (
            O => \N__30943\,
            I => \N__30871\
        );

    \I__6512\ : CEMux
    port map (
            O => \N__30942\,
            I => \N__30871\
        );

    \I__6511\ : Glb2LocalMux
    port map (
            O => \N__30939\,
            I => \N__30871\
        );

    \I__6510\ : Glb2LocalMux
    port map (
            O => \N__30936\,
            I => \N__30871\
        );

    \I__6509\ : Glb2LocalMux
    port map (
            O => \N__30933\,
            I => \N__30871\
        );

    \I__6508\ : Glb2LocalMux
    port map (
            O => \N__30930\,
            I => \N__30871\
        );

    \I__6507\ : Glb2LocalMux
    port map (
            O => \N__30927\,
            I => \N__30871\
        );

    \I__6506\ : Glb2LocalMux
    port map (
            O => \N__30924\,
            I => \N__30871\
        );

    \I__6505\ : Glb2LocalMux
    port map (
            O => \N__30921\,
            I => \N__30871\
        );

    \I__6504\ : Glb2LocalMux
    port map (
            O => \N__30918\,
            I => \N__30871\
        );

    \I__6503\ : GlobalMux
    port map (
            O => \N__30871\,
            I => \N__30868\
        );

    \I__6502\ : gio2CtrlBuf
    port map (
            O => \N__30868\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en_g\
        );

    \I__6501\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30862\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__30862\,
            I => \HDA_STRAP.count_1_12\
        );

    \I__6499\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30853\
        );

    \I__6498\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30853\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__30853\,
            I => \HDA_STRAP.count_1_9\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__30850\,
            I => \HDA_STRAP.countZ0Z_12_cascade_\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__30847\,
            I => \N__30844\
        );

    \I__6494\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30838\
        );

    \I__6493\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30838\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__30838\,
            I => \HDA_STRAP.count_1_0_8\
        );

    \I__6491\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30832\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__30832\,
            I => \HDA_STRAP.count_1_0_6\
        );

    \I__6489\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30823\
        );

    \I__6488\ : InMux
    port map (
            O => \N__30828\,
            I => \N__30823\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__30823\,
            I => \HDA_STRAP.count_1_15\
        );

    \I__6486\ : CascadeMux
    port map (
            O => \N__30820\,
            I => \HDA_STRAP.countZ0Z_6_cascade_\
        );

    \I__6485\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30814\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__30814\,
            I => \HDA_STRAP.un25_clk_100khz_6\
        );

    \I__6483\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30805\
        );

    \I__6482\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30805\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__30805\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__6480\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30799\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__30799\,
            I => \HDA_STRAP.un25_clk_100khz_0\
        );

    \I__6478\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30793\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__30793\,
            I => \N__30790\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__30790\,
            I => \VPP_VDDQ.un1_count_2_1_axb_14\
        );

    \I__6475\ : CascadeMux
    port map (
            O => \N__30787\,
            I => \N__30784\
        );

    \I__6474\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30779\
        );

    \I__6473\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30774\
        );

    \I__6472\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30774\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30769\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__30774\,
            I => \N__30769\
        );

    \I__6469\ : Odrv4
    port map (
            O => \N__30769\,
            I => \VPP_VDDQ.count_2_rst_10\
        );

    \I__6468\ : InMux
    port map (
            O => \N__30766\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__6467\ : InMux
    port map (
            O => \N__30763\,
            I => \N__30760\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__30760\,
            I => \N__30757\
        );

    \I__6465\ : Span4Mux_v
    port map (
            O => \N__30757\,
            I => \N__30753\
        );

    \I__6464\ : InMux
    port map (
            O => \N__30756\,
            I => \N__30750\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__30753\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__30750\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__6461\ : InMux
    port map (
            O => \N__30745\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30742\,
            I => \N__30736\
        );

    \I__6459\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30736\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__30736\,
            I => \N__30733\
        );

    \I__6457\ : Span4Mux_s2_v
    port map (
            O => \N__30733\,
            I => \N__30730\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__30730\,
            I => \VPP_VDDQ.count_2_rst_9\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__30727\,
            I => \N__30724\
        );

    \I__6454\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30721\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30717\
        );

    \I__6452\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30714\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__30717\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__30714\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__30709\,
            I => \HDA_STRAP.count_1_0_cascade_\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__30706\,
            I => \HDA_STRAP.countZ0Z_0_cascade_\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__30703\,
            I => \HDA_STRAP.un25_clk_100khz_13_cascade_\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__30700\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_\
        );

    \I__6445\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30694\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__30694\,
            I => \HDA_STRAP.count_1_0_0\
        );

    \I__6443\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30688\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__30688\,
            I => \HDA_STRAP.un25_clk_100khz_7\
        );

    \I__6441\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30679\
        );

    \I__6440\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30679\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__30679\,
            I => \N__30676\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__30676\,
            I => \VPP_VDDQ.count_2_rst_2\
        );

    \I__6437\ : InMux
    port map (
            O => \N__30673\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__6436\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30667\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__30667\,
            I => \N__30664\
        );

    \I__6434\ : Odrv12
    port map (
            O => \N__30664\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__6433\ : CascadeMux
    port map (
            O => \N__30661\,
            I => \N__30658\
        );

    \I__6432\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30655\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30650\
        );

    \I__6430\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30645\
        );

    \I__6429\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30645\
        );

    \I__6428\ : Span4Mux_v
    port map (
            O => \N__30650\,
            I => \N__30640\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__30645\,
            I => \N__30640\
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__30640\,
            I => \VPP_VDDQ.count_2_rst_1\
        );

    \I__6425\ : InMux
    port map (
            O => \N__30637\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__6424\ : InMux
    port map (
            O => \N__30634\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__6423\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30628\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__30628\,
            I => \N__30624\
        );

    \I__6421\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30621\
        );

    \I__6420\ : Span4Mux_s3_v
    port map (
            O => \N__30624\,
            I => \N__30618\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__30621\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__30618\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__6417\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30607\
        );

    \I__6416\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30607\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__30607\,
            I => \N__30604\
        );

    \I__6414\ : Span4Mux_h
    port map (
            O => \N__30604\,
            I => \N__30601\
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__30601\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\
        );

    \I__6412\ : InMux
    port map (
            O => \N__30598\,
            I => \bfn_11_3_0_\
        );

    \I__6411\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30592\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__30592\,
            I => \N__30589\
        );

    \I__6409\ : Span4Mux_s2_h
    port map (
            O => \N__30589\,
            I => \N__30586\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__30586\,
            I => \VPP_VDDQ.un1_count_2_1_axb_10\
        );

    \I__6407\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30574\
        );

    \I__6406\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30574\
        );

    \I__6405\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30574\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__30574\,
            I => \N__30571\
        );

    \I__6403\ : Span4Mux_h
    port map (
            O => \N__30571\,
            I => \N__30568\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__30568\,
            I => \VPP_VDDQ.count_2_rst_14\
        );

    \I__6401\ : InMux
    port map (
            O => \N__30565\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__6400\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30559\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30555\
        );

    \I__6398\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30552\
        );

    \I__6397\ : Span4Mux_s2_h
    port map (
            O => \N__30555\,
            I => \N__30549\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__30552\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__30549\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__6394\ : InMux
    port map (
            O => \N__30544\,
            I => \N__30540\
        );

    \I__6393\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30537\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30532\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30532\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__30532\,
            I => \N__30529\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__30529\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__6388\ : InMux
    port map (
            O => \N__30526\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__6387\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30520\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__30520\,
            I => \N__30517\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__30517\,
            I => \VPP_VDDQ.un1_count_2_1_axb_12\
        );

    \I__6384\ : InMux
    port map (
            O => \N__30514\,
            I => \N__30505\
        );

    \I__6383\ : InMux
    port map (
            O => \N__30513\,
            I => \N__30505\
        );

    \I__6382\ : InMux
    port map (
            O => \N__30512\,
            I => \N__30505\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__30505\,
            I => \N__30502\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__30502\,
            I => \VPP_VDDQ.count_2_rst_12\
        );

    \I__6379\ : InMux
    port map (
            O => \N__30499\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__6378\ : InMux
    port map (
            O => \N__30496\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__6377\ : CascadeMux
    port map (
            O => \N__30493\,
            I => \VPP_VDDQ.count_2_rst_5_cascade_\
        );

    \I__6376\ : CascadeMux
    port map (
            O => \N__30490\,
            I => \VPP_VDDQ.count_2Z0Z_3_cascade_\
        );

    \I__6375\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30484\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__30484\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__30481\,
            I => \N__30477\
        );

    \I__6372\ : CascadeMux
    port map (
            O => \N__30480\,
            I => \N__30474\
        );

    \I__6371\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30471\
        );

    \I__6370\ : InMux
    port map (
            O => \N__30474\,
            I => \N__30468\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__30471\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__30468\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2\
        );

    \I__6367\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30457\
        );

    \I__6366\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30457\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__30457\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\
        );

    \I__6364\ : InMux
    port map (
            O => \N__30454\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__30451\,
            I => \N__30447\
        );

    \I__6362\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30443\
        );

    \I__6361\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30440\
        );

    \I__6360\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30437\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__30443\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__30440\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__30437\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__6356\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30424\
        );

    \I__6355\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30424\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__30424\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\
        );

    \I__6353\ : InMux
    port map (
            O => \N__30421\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__6352\ : InMux
    port map (
            O => \N__30418\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__6351\ : InMux
    port map (
            O => \N__30415\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__30412\,
            I => \POWERLED.dutycycleZ0Z_11_cascade_\
        );

    \I__6349\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30406\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__30406\,
            I => \POWERLED.dutycycle_RNIZ0Z_10\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__30403\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__30400\,
            I => \POWERLED.un1_dutycycle_53_axb_12_cascade_\
        );

    \I__6345\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30392\
        );

    \I__6344\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30389\
        );

    \I__6343\ : InMux
    port map (
            O => \N__30395\,
            I => \N__30383\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__30392\,
            I => \N__30378\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30378\
        );

    \I__6340\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30375\
        );

    \I__6339\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30370\
        );

    \I__6338\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30367\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__30383\,
            I => \N__30362\
        );

    \I__6336\ : Span4Mux_v
    port map (
            O => \N__30378\,
            I => \N__30362\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__30375\,
            I => \N__30359\
        );

    \I__6334\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30354\
        );

    \I__6333\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30354\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__30370\,
            I => \N__30349\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__30367\,
            I => \N__30349\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__30362\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__30359\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__30354\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__30349\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6326\ : CascadeMux
    port map (
            O => \N__30340\,
            I => \N__30337\
        );

    \I__6325\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30334\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__30331\,
            I => \POWERLED.dutycycle_RNIZ0Z_15\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__30328\,
            I => \POWERLED.un1_dutycycle_53_axb_14_cascade_\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30322\
        );

    \I__6320\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30319\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__30319\,
            I => \N__30316\
        );

    \I__6318\ : Odrv12
    port map (
            O => \N__30316\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_14\
        );

    \I__6317\ : InMux
    port map (
            O => \N__30313\,
            I => \N__30310\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__30310\,
            I => \VPP_VDDQ.count_2_rst_6\
        );

    \I__6315\ : CascadeMux
    port map (
            O => \N__30307\,
            I => \VPP_VDDQ.count_2_rst_6_cascade_\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__30304\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2_cascade_\
        );

    \I__6313\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30295\
        );

    \I__6312\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30295\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__30295\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__30292\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__30289\,
            I => \POWERLED.g0_4_1_cascade_\
        );

    \I__6308\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30283\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__30283\,
            I => \POWERLED.un1_dutycycle_53_25_1_1\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__30280\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_7_cascade_\
        );

    \I__6305\ : InMux
    port map (
            O => \N__30277\,
            I => \N__30267\
        );

    \I__6304\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30267\
        );

    \I__6303\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30262\
        );

    \I__6302\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30257\
        );

    \I__6301\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30257\
        );

    \I__6300\ : CascadeMux
    port map (
            O => \N__30272\,
            I => \N__30254\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30251\
        );

    \I__6298\ : InMux
    port map (
            O => \N__30266\,
            I => \N__30247\
        );

    \I__6297\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30244\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__30262\,
            I => \N__30236\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30233\
        );

    \I__6294\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30230\
        );

    \I__6293\ : Span4Mux_h
    port map (
            O => \N__30251\,
            I => \N__30227\
        );

    \I__6292\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30224\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__30247\,
            I => \N__30219\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__30244\,
            I => \N__30219\
        );

    \I__6289\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30210\
        );

    \I__6288\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30210\
        );

    \I__6287\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30210\
        );

    \I__6286\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30210\
        );

    \I__6285\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30207\
        );

    \I__6284\ : Span4Mux_h
    port map (
            O => \N__30236\,
            I => \N__30200\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__30233\,
            I => \N__30200\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__30230\,
            I => \N__30200\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__30227\,
            I => \tmp_1_rep1_RNIC08FV_0\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__30224\,
            I => \tmp_1_rep1_RNIC08FV_0\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__30219\,
            I => \tmp_1_rep1_RNIC08FV_0\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__30210\,
            I => \tmp_1_rep1_RNIC08FV_0\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__30207\,
            I => \tmp_1_rep1_RNIC08FV_0\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__30200\,
            I => \tmp_1_rep1_RNIC08FV_0\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__30187\,
            I => \N__30184\
        );

    \I__6274\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30181\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__6272\ : Odrv12
    port map (
            O => \N__30178\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_9\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__30175\,
            I => \N__30163\
        );

    \I__6270\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30156\
        );

    \I__6269\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30156\
        );

    \I__6268\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30156\
        );

    \I__6267\ : CascadeMux
    port map (
            O => \N__30171\,
            I => \N__30150\
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__30170\,
            I => \N__30147\
        );

    \I__6265\ : InMux
    port map (
            O => \N__30169\,
            I => \N__30143\
        );

    \I__6264\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30134\
        );

    \I__6263\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30134\
        );

    \I__6262\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30134\
        );

    \I__6261\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30130\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__30156\,
            I => \N__30127\
        );

    \I__6259\ : InMux
    port map (
            O => \N__30155\,
            I => \N__30120\
        );

    \I__6258\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30120\
        );

    \I__6257\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30120\
        );

    \I__6256\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30113\
        );

    \I__6255\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30113\
        );

    \I__6254\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30113\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__30143\,
            I => \N__30110\
        );

    \I__6252\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30107\
        );

    \I__6251\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30104\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30100\
        );

    \I__6249\ : CascadeMux
    port map (
            O => \N__30133\,
            I => \N__30097\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__30130\,
            I => \N__30094\
        );

    \I__6247\ : Span4Mux_s1_v
    port map (
            O => \N__30127\,
            I => \N__30085\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__30120\,
            I => \N__30085\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__30113\,
            I => \N__30085\
        );

    \I__6244\ : Span4Mux_s1_v
    port map (
            O => \N__30110\,
            I => \N__30082\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30077\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__30104\,
            I => \N__30077\
        );

    \I__6241\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30074\
        );

    \I__6240\ : Span4Mux_s1_v
    port map (
            O => \N__30100\,
            I => \N__30071\
        );

    \I__6239\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30066\
        );

    \I__6238\ : Span4Mux_v
    port map (
            O => \N__30094\,
            I => \N__30063\
        );

    \I__6237\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30060\
        );

    \I__6236\ : InMux
    port map (
            O => \N__30092\,
            I => \N__30057\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__30085\,
            I => \N__30054\
        );

    \I__6234\ : Span4Mux_v
    port map (
            O => \N__30082\,
            I => \N__30051\
        );

    \I__6233\ : Span4Mux_v
    port map (
            O => \N__30077\,
            I => \N__30044\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__30074\,
            I => \N__30044\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__30071\,
            I => \N__30044\
        );

    \I__6230\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30039\
        );

    \I__6229\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30039\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__30066\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6227\ : Odrv4
    port map (
            O => \N__30063\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__30060\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__30057\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__30054\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6223\ : Odrv4
    port map (
            O => \N__30051\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6222\ : Odrv4
    port map (
            O => \N__30044\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__30039\,
            I => \POWERLED.func_m1_0_a2Z0Z_0\
        );

    \I__6220\ : InMux
    port map (
            O => \N__30022\,
            I => \N__30018\
        );

    \I__6219\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30015\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__30018\,
            I => \N__30012\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__30009\
        );

    \I__6216\ : Span4Mux_s2_v
    port map (
            O => \N__30012\,
            I => \N__30006\
        );

    \I__6215\ : Odrv4
    port map (
            O => \N__30009\,
            I => \POWERLED.N_235_N\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__30006\,
            I => \POWERLED.N_235_N\
        );

    \I__6213\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29998\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__29998\,
            I => \POWERLED.dutycycle_eena_9\
        );

    \I__6211\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29989\
        );

    \I__6210\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29989\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29986\
        );

    \I__6208\ : Odrv12
    port map (
            O => \N__29986\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1\
        );

    \I__6207\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29977\
        );

    \I__6206\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29977\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__29977\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__29974\,
            I => \POWERLED.dutycycle_eena_9_cascade_\
        );

    \I__6203\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29966\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__29970\,
            I => \N__29958\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \N__29952\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__29966\,
            I => \N__29938\
        );

    \I__6199\ : IoInMux
    port map (
            O => \N__29965\,
            I => \N__29935\
        );

    \I__6198\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29929\
        );

    \I__6197\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29924\
        );

    \I__6196\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29924\
        );

    \I__6195\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29915\
        );

    \I__6194\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29915\
        );

    \I__6193\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29915\
        );

    \I__6192\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29915\
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__29955\,
            I => \N__29912\
        );

    \I__6190\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29908\
        );

    \I__6189\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29905\
        );

    \I__6188\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29902\
        );

    \I__6187\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29897\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29897\
        );

    \I__6185\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29894\
        );

    \I__6184\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29889\
        );

    \I__6183\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29889\
        );

    \I__6182\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29886\
        );

    \I__6181\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29883\
        );

    \I__6180\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29880\
        );

    \I__6179\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29877\
        );

    \I__6178\ : Span4Mux_v
    port map (
            O => \N__29938\,
            I => \N__29874\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__29935\,
            I => \N__29871\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29866\
        );

    \I__6175\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29866\
        );

    \I__6174\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29863\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__29929\,
            I => \N__29860\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__29924\,
            I => \N__29855\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__29915\,
            I => \N__29855\
        );

    \I__6170\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29850\
        );

    \I__6169\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29850\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__29908\,
            I => \N__29847\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__29905\,
            I => \N__29844\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__29902\,
            I => \N__29841\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__29897\,
            I => \N__29832\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29832\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__29889\,
            I => \N__29832\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__29886\,
            I => \N__29832\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29829\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29826\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29823\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__29874\,
            I => \N__29818\
        );

    \I__6157\ : Span4Mux_s1_h
    port map (
            O => \N__29871\,
            I => \N__29818\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29815\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29806\
        );

    \I__6154\ : Span4Mux_h
    port map (
            O => \N__29860\,
            I => \N__29806\
        );

    \I__6153\ : Span4Mux_s2_v
    port map (
            O => \N__29855\,
            I => \N__29806\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__29850\,
            I => \N__29806\
        );

    \I__6151\ : Span4Mux_s2_v
    port map (
            O => \N__29847\,
            I => \N__29801\
        );

    \I__6150\ : Span4Mux_s2_v
    port map (
            O => \N__29844\,
            I => \N__29801\
        );

    \I__6149\ : Span4Mux_s2_v
    port map (
            O => \N__29841\,
            I => \N__29796\
        );

    \I__6148\ : Span4Mux_s2_v
    port map (
            O => \N__29832\,
            I => \N__29796\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__29829\,
            I => \N__29793\
        );

    \I__6146\ : Span4Mux_s3_v
    port map (
            O => \N__29826\,
            I => \N__29790\
        );

    \I__6145\ : Span4Mux_h
    port map (
            O => \N__29823\,
            I => \N__29785\
        );

    \I__6144\ : Span4Mux_h
    port map (
            O => \N__29818\,
            I => \N__29785\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__29815\,
            I => \N__29778\
        );

    \I__6142\ : Span4Mux_v
    port map (
            O => \N__29806\,
            I => \N__29778\
        );

    \I__6141\ : Span4Mux_v
    port map (
            O => \N__29801\,
            I => \N__29778\
        );

    \I__6140\ : Span4Mux_v
    port map (
            O => \N__29796\,
            I => \N__29775\
        );

    \I__6139\ : Odrv4
    port map (
            O => \N__29793\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__29790\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6137\ : Odrv4
    port map (
            O => \N__29785\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6136\ : Odrv4
    port map (
            O => \N__29778\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__29775\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6134\ : InMux
    port map (
            O => \N__29764\,
            I => \POWERLED.CO2\
        );

    \I__6133\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29755\
        );

    \I__6132\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29755\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29752\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__29752\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__6128\ : InMux
    port map (
            O => \N__29746\,
            I => \N__29743\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__29743\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__6126\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29736\
        );

    \I__6125\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29733\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__29736\,
            I => \N__29723\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__29733\,
            I => \N__29723\
        );

    \I__6122\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29720\
        );

    \I__6121\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29715\
        );

    \I__6120\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29715\
        );

    \I__6119\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29712\
        );

    \I__6118\ : CascadeMux
    port map (
            O => \N__29728\,
            I => \N__29709\
        );

    \I__6117\ : Span4Mux_s3_v
    port map (
            O => \N__29723\,
            I => \N__29706\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__29720\,
            I => \N__29701\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29701\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__29712\,
            I => \N__29698\
        );

    \I__6113\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29695\
        );

    \I__6112\ : Span4Mux_v
    port map (
            O => \N__29706\,
            I => \N__29690\
        );

    \I__6111\ : Span4Mux_s3_v
    port map (
            O => \N__29701\,
            I => \N__29690\
        );

    \I__6110\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29687\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29684\
        );

    \I__6108\ : Odrv4
    port map (
            O => \N__29690\,
            I => \POWERLED.N_428\
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__29687\,
            I => \POWERLED.N_428\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__29684\,
            I => \POWERLED.N_428\
        );

    \I__6105\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29674\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__29674\,
            I => \N__29671\
        );

    \I__6103\ : Span4Mux_h
    port map (
            O => \N__29671\,
            I => \N__29668\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__29668\,
            I => \POWERLED.un1_dutycycle_53_axb_13_1\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__6100\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29659\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__29659\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_13\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__29656\,
            I => \N__29653\
        );

    \I__6097\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29650\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__29650\,
            I => \N__29647\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__29647\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__29644\,
            I => \N__29640\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__29643\,
            I => \N__29635\
        );

    \I__6092\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29628\
        );

    \I__6091\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29628\
        );

    \I__6090\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29628\
        );

    \I__6089\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29625\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__29628\,
            I => \N__29622\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__29625\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__29622\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__29617\,
            I => \N__29613\
        );

    \I__6084\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29607\
        );

    \I__6083\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29607\
        );

    \I__6082\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29604\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__29607\,
            I => \N__29601\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__29604\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__29601\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__6078\ : CascadeMux
    port map (
            O => \N__29596\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_\
        );

    \I__6077\ : CascadeMux
    port map (
            O => \N__29593\,
            I => \N__29590\
        );

    \I__6076\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29587\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__29587\,
            I => \N__29584\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__29584\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_7\
        );

    \I__6073\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29577\
        );

    \I__6072\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29574\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__29577\,
            I => \N__29571\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__29574\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__6069\ : Odrv4
    port map (
            O => \N__29571\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__29566\,
            I => \N__29563\
        );

    \I__6067\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29560\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__29560\,
            I => \N__29556\
        );

    \I__6065\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29553\
        );

    \I__6064\ : Span4Mux_s3_h
    port map (
            O => \N__29556\,
            I => \N__29550\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__29553\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__6062\ : Odrv4
    port map (
            O => \N__29550\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__6061\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29541\
        );

    \I__6060\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29538\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29535\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__29538\,
            I => \POWERLED.dutycycle_en_6\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__29535\,
            I => \POWERLED.dutycycle_en_6\
        );

    \I__6056\ : InMux
    port map (
            O => \N__29530\,
            I => \bfn_9_13_0_\
        );

    \I__6055\ : InMux
    port map (
            O => \N__29527\,
            I => \POWERLED.un1_dutycycle_53_cry_8\
        );

    \I__6054\ : InMux
    port map (
            O => \N__29524\,
            I => \POWERLED.un1_dutycycle_53_cry_9\
        );

    \I__6053\ : InMux
    port map (
            O => \N__29521\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__6052\ : InMux
    port map (
            O => \N__29518\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__6051\ : InMux
    port map (
            O => \N__29515\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__6050\ : InMux
    port map (
            O => \N__29512\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__6048\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29503\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29500\
        );

    \I__6046\ : Span4Mux_h
    port map (
            O => \N__29500\,
            I => \N__29497\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__29497\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_15\
        );

    \I__6044\ : InMux
    port map (
            O => \N__29494\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__6043\ : InMux
    port map (
            O => \N__29491\,
            I => \bfn_9_14_0_\
        );

    \I__6042\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29485\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__29485\,
            I => \N__29481\
        );

    \I__6040\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29478\
        );

    \I__6039\ : Span4Mux_v
    port map (
            O => \N__29481\,
            I => \N__29475\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__29478\,
            I => \N__29472\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__29475\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__6036\ : Odrv12
    port map (
            O => \N__29472\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__6035\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29463\
        );

    \I__6034\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29460\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__29463\,
            I => \N__29455\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29455\
        );

    \I__6031\ : Span4Mux_v
    port map (
            O => \N__29455\,
            I => \N__29452\
        );

    \I__6030\ : Odrv4
    port map (
            O => \N__29452\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__6029\ : InMux
    port map (
            O => \N__29449\,
            I => \POWERLED.un1_dutycycle_53_cry_0\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__29446\,
            I => \N__29443\
        );

    \I__6027\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29440\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29437\
        );

    \I__6025\ : Span4Mux_v
    port map (
            O => \N__29437\,
            I => \N__29434\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__29434\,
            I => \POWERLED.dutycycle_RNIZ0Z_2\
        );

    \I__6023\ : InMux
    port map (
            O => \N__29431\,
            I => \N__29428\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__29428\,
            I => \N__29424\
        );

    \I__6021\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29421\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__29424\,
            I => \N__29418\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__29421\,
            I => \N__29415\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__29418\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__6017\ : Odrv12
    port map (
            O => \N__29415\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__6016\ : InMux
    port map (
            O => \N__29410\,
            I => \POWERLED.un1_dutycycle_53_cry_1\
        );

    \I__6015\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29404\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__29404\,
            I => \N__29401\
        );

    \I__6013\ : Span4Mux_s3_h
    port map (
            O => \N__29401\,
            I => \N__29398\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__29398\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_2\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__29395\,
            I => \N__29388\
        );

    \I__6010\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29384\
        );

    \I__6009\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29378\
        );

    \I__6008\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29378\
        );

    \I__6007\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29375\
        );

    \I__6006\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29370\
        );

    \I__6005\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29370\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__29384\,
            I => \N__29366\
        );

    \I__6003\ : CascadeMux
    port map (
            O => \N__29383\,
            I => \N__29363\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__29378\,
            I => \N__29358\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__29375\,
            I => \N__29358\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__29370\,
            I => \N__29355\
        );

    \I__5999\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29352\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__29366\,
            I => \N__29349\
        );

    \I__5997\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29346\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__29358\,
            I => \N__29340\
        );

    \I__5995\ : Span4Mux_h
    port map (
            O => \N__29355\,
            I => \N__29340\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__29352\,
            I => \N__29337\
        );

    \I__5993\ : Span4Mux_h
    port map (
            O => \N__29349\,
            I => \N__29332\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29329\
        );

    \I__5991\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29326\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__29340\,
            I => \N__29323\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__29337\,
            I => \N__29320\
        );

    \I__5988\ : InMux
    port map (
            O => \N__29336\,
            I => \N__29315\
        );

    \I__5987\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29315\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__29332\,
            I => \POWERLED.dutycycle\
        );

    \I__5985\ : Odrv4
    port map (
            O => \N__29329\,
            I => \POWERLED.dutycycle\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__29326\,
            I => \POWERLED.dutycycle\
        );

    \I__5983\ : Odrv4
    port map (
            O => \N__29323\,
            I => \POWERLED.dutycycle\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__29320\,
            I => \POWERLED.dutycycle\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__29315\,
            I => \POWERLED.dutycycle\
        );

    \I__5980\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29299\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__29299\,
            I => \N__29295\
        );

    \I__5978\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29292\
        );

    \I__5977\ : Span4Mux_h
    port map (
            O => \N__29295\,
            I => \N__29289\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__29292\,
            I => \N__29286\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__29289\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__29286\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__5973\ : InMux
    port map (
            O => \N__29281\,
            I => \POWERLED.un1_dutycycle_53_cry_2\
        );

    \I__5972\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29275\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__29272\,
            I => \N__29269\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__29269\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_3\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__5967\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29259\
        );

    \I__5966\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29256\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__29259\,
            I => \N__29253\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__29256\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_7\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__29253\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_7\
        );

    \I__5962\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29245\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29242\
        );

    \I__5960\ : Span4Mux_v
    port map (
            O => \N__29242\,
            I => \N__29238\
        );

    \I__5959\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29235\
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__29238\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__29235\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__5956\ : InMux
    port map (
            O => \N__29230\,
            I => \POWERLED.un1_dutycycle_53_cry_3\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__29227\,
            I => \N__29224\
        );

    \I__5954\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29221\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29218\
        );

    \I__5952\ : Span4Mux_s3_h
    port map (
            O => \N__29218\,
            I => \N__29215\
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__29215\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_8\
        );

    \I__5950\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29206\
        );

    \I__5949\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29206\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__29206\,
            I => \N__29203\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__29203\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__5946\ : InMux
    port map (
            O => \N__29200\,
            I => \POWERLED.un1_dutycycle_53_cry_4\
        );

    \I__5945\ : InMux
    port map (
            O => \N__29197\,
            I => \N__29194\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__29194\,
            I => \N__29190\
        );

    \I__5943\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29187\
        );

    \I__5942\ : Odrv4
    port map (
            O => \N__29190\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__29187\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__5940\ : InMux
    port map (
            O => \N__29182\,
            I => \POWERLED.un1_dutycycle_53_cry_5\
        );

    \I__5939\ : InMux
    port map (
            O => \N__29179\,
            I => \POWERLED.un1_dutycycle_53_cry_6\
        );

    \I__5938\ : InMux
    port map (
            O => \N__29176\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__29173\,
            I => \N__29170\
        );

    \I__5936\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29162\
        );

    \I__5935\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29162\
        );

    \I__5934\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29157\
        );

    \I__5933\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29157\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__29162\,
            I => \N__29152\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__29157\,
            I => \N__29152\
        );

    \I__5930\ : Span4Mux_v
    port map (
            O => \N__29152\,
            I => \N__29148\
        );

    \I__5929\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29145\
        );

    \I__5928\ : Odrv4
    port map (
            O => \N__29148\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__29145\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__29140\,
            I => \N__29136\
        );

    \I__5925\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29128\
        );

    \I__5924\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29128\
        );

    \I__5923\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29128\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__29128\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__5921\ : InMux
    port map (
            O => \N__29125\,
            I => \N__29122\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__29122\,
            I => \N__29119\
        );

    \I__5919\ : Span12Mux_s4_v
    port map (
            O => \N__29119\,
            I => \N__29115\
        );

    \I__5918\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29112\
        );

    \I__5917\ : Odrv12
    port map (
            O => \N__29115\,
            I => \POWERLED.g0_i_o3_0\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__29112\,
            I => \POWERLED.g0_i_o3_0\
        );

    \I__5915\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29103\
        );

    \I__5914\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29100\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29097\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__29100\,
            I => \N__29093\
        );

    \I__5911\ : Span4Mux_v
    port map (
            O => \N__29097\,
            I => \N__29089\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__29096\,
            I => \N__29086\
        );

    \I__5909\ : Span4Mux_v
    port map (
            O => \N__29093\,
            I => \N__29083\
        );

    \I__5908\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29080\
        );

    \I__5907\ : Span4Mux_h
    port map (
            O => \N__29089\,
            I => \N__29077\
        );

    \I__5906\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29074\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__29083\,
            I => \N__29069\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29069\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__29077\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__29074\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5901\ : Odrv4
    port map (
            O => \N__29069\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__29062\,
            I => \N__29059\
        );

    \I__5899\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29056\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__29056\,
            I => \N__29052\
        );

    \I__5897\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29049\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__29052\,
            I => \N__29046\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29043\
        );

    \I__5894\ : Span4Mux_h
    port map (
            O => \N__29046\,
            I => \N__29040\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__29043\,
            I => \N__29037\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__29040\,
            I => \POWERLED.N_8\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__29037\,
            I => \POWERLED.N_8\
        );

    \I__5890\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29029\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__29029\,
            I => \N__29026\
        );

    \I__5888\ : Span4Mux_v
    port map (
            O => \N__29026\,
            I => \N__29023\
        );

    \I__5887\ : Span4Mux_h
    port map (
            O => \N__29023\,
            I => \N__29019\
        );

    \I__5886\ : InMux
    port map (
            O => \N__29022\,
            I => \N__29016\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__29019\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__29016\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__5883\ : SRMux
    port map (
            O => \N__29011\,
            I => \N__29008\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__29008\,
            I => \N__29005\
        );

    \I__5881\ : Span4Mux_v
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__5880\ : Span4Mux_s3_h
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__28999\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__5878\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \POWERLED.mult1_un40_sum_i_5_cascade_\
        );

    \I__5877\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__5875\ : Span4Mux_v
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__5874\ : Span4Mux_h
    port map (
            O => \N__28984\,
            I => \N__28981\
        );

    \I__5873\ : Span4Mux_v
    port map (
            O => \N__28981\,
            I => \N__28978\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__28978\,
            I => \RSMRST_PWRGD.count_4_7\
        );

    \I__5871\ : CEMux
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28966\
        );

    \I__5869\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28962\
        );

    \I__5868\ : CEMux
    port map (
            O => \N__28970\,
            I => \N__28956\
        );

    \I__5867\ : CEMux
    port map (
            O => \N__28969\,
            I => \N__28951\
        );

    \I__5866\ : Span4Mux_h
    port map (
            O => \N__28966\,
            I => \N__28948\
        );

    \I__5865\ : CEMux
    port map (
            O => \N__28965\,
            I => \N__28945\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28942\
        );

    \I__5863\ : CEMux
    port map (
            O => \N__28961\,
            I => \N__28938\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__28960\,
            I => \N__28935\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__28959\,
            I => \N__28925\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28920\
        );

    \I__5859\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28915\
        );

    \I__5858\ : CEMux
    port map (
            O => \N__28954\,
            I => \N__28915\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28910\
        );

    \I__5856\ : Sp12to4
    port map (
            O => \N__28948\,
            I => \N__28910\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28906\
        );

    \I__5854\ : Span4Mux_h
    port map (
            O => \N__28942\,
            I => \N__28903\
        );

    \I__5853\ : CEMux
    port map (
            O => \N__28941\,
            I => \N__28895\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__28938\,
            I => \N__28892\
        );

    \I__5851\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28889\
        );

    \I__5850\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28884\
        );

    \I__5849\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28884\
        );

    \I__5848\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28875\
        );

    \I__5847\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28875\
        );

    \I__5846\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28875\
        );

    \I__5845\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28875\
        );

    \I__5844\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28866\
        );

    \I__5843\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28866\
        );

    \I__5842\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28866\
        );

    \I__5841\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28866\
        );

    \I__5840\ : Span4Mux_s1_h
    port map (
            O => \N__28920\,
            I => \N__28861\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__28915\,
            I => \N__28856\
        );

    \I__5838\ : Span12Mux_s7_v
    port map (
            O => \N__28910\,
            I => \N__28856\
        );

    \I__5837\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28853\
        );

    \I__5836\ : Span4Mux_v
    port map (
            O => \N__28906\,
            I => \N__28848\
        );

    \I__5835\ : Span4Mux_h
    port map (
            O => \N__28903\,
            I => \N__28848\
        );

    \I__5834\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28837\
        );

    \I__5833\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28837\
        );

    \I__5832\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28837\
        );

    \I__5831\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28837\
        );

    \I__5830\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28837\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__28895\,
            I => \N__28824\
        );

    \I__5828\ : Span4Mux_h
    port map (
            O => \N__28892\,
            I => \N__28824\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__28889\,
            I => \N__28824\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28824\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__28875\,
            I => \N__28824\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__28866\,
            I => \N__28824\
        );

    \I__5823\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28819\
        );

    \I__5822\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28819\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__28861\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5820\ : Odrv12
    port map (
            O => \N__28856\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__28853\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__28848\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__28837\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__28824\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__28819\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__5814\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28801\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28797\
        );

    \I__5812\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28794\
        );

    \I__5811\ : Span4Mux_v
    port map (
            O => \N__28797\,
            I => \N__28791\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__28794\,
            I => \N__28788\
        );

    \I__5809\ : Span4Mux_h
    port map (
            O => \N__28791\,
            I => \N__28785\
        );

    \I__5808\ : Span4Mux_h
    port map (
            O => \N__28788\,
            I => \N__28782\
        );

    \I__5807\ : Span4Mux_h
    port map (
            O => \N__28785\,
            I => \N__28779\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__28782\,
            I => \RSMRST_PWRGD.count_rst_12\
        );

    \I__5805\ : Odrv4
    port map (
            O => \N__28779\,
            I => \RSMRST_PWRGD.count_rst_12\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__28774\,
            I => \N__28771\
        );

    \I__5803\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28768\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28765\
        );

    \I__5801\ : Span4Mux_v
    port map (
            O => \N__28765\,
            I => \N__28761\
        );

    \I__5800\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28758\
        );

    \I__5799\ : Sp12to4
    port map (
            O => \N__28761\,
            I => \N__28753\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__28758\,
            I => \N__28753\
        );

    \I__5797\ : Span12Mux_s8_h
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__5796\ : Odrv12
    port map (
            O => \N__28750\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__5795\ : CascadeMux
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__5794\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28741\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__28741\,
            I => \N__28738\
        );

    \I__5792\ : Span4Mux_h
    port map (
            O => \N__28738\,
            I => \N__28735\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__28735\,
            I => \POWERLED.mult1_un89_sum_i_8\
        );

    \I__5790\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28728\
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__28731\,
            I => \N__28725\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__28728\,
            I => \N__28720\
        );

    \I__5787\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28715\
        );

    \I__5786\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28715\
        );

    \I__5785\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28712\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__28720\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__28715\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__28712\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__5781\ : CascadeMux
    port map (
            O => \N__28705\,
            I => \N__28702\
        );

    \I__5780\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28699\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__28699\,
            I => \POWERLED.un85_clk_100khz_2\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__28696\,
            I => \N__28693\
        );

    \I__5777\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__28690\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__5775\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__5773\ : Span4Mux_v
    port map (
            O => \N__28681\,
            I => \N__28678\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__28678\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__5771\ : InMux
    port map (
            O => \N__28675\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__28672\,
            I => \N__28669\
        );

    \I__5769\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28666\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28663\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__28663\,
            I => \N__28660\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__28660\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__5765\ : InMux
    port map (
            O => \N__28657\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__5764\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28651\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__5762\ : Span4Mux_v
    port map (
            O => \N__28648\,
            I => \N__28645\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__28645\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__5760\ : InMux
    port map (
            O => \N__28642\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__28639\,
            I => \N__28636\
        );

    \I__5758\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28633\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__5756\ : Span4Mux_v
    port map (
            O => \N__28630\,
            I => \N__28627\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__28627\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__5754\ : InMux
    port map (
            O => \N__28624\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__5753\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28615\
        );

    \I__5751\ : Span4Mux_v
    port map (
            O => \N__28615\,
            I => \N__28612\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__28612\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__5749\ : InMux
    port map (
            O => \N__28609\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__28606\,
            I => \N__28603\
        );

    \I__5747\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__28600\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \N__28594\
        );

    \I__5744\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28591\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__28591\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__5742\ : InMux
    port map (
            O => \N__28588\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__5741\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__28582\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__28579\,
            I => \N__28576\
        );

    \I__5738\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28573\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__28573\,
            I => \N__28570\
        );

    \I__5736\ : Odrv4
    port map (
            O => \N__28570\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__5735\ : InMux
    port map (
            O => \N__28567\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__28564\,
            I => \N__28560\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28552\
        );

    \I__5732\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28552\
        );

    \I__5731\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28552\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__28552\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__5728\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28543\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__28543\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__5726\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__28537\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__5724\ : InMux
    port map (
            O => \N__28534\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__5723\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28528\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__28528\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__5721\ : InMux
    port map (
            O => \N__28525\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__28522\,
            I => \N__28517\
        );

    \I__5719\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28512\
        );

    \I__5718\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28505\
        );

    \I__5717\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28505\
        );

    \I__5716\ : InMux
    port map (
            O => \N__28516\,
            I => \N__28505\
        );

    \I__5715\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28502\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__28512\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__28505\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__28502\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__28495\,
            I => \N__28492\
        );

    \I__5710\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__28486\,
            I => \N__28483\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__28483\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__5705\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__5703\ : Span4Mux_v
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__5702\ : Odrv4
    port map (
            O => \N__28468\,
            I => \POWERLED.mult1_un82_sum_i_8\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__28465\,
            I => \N__28462\
        );

    \I__5700\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28459\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__28459\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__5698\ : InMux
    port map (
            O => \N__28456\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__5697\ : InMux
    port map (
            O => \N__28453\,
            I => \N__28450\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__28450\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__5695\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28443\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__28446\,
            I => \N__28439\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__28443\,
            I => \N__28434\
        );

    \I__5692\ : InMux
    port map (
            O => \N__28442\,
            I => \N__28431\
        );

    \I__5691\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28426\
        );

    \I__5690\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28426\
        );

    \I__5689\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28423\
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__28434\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__28431\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__28426\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__28423\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__5684\ : InMux
    port map (
            O => \N__28414\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__28411\,
            I => \N__28407\
        );

    \I__5682\ : InMux
    port map (
            O => \N__28410\,
            I => \N__28399\
        );

    \I__5681\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28399\
        );

    \I__5680\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28399\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__28399\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__28396\,
            I => \N__28393\
        );

    \I__5677\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28390\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__28390\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__5675\ : InMux
    port map (
            O => \N__28387\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__5674\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28381\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__28381\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__5672\ : InMux
    port map (
            O => \N__28378\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__28375\,
            I => \POWERLED.mult1_un152_sum_s_8_cascade_\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__28372\,
            I => \N__28369\
        );

    \I__5669\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28366\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__28366\,
            I => \N__28363\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__28363\,
            I => \N__28360\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__28360\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__5665\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28354\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__28354\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__5663\ : InMux
    port map (
            O => \N__28351\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__5662\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28345\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__28345\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__5660\ : InMux
    port map (
            O => \N__28342\,
            I => \N__28339\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__28339\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__5658\ : InMux
    port map (
            O => \N__28336\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__5657\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__28330\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__5655\ : InMux
    port map (
            O => \N__28327\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__28324\,
            I => \N__28321\
        );

    \I__5653\ : InMux
    port map (
            O => \N__28321\,
            I => \N__28318\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__28318\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__5651\ : InMux
    port map (
            O => \N__28315\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__5650\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28309\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__28309\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__5648\ : InMux
    port map (
            O => \N__28306\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__28303\,
            I => \N__28300\
        );

    \I__5646\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__28297\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__5644\ : InMux
    port map (
            O => \N__28294\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__5643\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28288\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__28288\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__5641\ : InMux
    port map (
            O => \N__28285\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__5640\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28278\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__28281\,
            I => \N__28275\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__28278\,
            I => \N__28269\
        );

    \I__5637\ : InMux
    port map (
            O => \N__28275\,
            I => \N__28262\
        );

    \I__5636\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28262\
        );

    \I__5635\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28262\
        );

    \I__5634\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28259\
        );

    \I__5633\ : Odrv4
    port map (
            O => \N__28269\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__28262\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__28259\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__5630\ : CascadeMux
    port map (
            O => \N__28252\,
            I => \N__28248\
        );

    \I__5629\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28240\
        );

    \I__5628\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28240\
        );

    \I__5627\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28240\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__28240\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__5624\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28231\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__28228\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__5621\ : InMux
    port map (
            O => \N__28225\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__5620\ : InMux
    port map (
            O => \N__28222\,
            I => \N__28219\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__28219\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__5618\ : InMux
    port map (
            O => \N__28216\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__5617\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__5615\ : Span4Mux_h
    port map (
            O => \N__28207\,
            I => \N__28200\
        );

    \I__5614\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28191\
        );

    \I__5613\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28191\
        );

    \I__5612\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28191\
        );

    \I__5611\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28191\
        );

    \I__5610\ : Sp12to4
    port map (
            O => \N__28200\,
            I => \N__28186\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__28191\,
            I => \N__28186\
        );

    \I__5608\ : Span12Mux_v
    port map (
            O => \N__28186\,
            I => \N__28183\
        );

    \I__5607\ : Odrv12
    port map (
            O => \N__28183\,
            I => v33dsw_ok
        );

    \I__5606\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28172\
        );

    \I__5605\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28161\
        );

    \I__5604\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28161\
        );

    \I__5603\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28161\
        );

    \I__5602\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28161\
        );

    \I__5601\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28161\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__28172\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__28161\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__5598\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28148\
        );

    \I__5597\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28137\
        );

    \I__5596\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28137\
        );

    \I__5595\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28137\
        );

    \I__5594\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28137\
        );

    \I__5593\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28137\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__28148\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__28137\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__5590\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28129\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__28129\,
            I => \DSW_PWRGD.curr_state10\
        );

    \I__5588\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28123\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__28123\,
            I => \N__28120\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__28120\,
            I => \N__28117\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__28117\,
            I => vccst_cpu_ok
        );

    \I__5584\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28111\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__28111\,
            I => \N__28108\
        );

    \I__5582\ : Span4Mux_v
    port map (
            O => \N__28108\,
            I => \N__28105\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__28105\,
            I => v5s_ok
        );

    \I__5580\ : CascadeMux
    port map (
            O => \N__28102\,
            I => \N__28099\
        );

    \I__5579\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28096\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__28096\,
            I => \N__28093\
        );

    \I__5577\ : Span4Mux_v
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__5576\ : IoSpan4Mux
    port map (
            O => \N__28090\,
            I => \N__28087\
        );

    \I__5575\ : IoSpan4Mux
    port map (
            O => \N__28087\,
            I => \N__28084\
        );

    \I__5574\ : Odrv4
    port map (
            O => \N__28084\,
            I => v33s_ok
        );

    \I__5573\ : IoInMux
    port map (
            O => \N__28081\,
            I => \N__28078\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__28078\,
            I => \N__28075\
        );

    \I__5571\ : IoSpan4Mux
    port map (
            O => \N__28075\,
            I => \N__28072\
        );

    \I__5570\ : Span4Mux_s3_h
    port map (
            O => \N__28072\,
            I => \N__28069\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__28069\,
            I => \N__28065\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__28068\,
            I => \N__28061\
        );

    \I__5567\ : Span4Mux_v
    port map (
            O => \N__28065\,
            I => \N__28058\
        );

    \I__5566\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28055\
        );

    \I__5565\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28052\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__28058\,
            I => dsw_pwrok
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__28055\,
            I => dsw_pwrok
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__28052\,
            I => dsw_pwrok
        );

    \I__5561\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28038\
        );

    \I__5560\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28038\
        );

    \I__5559\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28035\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__28038\,
            I => \N__28030\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__28035\,
            I => \N__28027\
        );

    \I__5556\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28022\
        );

    \I__5555\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28022\
        );

    \I__5554\ : Span4Mux_v
    port map (
            O => \N__28030\,
            I => \N__28019\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__28027\,
            I => \N__28016\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__28022\,
            I => \N__28013\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__28019\,
            I => \N__28007\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__28007\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__28013\,
            I => \N__28004\
        );

    \I__5548\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28001\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__28007\,
            I => \N_392\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__28004\,
            I => \N_392\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__28001\,
            I => \N_392\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__27994\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\
        );

    \I__5543\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27984\
        );

    \I__5542\ : IoInMux
    port map (
            O => \N__27990\,
            I => \N__27977\
        );

    \I__5541\ : IoInMux
    port map (
            O => \N__27989\,
            I => \N__27974\
        );

    \I__5540\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27968\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__27987\,
            I => \N__27964\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27961\
        );

    \I__5537\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27952\
        );

    \I__5536\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27952\
        );

    \I__5535\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27952\
        );

    \I__5534\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27952\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__27977\,
            I => \N__27947\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__27974\,
            I => \N__27947\
        );

    \I__5531\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27939\
        );

    \I__5530\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27939\
        );

    \I__5529\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27939\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27936\
        );

    \I__5527\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27929\
        );

    \I__5526\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27926\
        );

    \I__5525\ : Span4Mux_h
    port map (
            O => \N__27961\,
            I => \N__27923\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__27952\,
            I => \N__27920\
        );

    \I__5523\ : IoSpan4Mux
    port map (
            O => \N__27947\,
            I => \N__27917\
        );

    \I__5522\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27914\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27911\
        );

    \I__5520\ : Span4Mux_v
    port map (
            O => \N__27936\,
            I => \N__27908\
        );

    \I__5519\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27899\
        );

    \I__5518\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27899\
        );

    \I__5517\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27899\
        );

    \I__5516\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27899\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27894\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27894\
        );

    \I__5513\ : Sp12to4
    port map (
            O => \N__27923\,
            I => \N__27889\
        );

    \I__5512\ : Span12Mux_s2_v
    port map (
            O => \N__27920\,
            I => \N__27889\
        );

    \I__5511\ : Span4Mux_s3_h
    port map (
            O => \N__27917\,
            I => \N__27882\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__27914\,
            I => \N__27882\
        );

    \I__5509\ : Span4Mux_s3_h
    port map (
            O => \N__27911\,
            I => \N__27882\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__27908\,
            I => \N__27875\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27875\
        );

    \I__5506\ : Span4Mux_h
    port map (
            O => \N__27894\,
            I => \N__27875\
        );

    \I__5505\ : Odrv12
    port map (
            O => \N__27889\,
            I => v5s_enn
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__27882\,
            I => v5s_enn
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__27875\,
            I => v5s_enn
        );

    \I__5502\ : IoInMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__5500\ : IoSpan4Mux
    port map (
            O => \N__27862\,
            I => \N__27859\
        );

    \I__5499\ : Sp12to4
    port map (
            O => \N__27859\,
            I => \N__27856\
        );

    \I__5498\ : Odrv12
    port map (
            O => \N__27856\,
            I => vccin_en
        );

    \I__5497\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27850\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__27850\,
            I => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0\
        );

    \I__5495\ : InMux
    port map (
            O => \N__27847\,
            I => \N__27819\
        );

    \I__5494\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27819\
        );

    \I__5493\ : InMux
    port map (
            O => \N__27845\,
            I => \N__27819\
        );

    \I__5492\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27819\
        );

    \I__5491\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27810\
        );

    \I__5490\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27810\
        );

    \I__5489\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27810\
        );

    \I__5488\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27810\
        );

    \I__5487\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27801\
        );

    \I__5486\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27801\
        );

    \I__5485\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27801\
        );

    \I__5484\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27801\
        );

    \I__5483\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27794\
        );

    \I__5482\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27794\
        );

    \I__5481\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27794\
        );

    \I__5480\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27789\
        );

    \I__5479\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27789\
        );

    \I__5478\ : InMux
    port map (
            O => \N__27830\,
            I => \N__27784\
        );

    \I__5477\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27784\
        );

    \I__5476\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27781\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27778\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__27810\,
            I => \N__27773\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__27801\,
            I => \N__27773\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__27794\,
            I => \N__27768\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27768\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27763\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27763\
        );

    \I__5468\ : Span4Mux_v
    port map (
            O => \N__27778\,
            I => \N__27756\
        );

    \I__5467\ : Span4Mux_v
    port map (
            O => \N__27773\,
            I => \N__27756\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__27768\,
            I => \N__27756\
        );

    \I__5465\ : Span12Mux_s9_v
    port map (
            O => \N__27763\,
            I => \N__27753\
        );

    \I__5464\ : Span4Mux_v
    port map (
            O => \N__27756\,
            I => \N__27750\
        );

    \I__5463\ : Odrv12
    port map (
            O => \N__27753\,
            I => \un4_counter_7_c_RNIBJDJ\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__27750\,
            I => \un4_counter_7_c_RNIBJDJ\
        );

    \I__5461\ : SRMux
    port map (
            O => \N__27745\,
            I => \N__27741\
        );

    \I__5460\ : SRMux
    port map (
            O => \N__27744\,
            I => \N__27738\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27734\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__27738\,
            I => \N__27731\
        );

    \I__5457\ : SRMux
    port map (
            O => \N__27737\,
            I => \N__27728\
        );

    \I__5456\ : Span4Mux_v
    port map (
            O => \N__27734\,
            I => \N__27724\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__27731\,
            I => \N__27721\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__27728\,
            I => \N__27718\
        );

    \I__5453\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27715\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__27724\,
            I => \un4_counter_7_c_RNI09TK5\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__27721\,
            I => \un4_counter_7_c_RNI09TK5\
        );

    \I__5450\ : Odrv12
    port map (
            O => \N__27718\,
            I => \un4_counter_7_c_RNI09TK5\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__27715\,
            I => \un4_counter_7_c_RNI09TK5\
        );

    \I__5448\ : CascadeMux
    port map (
            O => \N__27706\,
            I => \N__27703\
        );

    \I__5447\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27700\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__27700\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__5444\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27691\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__27691\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__5442\ : InMux
    port map (
            O => \N__27688\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__5441\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27679\
        );

    \I__5440\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27679\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__27679\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__5438\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27670\
        );

    \I__5437\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27670\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__27670\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__5435\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27664\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__27664\,
            I => \VPP_VDDQ.un29_clk_100khz_3\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__27661\,
            I => \N__27658\
        );

    \I__5432\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27655\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__27655\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__5430\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27649\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__27649\,
            I => \VPP_VDDQ.un29_clk_100khz_1\
        );

    \I__5428\ : CascadeMux
    port map (
            O => \N__27646\,
            I => \N__27643\
        );

    \I__5427\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27636\
        );

    \I__5426\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27636\
        );

    \I__5425\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27633\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27630\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__27633\,
            I => \N__27627\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__27630\,
            I => \N__27624\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__27627\,
            I => \N__27621\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__27624\,
            I => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__27621\,
            I => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__27616\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_\
        );

    \I__5417\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27607\
        );

    \I__5416\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27607\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__27607\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__5414\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27601\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__27601\,
            I => \VPP_VDDQ.count_2_0_6\
        );

    \I__5412\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27595\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__27595\,
            I => \VPP_VDDQ.count_3_13\
        );

    \I__5410\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27588\
        );

    \I__5409\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27585\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27582\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__27585\,
            I => \VPP_VDDQ.count_rst_2\
        );

    \I__5406\ : Odrv4
    port map (
            O => \N__27582\,
            I => \VPP_VDDQ.count_rst_2\
        );

    \I__5405\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27574\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27570\
        );

    \I__5403\ : InMux
    port map (
            O => \N__27573\,
            I => \N__27567\
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__27570\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__27567\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__5400\ : CEMux
    port map (
            O => \N__27562\,
            I => \N__27555\
        );

    \I__5399\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27548\
        );

    \I__5398\ : CEMux
    port map (
            O => \N__27560\,
            I => \N__27548\
        );

    \I__5397\ : CEMux
    port map (
            O => \N__27559\,
            I => \N__27545\
        );

    \I__5396\ : CEMux
    port map (
            O => \N__27558\,
            I => \N__27542\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__27555\,
            I => \N__27539\
        );

    \I__5394\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27534\
        );

    \I__5393\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27534\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__27548\,
            I => \N__27522\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27514\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27514\
        );

    \I__5389\ : Span4Mux_s2_v
    port map (
            O => \N__27539\,
            I => \N__27511\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__27534\,
            I => \N__27508\
        );

    \I__5387\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27499\
        );

    \I__5386\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27499\
        );

    \I__5385\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27499\
        );

    \I__5384\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27499\
        );

    \I__5383\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27490\
        );

    \I__5382\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27490\
        );

    \I__5381\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27490\
        );

    \I__5380\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27490\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__27525\,
            I => \N__27485\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__27522\,
            I => \N__27481\
        );

    \I__5377\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27474\
        );

    \I__5376\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27474\
        );

    \I__5375\ : CEMux
    port map (
            O => \N__27519\,
            I => \N__27474\
        );

    \I__5374\ : Span4Mux_s2_v
    port map (
            O => \N__27514\,
            I => \N__27471\
        );

    \I__5373\ : Span4Mux_s2_h
    port map (
            O => \N__27511\,
            I => \N__27466\
        );

    \I__5372\ : Span4Mux_s2_v
    port map (
            O => \N__27508\,
            I => \N__27466\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__27499\,
            I => \N__27461\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27461\
        );

    \I__5369\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27454\
        );

    \I__5368\ : CEMux
    port map (
            O => \N__27488\,
            I => \N__27454\
        );

    \I__5367\ : InMux
    port map (
            O => \N__27485\,
            I => \N__27454\
        );

    \I__5366\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27451\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__27481\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__27474\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__27471\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5362\ : Odrv4
    port map (
            O => \N__27466\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__27461\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__27454\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__27451\,
            I => \VPP_VDDQ.count_en\
        );

    \I__5358\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27433\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__27433\,
            I => \VPP_VDDQ.count_3_14\
        );

    \I__5356\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27426\
        );

    \I__5355\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27423\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__27426\,
            I => \N__27420\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__27423\,
            I => \VPP_VDDQ.count_rst_3\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__27420\,
            I => \VPP_VDDQ.count_rst_3\
        );

    \I__5351\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27411\
        );

    \I__5350\ : CascadeMux
    port map (
            O => \N__27414\,
            I => \N__27408\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27405\
        );

    \I__5348\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27402\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__27405\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__27402\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__5345\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27393\
        );

    \I__5344\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27390\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__27393\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__27390\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__27385\,
            I => \VPP_VDDQ.un29_clk_100khz_0_cascade_\
        );

    \I__5340\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27379\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__27379\,
            I => \VPP_VDDQ.un29_clk_100khz_2\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__27376\,
            I => \N__27372\
        );

    \I__5337\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27369\
        );

    \I__5336\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27366\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__27369\,
            I => \N__27361\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__27366\,
            I => \N__27361\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__27361\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__5332\ : CascadeMux
    port map (
            O => \N__27358\,
            I => \POWERLED.dutycycle_en_12_cascade_\
        );

    \I__5331\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27351\
        );

    \I__5330\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27348\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__27351\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__27348\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__5327\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27339\
        );

    \I__5326\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27336\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__27339\,
            I => \N__27333\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__27336\,
            I => \N__27330\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__27333\,
            I => \VPP_VDDQ.count_rst_1\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__27330\,
            I => \VPP_VDDQ.count_rst_1\
        );

    \I__5321\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27322\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27319\
        );

    \I__5319\ : Odrv12
    port map (
            O => \N__27319\,
            I => \VPP_VDDQ.count_3_12\
        );

    \I__5318\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27312\
        );

    \I__5317\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27309\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__27312\,
            I => \VPP_VDDQ.count_rst_12\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__27309\,
            I => \VPP_VDDQ.count_rst_12\
        );

    \I__5314\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27301\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__27301\,
            I => \VPP_VDDQ.count_3_7\
        );

    \I__5312\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27295\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__27295\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__27292\,
            I => \POWERLED.dutycycleZ0Z_7_cascade_\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__27289\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_7_cascade_\
        );

    \I__5308\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27280\
        );

    \I__5307\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27280\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__27280\,
            I => \N__27277\
        );

    \I__5305\ : Span4Mux_h
    port map (
            O => \N__27277\,
            I => \N__27274\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__27274\,
            I => \POWERLED.dutycycle_en_11\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__27271\,
            I => \POWERLED.N_156_N_cascade_\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__27268\,
            I => \N__27265\
        );

    \I__5301\ : InMux
    port map (
            O => \N__27265\,
            I => \N__27262\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__27262\,
            I => \POWERLED.N_158_N\
        );

    \I__5299\ : InMux
    port map (
            O => \N__27259\,
            I => \N__27249\
        );

    \I__5298\ : InMux
    port map (
            O => \N__27258\,
            I => \N__27249\
        );

    \I__5297\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27249\
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__27256\,
            I => \N__27242\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__27249\,
            I => \N__27238\
        );

    \I__5294\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27235\
        );

    \I__5293\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27230\
        );

    \I__5292\ : InMux
    port map (
            O => \N__27246\,
            I => \N__27230\
        );

    \I__5291\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27223\
        );

    \I__5290\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27223\
        );

    \I__5289\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27223\
        );

    \I__5288\ : Span4Mux_h
    port map (
            O => \N__27238\,
            I => \N__27218\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__27235\,
            I => \N__27218\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__27230\,
            I => \N__27213\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__27223\,
            I => \N__27213\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__27218\,
            I => \N__27210\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__27213\,
            I => \N__27207\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__27210\,
            I => \POWERLED.func_state_RNIHU7V2Z0Z_0\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__27207\,
            I => \POWERLED.func_state_RNIHU7V2Z0Z_0\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__27202\,
            I => \POWERLED.dutycycleZ0Z_13_cascade_\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__27199\,
            I => \POWERLED.N_161_N_cascade_\
        );

    \I__5278\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__27193\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__5275\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27179\
        );

    \I__5274\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27179\
        );

    \I__5273\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27176\
        );

    \I__5272\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27173\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27170\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__27176\,
            I => \N__27165\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__27173\,
            I => \N__27165\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__27170\,
            I => \N__27162\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__27165\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_0\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__27162\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_0\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__27157\,
            I => \POWERLED.N_361_cascade_\
        );

    \I__5264\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27148\
        );

    \I__5263\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27148\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__27148\,
            I => \POWERLED.dutycycle_RNI_9Z0Z_3\
        );

    \I__5261\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__27142\,
            I => \POWERLED.N_361\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__5258\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27130\
        );

    \I__5257\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27130\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__27130\,
            I => \N__27127\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__27127\,
            I => \POWERLED.N_369\
        );

    \I__5254\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27121\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__27121\,
            I => \POWERLED.d_i3_mux\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__27118\,
            I => \POWERLED.un1_i3_mux_cascade_\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__27115\,
            I => \N__27112\
        );

    \I__5250\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27106\
        );

    \I__5249\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27106\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__27106\,
            I => \N__27103\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__27103\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__27100\,
            I => \N__27096\
        );

    \I__5245\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27091\
        );

    \I__5244\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27091\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__27091\,
            I => \POWERLED.dutycycleZ1Z_3\
        );

    \I__5242\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27082\
        );

    \I__5241\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27082\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__27082\,
            I => \POWERLED.dutycycle_RNIQU4T5Z0Z_3\
        );

    \I__5239\ : CascadeMux
    port map (
            O => \N__27079\,
            I => \POWERLED.un1_dutycycle_172_m1_1_cascade_\
        );

    \I__5238\ : InMux
    port map (
            O => \N__27076\,
            I => \N__27073\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__27073\,
            I => \POWERLED.un1_dutycycle_172_m1\
        );

    \I__5236\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27064\
        );

    \I__5235\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27057\
        );

    \I__5234\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27057\
        );

    \I__5233\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27057\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__27064\,
            I => \N__27045\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__27057\,
            I => \N__27045\
        );

    \I__5230\ : InMux
    port map (
            O => \N__27056\,
            I => \N__27042\
        );

    \I__5229\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27039\
        );

    \I__5228\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27036\
        );

    \I__5227\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27027\
        );

    \I__5226\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27027\
        );

    \I__5225\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27027\
        );

    \I__5224\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27024\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__27045\,
            I => \N__27019\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__27042\,
            I => \N__27019\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27014\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__27036\,
            I => \N__27014\
        );

    \I__5219\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27006\
        );

    \I__5218\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27006\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27003\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__26996\
        );

    \I__5215\ : Span4Mux_h
    port map (
            O => \N__27019\,
            I => \N__26996\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__27014\,
            I => \N__26996\
        );

    \I__5213\ : InMux
    port map (
            O => \N__27013\,
            I => \N__26989\
        );

    \I__5212\ : InMux
    port map (
            O => \N__27012\,
            I => \N__26989\
        );

    \I__5211\ : InMux
    port map (
            O => \N__27011\,
            I => \N__26989\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__27006\,
            I => \POWERLED.N_2905_i\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__27003\,
            I => \POWERLED.N_2905_i\
        );

    \I__5208\ : Odrv4
    port map (
            O => \N__26996\,
            I => \POWERLED.N_2905_i\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__26989\,
            I => \POWERLED.N_2905_i\
        );

    \I__5206\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26971\
        );

    \I__5205\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26971\
        );

    \I__5204\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26964\
        );

    \I__5203\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26964\
        );

    \I__5202\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26961\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__26971\,
            I => \N__26958\
        );

    \I__5200\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26953\
        );

    \I__5199\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26953\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__26964\,
            I => \N__26950\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__26961\,
            I => \N__26947\
        );

    \I__5196\ : Span4Mux_h
    port map (
            O => \N__26958\,
            I => \N__26940\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26940\
        );

    \I__5194\ : Span4Mux_s3_v
    port map (
            O => \N__26950\,
            I => \N__26940\
        );

    \I__5193\ : Odrv12
    port map (
            O => \N__26947\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__26940\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__5191\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26932\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__26932\,
            I => \N__26928\
        );

    \I__5189\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26925\
        );

    \I__5188\ : Span4Mux_s3_v
    port map (
            O => \N__26928\,
            I => \N__26920\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__26925\,
            I => \N__26920\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__26920\,
            I => \POWERLED.N_19\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__26917\,
            I => \POWERLED.N_134_cascade_\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__5183\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__26908\,
            I => \POWERLED.un1_dutycycle_172_m0\
        );

    \I__5181\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26902\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__26902\,
            I => \N__26897\
        );

    \I__5179\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26892\
        );

    \I__5178\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26892\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__26897\,
            I => \POWERLED.g2_0_1_0\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__26892\,
            I => \POWERLED.g2_0_1_0\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__26887\,
            I => \POWERLED.un1_dutycycle_172_m0_cascade_\
        );

    \I__5174\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26880\
        );

    \I__5173\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26877\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__26880\,
            I => \POWERLED.N_15\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__26877\,
            I => \POWERLED.N_15\
        );

    \I__5170\ : InMux
    port map (
            O => \N__26872\,
            I => \N__26869\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__26869\,
            I => \POWERLED.N_10\
        );

    \I__5168\ : CascadeMux
    port map (
            O => \N__26866\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_\
        );

    \I__5167\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26860\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__26860\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_6\
        );

    \I__5165\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26850\
        );

    \I__5164\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26850\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__26855\,
            I => \N__26846\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26843\
        );

    \I__5161\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26840\
        );

    \I__5160\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26837\
        );

    \I__5159\ : Span4Mux_s3_v
    port map (
            O => \N__26843\,
            I => \N__26834\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26827\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__26837\,
            I => \N__26827\
        );

    \I__5156\ : Span4Mux_s3_h
    port map (
            O => \N__26834\,
            I => \N__26827\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__26827\,
            I => \tmp_1_rep1_RNI\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__26824\,
            I => \POWERLED.dutycycle_RNIZ0Z_1_cascade_\
        );

    \I__5153\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26814\
        );

    \I__5152\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26811\
        );

    \I__5151\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26806\
        );

    \I__5150\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26806\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__26817\,
            I => \N__26802\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__26814\,
            I => \N__26799\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__26811\,
            I => \N__26796\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__26806\,
            I => \N__26793\
        );

    \I__5145\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26788\
        );

    \I__5144\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26788\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__26799\,
            I => \N__26785\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__26796\,
            I => \N__26780\
        );

    \I__5141\ : Span4Mux_v
    port map (
            O => \N__26793\,
            I => \N__26780\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__26788\,
            I => \N__26777\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__26785\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__26780\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__26777\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__26770\,
            I => \N__26767\
        );

    \I__5135\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26764\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__26764\,
            I => \N__26761\
        );

    \I__5133\ : Odrv4
    port map (
            O => \N__26761\,
            I => \POWERLED.mult1_un75_sum_i_8\
        );

    \I__5132\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26755\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__26755\,
            I => \N__26752\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__26752\,
            I => \POWERLED.N_96_mux_i_i_2_1\
        );

    \I__5129\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26743\
        );

    \I__5128\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26743\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__26743\,
            I => \N__26740\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__26740\,
            I => \N_96_mux_i_i_2\
        );

    \I__5125\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26731\
        );

    \I__5124\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26731\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26728\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__26728\,
            I => \N_13\
        );

    \I__5121\ : CascadeMux
    port map (
            O => \N__26725\,
            I => \N__26722\
        );

    \I__5120\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26719\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26716\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__26716\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__26713\,
            I => \N__26710\
        );

    \I__5116\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26699\
        );

    \I__5115\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26699\
        );

    \I__5114\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26699\
        );

    \I__5113\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26696\
        );

    \I__5112\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26693\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__26699\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__26696\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__26693\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__26686\,
            I => \N__26683\
        );

    \I__5107\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26680\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__26677\,
            I => \N__26674\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__26674\,
            I => \POWERLED.mult1_un110_sum_i_8\
        );

    \I__5103\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26667\
        );

    \I__5102\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26664\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__26667\,
            I => \POWERLED.count_off_1_sqmuxa\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__26664\,
            I => \POWERLED.count_off_1_sqmuxa\
        );

    \I__5099\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26653\
        );

    \I__5098\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26653\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__26653\,
            I => \POWERLED.un1_dutycycle_172_m4\
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__26650\,
            I => \N__26647\
        );

    \I__5095\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26644\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26641\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__26641\,
            I => \POWERLED.mult1_un96_sum_i_8\
        );

    \I__5092\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26634\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__26637\,
            I => \N__26630\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__26634\,
            I => \N__26627\
        );

    \I__5089\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26624\
        );

    \I__5088\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26621\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__26627\,
            I => \N__26616\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26616\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__26621\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__26616\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__5083\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__26608\,
            I => \POWERLED.N_6117_i\
        );

    \I__5081\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26601\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__26604\,
            I => \N__26597\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__26601\,
            I => \N__26594\
        );

    \I__5078\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26591\
        );

    \I__5077\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26588\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__26594\,
            I => \N__26583\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26583\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__26588\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__26583\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__5072\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26575\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__26575\,
            I => \POWERLED.N_6118_i\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__26572\,
            I => \N__26569\
        );

    \I__5069\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26565\
        );

    \I__5068\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26562\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26559\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__26562\,
            I => \N__26555\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__26559\,
            I => \N__26552\
        );

    \I__5064\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26549\
        );

    \I__5063\ : Span4Mux_v
    port map (
            O => \N__26555\,
            I => \N__26546\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__26552\,
            I => \N__26541\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26541\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__26546\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__26541\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__5058\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26533\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__26533\,
            I => \POWERLED.N_6119_i\
        );

    \I__5056\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26526\
        );

    \I__5055\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26522\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__26526\,
            I => \N__26519\
        );

    \I__5053\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26516\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__26522\,
            I => \N__26513\
        );

    \I__5051\ : Span12Mux_s7_h
    port map (
            O => \N__26519\,
            I => \N__26508\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__26516\,
            I => \N__26508\
        );

    \I__5049\ : Odrv4
    port map (
            O => \N__26513\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__5048\ : Odrv12
    port map (
            O => \N__26508\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__5047\ : InMux
    port map (
            O => \N__26503\,
            I => \N__26500\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__26500\,
            I => \POWERLED.N_6120_i\
        );

    \I__5045\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26494\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26490\
        );

    \I__5043\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26486\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__26490\,
            I => \N__26483\
        );

    \I__5041\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26480\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26477\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__26483\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__26480\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__26477\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__5036\ : InMux
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__26467\,
            I => \POWERLED.N_6121_i\
        );

    \I__5034\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26461\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26458\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__26458\,
            I => \N__26453\
        );

    \I__5031\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26450\
        );

    \I__5030\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26447\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__26453\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__26450\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__26447\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__5026\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26437\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__26437\,
            I => \POWERLED.N_6122_i\
        );

    \I__5024\ : InMux
    port map (
            O => \N__26434\,
            I => \bfn_8_12_0_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26428\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__26428\,
            I => \N__26425\
        );

    \I__5021\ : Span12Mux_s7_h
    port map (
            O => \N__26425\,
            I => \N__26422\
        );

    \I__5020\ : Odrv12
    port map (
            O => \N__26422\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__26419\,
            I => \N__26416\
        );

    \I__5018\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26413\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26410\
        );

    \I__5016\ : Odrv12
    port map (
            O => \N__26410\,
            I => \POWERLED.un85_clk_100khz_3\
        );

    \I__5015\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26404\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26400\
        );

    \I__5013\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26397\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__26400\,
            I => \N__26393\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__26397\,
            I => \N__26390\
        );

    \I__5010\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26387\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__26393\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__26390\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__26387\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__5006\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26377\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__26377\,
            I => \POWERLED.N_6110_i\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__26374\,
            I => \N__26371\
        );

    \I__5003\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26368\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__26368\,
            I => \POWERLED.un85_clk_100khz_4\
        );

    \I__5001\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26362\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__26362\,
            I => \N__26359\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__26359\,
            I => \N__26354\
        );

    \I__4998\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26351\
        );

    \I__4997\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26348\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__26354\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__26351\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__26348\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__4993\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__26338\,
            I => \POWERLED.N_6111_i\
        );

    \I__4991\ : CascadeMux
    port map (
            O => \N__26335\,
            I => \N__26332\
        );

    \I__4990\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26329\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__26326\,
            I => \POWERLED.mult1_un131_sum_i_8\
        );

    \I__4987\ : InMux
    port map (
            O => \N__26323\,
            I => \N__26320\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__26320\,
            I => \N__26316\
        );

    \I__4985\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26312\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__26316\,
            I => \N__26309\
        );

    \I__4983\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26306\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__26312\,
            I => \N__26303\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__26309\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__26306\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__26303\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__4978\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26293\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__26293\,
            I => \POWERLED.N_6112_i\
        );

    \I__4976\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26287\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26284\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__26284\,
            I => \N__26279\
        );

    \I__4973\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26276\
        );

    \I__4972\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26273\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__26279\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__26276\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__26273\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__4968\ : CascadeMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__4967\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26260\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__26257\,
            I => \POWERLED.mult1_un124_sum_i_8\
        );

    \I__4964\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__26251\,
            I => \POWERLED.N_6113_i\
        );

    \I__4962\ : InMux
    port map (
            O => \N__26248\,
            I => \N__26245\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__26245\,
            I => \N__26242\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__26242\,
            I => \N__26237\
        );

    \I__4959\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26234\
        );

    \I__4958\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26231\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__26237\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__26234\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__26231\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__26224\,
            I => \N__26221\
        );

    \I__4953\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26218\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__26218\,
            I => \POWERLED.mult1_un117_sum_i_8\
        );

    \I__4951\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26212\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__26212\,
            I => \POWERLED.N_6114_i\
        );

    \I__4949\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26206\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__26206\,
            I => \N__26203\
        );

    \I__4947\ : Span4Mux_h
    port map (
            O => \N__26203\,
            I => \N__26198\
        );

    \I__4946\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26195\
        );

    \I__4945\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26192\
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__26198\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__26195\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__26192\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__4941\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__26182\,
            I => \POWERLED.N_6115_i\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__26179\,
            I => \N__26176\
        );

    \I__4938\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26173\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__26173\,
            I => \N__26170\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__26170\,
            I => \N__26167\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__26167\,
            I => \POWERLED.mult1_un103_sum_i_8\
        );

    \I__4934\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26161\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26158\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__26158\,
            I => \N__26153\
        );

    \I__4931\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26150\
        );

    \I__4930\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26147\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__26153\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__26150\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__26147\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__4926\ : InMux
    port map (
            O => \N__26140\,
            I => \N__26137\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__26137\,
            I => \POWERLED.N_6116_i\
        );

    \I__4924\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26127\
        );

    \I__4923\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26127\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__26132\,
            I => \N__26123\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__26127\,
            I => \N__26120\
        );

    \I__4920\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26115\
        );

    \I__4919\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26115\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__26120\,
            I => \N__26111\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26108\
        );

    \I__4916\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26105\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__26111\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__4914\ : Odrv12
    port map (
            O => \N__26108\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__26105\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__26098\,
            I => \N__26094\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__26097\,
            I => \N__26090\
        );

    \I__4910\ : InMux
    port map (
            O => \N__26094\,
            I => \N__26083\
        );

    \I__4909\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26083\
        );

    \I__4908\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26083\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__26083\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__26080\,
            I => \N__26077\
        );

    \I__4905\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26074\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__26074\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__26071\,
            I => \N__26067\
        );

    \I__4902\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26062\
        );

    \I__4901\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26062\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26056\
        );

    \I__4899\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26053\
        );

    \I__4898\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26050\
        );

    \I__4897\ : InMux
    port map (
            O => \N__26059\,
            I => \N__26047\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__26056\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__26053\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__26050\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__26047\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__4891\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26032\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__26029\,
            I => \POWERLED.un85_clk_100khz_0\
        );

    \I__4888\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26023\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__26023\,
            I => \N__26019\
        );

    \I__4886\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26013\
        );

    \I__4885\ : Span4Mux_v
    port map (
            O => \N__26019\,
            I => \N__26010\
        );

    \I__4884\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26003\
        );

    \I__4883\ : InMux
    port map (
            O => \N__26017\,
            I => \N__26003\
        );

    \I__4882\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26003\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__26013\,
            I => \N__26000\
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__26010\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__26003\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__26000\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__4877\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__25990\,
            I => \POWERLED.un1_count_cry_0_i\
        );

    \I__4875\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25984\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25980\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__25983\,
            I => \N__25977\
        );

    \I__4872\ : Span4Mux_v
    port map (
            O => \N__25980\,
            I => \N__25973\
        );

    \I__4871\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25970\
        );

    \I__4870\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25967\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__25973\,
            I => \N__25962\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__25970\,
            I => \N__25962\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__25967\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__25962\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__25957\,
            I => \N__25954\
        );

    \I__4864\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25951\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__25951\,
            I => \N__25948\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__25948\,
            I => \POWERLED.un85_clk_100khz_1\
        );

    \I__4861\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25942\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__25942\,
            I => \POWERLED.N_6108_i\
        );

    \I__4859\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25936\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__25936\,
            I => \N__25931\
        );

    \I__4857\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25928\
        );

    \I__4856\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25925\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__25931\,
            I => \N__25922\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__25928\,
            I => \N__25917\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__25925\,
            I => \N__25917\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__25922\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__25917\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__4850\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25909\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__25909\,
            I => \POWERLED.N_6109_i\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \N__25903\
        );

    \I__4847\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25900\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25897\
        );

    \I__4845\ : Odrv12
    port map (
            O => \N__25897\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__25894\,
            I => \N__25890\
        );

    \I__4843\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25882\
        );

    \I__4842\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25882\
        );

    \I__4841\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25882\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__25882\,
            I => \G_2898\
        );

    \I__4839\ : InMux
    port map (
            O => \N__25879\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__25876\,
            I => \N__25872\
        );

    \I__4837\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25867\
        );

    \I__4836\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25862\
        );

    \I__4835\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25862\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__25870\,
            I => \N__25859\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__25867\,
            I => \N__25855\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25852\
        );

    \I__4831\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25847\
        );

    \I__4830\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25847\
        );

    \I__4829\ : Span4Mux_v
    port map (
            O => \N__25855\,
            I => \N__25842\
        );

    \I__4828\ : Span4Mux_v
    port map (
            O => \N__25852\,
            I => \N__25842\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__25847\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__25842\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__4825\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__25834\,
            I => \N__25831\
        );

    \I__4823\ : Odrv12
    port map (
            O => \N__25831\,
            I => \POWERLED.curr_state_3_0\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__4821\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25822\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__25822\,
            I => \N__25819\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__25819\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__4818\ : InMux
    port map (
            O => \N__25816\,
            I => \POWERLED.mult1_un138_sum_cry_5_c\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__25813\,
            I => \N__25810\
        );

    \I__4816\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25807\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__25807\,
            I => \N__25804\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__25804\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__4813\ : InMux
    port map (
            O => \N__25801\,
            I => \POWERLED.mult1_un138_sum_cry_6_c\
        );

    \I__4812\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25795\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__25795\,
            I => \N__25792\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__25792\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__4809\ : InMux
    port map (
            O => \N__25789\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__4808\ : CEMux
    port map (
            O => \N__25786\,
            I => \N__25783\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__25783\,
            I => \N__25780\
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__25780\,
            I => \DSW_PWRGD.N_22_0\
        );

    \I__4805\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25773\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__25776\,
            I => \N__25770\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25766\
        );

    \I__4802\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25761\
        );

    \I__4801\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25761\
        );

    \I__4800\ : Span4Mux_h
    port map (
            O => \N__25766\,
            I => \N__25757\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__25761\,
            I => \N__25740\
        );

    \I__4798\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25737\
        );

    \I__4797\ : Span4Mux_h
    port map (
            O => \N__25757\,
            I => \N__25734\
        );

    \I__4796\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25727\
        );

    \I__4795\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25727\
        );

    \I__4794\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25727\
        );

    \I__4793\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25718\
        );

    \I__4792\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25718\
        );

    \I__4791\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25718\
        );

    \I__4790\ : InMux
    port map (
            O => \N__25750\,
            I => \N__25718\
        );

    \I__4789\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25711\
        );

    \I__4788\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25711\
        );

    \I__4787\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25711\
        );

    \I__4786\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25702\
        );

    \I__4785\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25702\
        );

    \I__4784\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25702\
        );

    \I__4783\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25702\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__25740\,
            I => \N__25699\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__25737\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__25734\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__25727\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__25718\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__25711\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__25702\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__25699\,
            I => \POWERLED.func_state_RNI1E8A4_0_0\
        );

    \I__4774\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25681\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__25681\,
            I => \N__25677\
        );

    \I__4772\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25672\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__25677\,
            I => \N__25669\
        );

    \I__4770\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25662\
        );

    \I__4769\ : InMux
    port map (
            O => \N__25675\,
            I => \N__25662\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__25672\,
            I => \N__25657\
        );

    \I__4767\ : Span4Mux_h
    port map (
            O => \N__25669\,
            I => \N__25657\
        );

    \I__4766\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25654\
        );

    \I__4765\ : InMux
    port map (
            O => \N__25667\,
            I => \N__25651\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__25662\,
            I => \N__25648\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__25657\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__25654\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__25651\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__25648\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4759\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25636\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25633\
        );

    \I__4757\ : Span4Mux_s3_h
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__25630\,
            I => \N__25627\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__25627\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__4754\ : CEMux
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25614\
        );

    \I__4752\ : CEMux
    port map (
            O => \N__25620\,
            I => \N__25611\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__25619\,
            I => \N__25608\
        );

    \I__4750\ : CEMux
    port map (
            O => \N__25618\,
            I => \N__25605\
        );

    \I__4749\ : CEMux
    port map (
            O => \N__25617\,
            I => \N__25602\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__25614\,
            I => \N__25599\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__25611\,
            I => \N__25596\
        );

    \I__4746\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25593\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__25605\,
            I => \N__25574\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__25602\,
            I => \N__25574\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__25599\,
            I => \N__25571\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__25596\,
            I => \N__25564\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__25593\,
            I => \N__25561\
        );

    \I__4740\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25554\
        );

    \I__4739\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25554\
        );

    \I__4738\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25554\
        );

    \I__4737\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25545\
        );

    \I__4736\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25545\
        );

    \I__4735\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25545\
        );

    \I__4734\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25545\
        );

    \I__4733\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25536\
        );

    \I__4732\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25536\
        );

    \I__4731\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25536\
        );

    \I__4730\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25536\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__25581\,
            I => \N__25533\
        );

    \I__4728\ : CEMux
    port map (
            O => \N__25580\,
            I => \N__25530\
        );

    \I__4727\ : CEMux
    port map (
            O => \N__25579\,
            I => \N__25527\
        );

    \I__4726\ : Sp12to4
    port map (
            O => \N__25574\,
            I => \N__25524\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__25571\,
            I => \N__25521\
        );

    \I__4724\ : CEMux
    port map (
            O => \N__25570\,
            I => \N__25512\
        );

    \I__4723\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25512\
        );

    \I__4722\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25512\
        );

    \I__4721\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25512\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__25564\,
            I => \N__25503\
        );

    \I__4719\ : Span4Mux_s1_h
    port map (
            O => \N__25561\,
            I => \N__25503\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__25554\,
            I => \N__25503\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__25545\,
            I => \N__25503\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__25536\,
            I => \N__25500\
        );

    \I__4715\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25497\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__25530\,
            I => \POWERLED.count_clk_en\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__25527\,
            I => \POWERLED.count_clk_en\
        );

    \I__4712\ : Odrv12
    port map (
            O => \N__25524\,
            I => \POWERLED.count_clk_en\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__25521\,
            I => \POWERLED.count_clk_en\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__25512\,
            I => \POWERLED.count_clk_en\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__25503\,
            I => \POWERLED.count_clk_en\
        );

    \I__4708\ : Odrv12
    port map (
            O => \N__25500\,
            I => \POWERLED.count_clk_en\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__25497\,
            I => \POWERLED.count_clk_en\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__25480\,
            I => \N__25476\
        );

    \I__4705\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25468\
        );

    \I__4704\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25468\
        );

    \I__4703\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25468\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__25468\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__25465\,
            I => \DSW_PWRGD.i3_mux_0_cascade_\
        );

    \I__4700\ : CascadeMux
    port map (
            O => \N__25462\,
            I => \N__25457\
        );

    \I__4699\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25454\
        );

    \I__4698\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25449\
        );

    \I__4697\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25449\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__25454\,
            I => \N__25444\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25444\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__25444\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__25441\,
            I => \DSW_PWRGD.N_6_cascade_\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__25438\,
            I => \N__25434\
        );

    \I__4691\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25431\
        );

    \I__4690\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25428\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__25431\,
            I => \DSW_PWRGD.un1_curr_state10_0\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__25428\,
            I => \DSW_PWRGD.un1_curr_state10_0\
        );

    \I__4687\ : InMux
    port map (
            O => \N__25423\,
            I => \POWERLED.mult1_un138_sum_cry_2_c\
        );

    \I__4686\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25417\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__25417\,
            I => \N__25414\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__25414\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__4683\ : InMux
    port map (
            O => \N__25411\,
            I => \POWERLED.mult1_un138_sum_cry_3_c\
        );

    \I__4682\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__25405\,
            I => \N__25402\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__25402\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__4679\ : InMux
    port map (
            O => \N__25399\,
            I => \POWERLED.mult1_un138_sum_cry_4_c\
        );

    \I__4678\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25392\
        );

    \I__4677\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25389\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__25392\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__25389\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__4674\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25378\
        );

    \I__4673\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25378\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__25378\,
            I => \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6CZ0\
        );

    \I__4671\ : InMux
    port map (
            O => \N__25375\,
            I => \VPP_VDDQ.un4_count_1_cry_10\
        );

    \I__4670\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25368\
        );

    \I__4669\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25365\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__25368\,
            I => \N__25362\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__25365\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__4666\ : Odrv4
    port map (
            O => \N__25362\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__4665\ : InMux
    port map (
            O => \N__25357\,
            I => \VPP_VDDQ.un4_count_1_cry_11\
        );

    \I__4664\ : InMux
    port map (
            O => \N__25354\,
            I => \VPP_VDDQ.un4_count_1_cry_12\
        );

    \I__4663\ : InMux
    port map (
            O => \N__25351\,
            I => \VPP_VDDQ.un4_count_1_cry_13\
        );

    \I__4662\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25345\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25341\
        );

    \I__4660\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25338\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__25341\,
            I => \N__25335\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__25338\,
            I => \N__25332\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__25335\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__4656\ : Odrv12
    port map (
            O => \N__25332\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__4655\ : InMux
    port map (
            O => \N__25327\,
            I => \VPP_VDDQ.un4_count_1_cry_14\
        );

    \I__4654\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25318\
        );

    \I__4653\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25318\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__25318\,
            I => \N__25315\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__25315\,
            I => \N__25312\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__25312\,
            I => \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0\
        );

    \I__4649\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25305\
        );

    \I__4648\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25302\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__25305\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__25302\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__4645\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25293\
        );

    \I__4644\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25290\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__25293\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__25290\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__25285\,
            I => \N__25281\
        );

    \I__4640\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25278\
        );

    \I__4639\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25275\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__25278\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__25275\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__4636\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25266\
        );

    \I__4635\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25263\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__25266\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__25263\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__4632\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25255\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__25252\,
            I => \DSW_PWRGD.un4_count_9\
        );

    \I__4629\ : IoInMux
    port map (
            O => \N__25249\,
            I => \N__25246\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__25246\,
            I => \N__25243\
        );

    \I__4627\ : IoSpan4Mux
    port map (
            O => \N__25243\,
            I => \N__25240\
        );

    \I__4626\ : Span4Mux_s1_h
    port map (
            O => \N__25240\,
            I => \N__25236\
        );

    \I__4625\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25233\
        );

    \I__4624\ : Span4Mux_h
    port map (
            O => \N__25236\,
            I => \N__25227\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__25233\,
            I => \N__25227\
        );

    \I__4622\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25224\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__25227\,
            I => \N__25221\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__25224\,
            I => \N__25218\
        );

    \I__4619\ : Span4Mux_v
    port map (
            O => \N__25221\,
            I => \N__25215\
        );

    \I__4618\ : Span12Mux_v
    port map (
            O => \N__25218\,
            I => \N__25212\
        );

    \I__4617\ : Span4Mux_h
    port map (
            O => \N__25215\,
            I => \N__25209\
        );

    \I__4616\ : Odrv12
    port map (
            O => \N__25212\,
            I => v33a_ok
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__25209\,
            I => v33a_ok
        );

    \I__4614\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25201\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25198\
        );

    \I__4612\ : Odrv12
    port map (
            O => \N__25198\,
            I => v5a_ok
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__25195\,
            I => \N__25191\
        );

    \I__4610\ : IoInMux
    port map (
            O => \N__25194\,
            I => \N__25188\
        );

    \I__4609\ : InMux
    port map (
            O => \N__25191\,
            I => \N__25185\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__25188\,
            I => \N__25182\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__25185\,
            I => \N__25179\
        );

    \I__4606\ : Span4Mux_s2_h
    port map (
            O => \N__25182\,
            I => \N__25176\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__25179\,
            I => \N__25173\
        );

    \I__4604\ : Sp12to4
    port map (
            O => \N__25176\,
            I => \N__25170\
        );

    \I__4603\ : Span4Mux_v
    port map (
            O => \N__25173\,
            I => \N__25167\
        );

    \I__4602\ : Span12Mux_s11_v
    port map (
            O => \N__25170\,
            I => \N__25164\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__25167\,
            I => \N__25161\
        );

    \I__4600\ : Odrv12
    port map (
            O => \N__25164\,
            I => v1p8a_ok
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__25161\,
            I => v1p8a_ok
        );

    \I__4598\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25153\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25149\
        );

    \I__4596\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25146\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__25149\,
            I => \N__25143\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__25146\,
            I => \N__25140\
        );

    \I__4593\ : Span4Mux_v
    port map (
            O => \N__25143\,
            I => \N__25135\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__25140\,
            I => \N__25135\
        );

    \I__4591\ : Span4Mux_v
    port map (
            O => \N__25135\,
            I => \N__25132\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__25132\,
            I => slp_susn
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__4588\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25122\
        );

    \I__4587\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25119\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__25122\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__25119\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4584\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25108\
        );

    \I__4583\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25108\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__25108\,
            I => \VPP_VDDQ.count_rst_8\
        );

    \I__4581\ : InMux
    port map (
            O => \N__25105\,
            I => \VPP_VDDQ.un4_count_1_cry_2_cZ0\
        );

    \I__4580\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25098\
        );

    \I__4579\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25095\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__25098\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__25095\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4576\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25084\
        );

    \I__4575\ : InMux
    port map (
            O => \N__25089\,
            I => \N__25084\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__25084\,
            I => \VPP_VDDQ.count_rst_9\
        );

    \I__4573\ : InMux
    port map (
            O => \N__25081\,
            I => \VPP_VDDQ.un4_count_1_cry_3_cZ0\
        );

    \I__4572\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25074\
        );

    \I__4571\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25071\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__25074\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__25071\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__4568\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__4567\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25060\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__25060\,
            I => \VPP_VDDQ.count_rst_10\
        );

    \I__4565\ : InMux
    port map (
            O => \N__25057\,
            I => \VPP_VDDQ.un4_count_1_cry_4_cZ0\
        );

    \I__4564\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25051\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__25051\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4562\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25042\
        );

    \I__4561\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25042\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__25042\,
            I => \VPP_VDDQ.count_rst_11\
        );

    \I__4559\ : InMux
    port map (
            O => \N__25039\,
            I => \VPP_VDDQ.un4_count_1_cry_5\
        );

    \I__4558\ : InMux
    port map (
            O => \N__25036\,
            I => \N__25032\
        );

    \I__4557\ : InMux
    port map (
            O => \N__25035\,
            I => \N__25029\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__25032\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__25029\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4554\ : InMux
    port map (
            O => \N__25024\,
            I => \VPP_VDDQ.un4_count_1_cry_6_cZ0\
        );

    \I__4553\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__25018\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__4551\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__4550\ : InMux
    port map (
            O => \N__25014\,
            I => \N__25009\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__25009\,
            I => \VPP_VDDQ.count_rst_13\
        );

    \I__4548\ : InMux
    port map (
            O => \N__25006\,
            I => \bfn_8_3_0_\
        );

    \I__4547\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24987\
        );

    \I__4546\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24987\
        );

    \I__4545\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24984\
        );

    \I__4544\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24981\
        );

    \I__4543\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24978\
        );

    \I__4542\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24971\
        );

    \I__4541\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24971\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24971\
        );

    \I__4539\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24962\
        );

    \I__4538\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24962\
        );

    \I__4537\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24962\
        );

    \I__4536\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24962\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__24987\,
            I => \N__24959\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__24984\,
            I => \VPP_VDDQ.count_RNI_1_10\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__24981\,
            I => \VPP_VDDQ.count_RNI_1_10\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24978\,
            I => \VPP_VDDQ.count_RNI_1_10\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__24971\,
            I => \VPP_VDDQ.count_RNI_1_10\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__24962\,
            I => \VPP_VDDQ.count_RNI_1_10\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__24959\,
            I => \VPP_VDDQ.count_RNI_1_10\
        );

    \I__4528\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24942\
        );

    \I__4527\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24939\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__24942\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__24939\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__4524\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24928\
        );

    \I__4523\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24928\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__24928\,
            I => \VPP_VDDQ.count_rst_14\
        );

    \I__4521\ : InMux
    port map (
            O => \N__24925\,
            I => \VPP_VDDQ.un4_count_1_cry_8_cZ0\
        );

    \I__4520\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24918\
        );

    \I__4519\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24915\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__24918\,
            I => \N__24912\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__24915\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__24912\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__4515\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24901\
        );

    \I__4514\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24901\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__24901\,
            I => \N__24898\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__24898\,
            I => \VPP_VDDQ.count_rst\
        );

    \I__4511\ : InMux
    port map (
            O => \N__24895\,
            I => \VPP_VDDQ.un4_count_1_cry_9\
        );

    \I__4510\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__24889\,
            I => \VPP_VDDQ.count_3_3\
        );

    \I__4508\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__24883\,
            I => \VPP_VDDQ.count_3_4\
        );

    \I__4506\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24877\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__24877\,
            I => \VPP_VDDQ.count_3_5\
        );

    \I__4504\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24871\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__24871\,
            I => \VPP_VDDQ.un4_count_1_axb_0\
        );

    \I__4502\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24864\
        );

    \I__4501\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24861\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__24864\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__24861\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__4498\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24850\
        );

    \I__4497\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24850\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__24850\,
            I => \VPP_VDDQ.count_rst_6\
        );

    \I__4495\ : InMux
    port map (
            O => \N__24847\,
            I => \VPP_VDDQ.un4_count_1_cry_0\
        );

    \I__4494\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24840\
        );

    \I__4493\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24837\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__24840\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__24837\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__4490\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__4489\ : InMux
    port map (
            O => \N__24831\,
            I => \N__24826\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__24826\,
            I => \VPP_VDDQ.count_rst_7\
        );

    \I__4487\ : InMux
    port map (
            O => \N__24823\,
            I => \VPP_VDDQ.un4_count_1_cry_1\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__24820\,
            I => \N__24816\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__24819\,
            I => \N__24813\
        );

    \I__4484\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24809\
        );

    \I__4483\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24806\
        );

    \I__4482\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24803\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24798\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__24806\,
            I => \N__24798\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__24803\,
            I => \POWERLED.N_332_N\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__24798\,
            I => \POWERLED.N_332_N\
        );

    \I__4477\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24790\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__24790\,
            I => \POWERLED.N_116_f0\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__24787\,
            I => \POWERLED.N_116_f0_cascade_\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__24784\,
            I => \N__24781\
        );

    \I__4473\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24772\
        );

    \I__4472\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24772\
        );

    \I__4471\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24772\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__24772\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__4468\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24763\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__24763\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\
        );

    \I__4466\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24754\
        );

    \I__4465\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24754\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__24754\,
            I => \POWERLED.dutycycle_e_1_9\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__24751\,
            I => \POWERLED.dutycycleZ0Z_6_cascade_\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__24748\,
            I => \POWERLED.N_157_N_cascade_\
        );

    \I__4461\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24742\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__24742\,
            I => \POWERLED.dutycycle_en_4\
        );

    \I__4459\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24733\
        );

    \I__4458\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24733\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__24733\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__24730\,
            I => \POWERLED.dutycycle_en_4_cascade_\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__24727\,
            I => \N__24723\
        );

    \I__4454\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24718\
        );

    \I__4453\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24718\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__24718\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__4451\ : InMux
    port map (
            O => \N__24715\,
            I => \N__24712\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__24712\,
            I => \VPP_VDDQ.un13_clk_100khz_10\
        );

    \I__4449\ : InMux
    port map (
            O => \N__24709\,
            I => \N__24706\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__24706\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__24703\,
            I => \POWERLED.dutycycle_RNI554R1Z0Z_8_cascade_\
        );

    \I__4446\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24697\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__24697\,
            I => \POWERLED.func_state_RNI778D2Z0Z_1\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__24694\,
            I => \POWERLED.func_state_RNI778D2Z0Z_1_cascade_\
        );

    \I__4443\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24688\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__24688\,
            I => \POWERLED.dutycycle_RNIKGV14Z0Z_8\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__24685\,
            I => \POWERLED.dutycycle_RNIKGV14Z0Z_8_cascade_\
        );

    \I__4440\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24679\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__24679\,
            I => \POWERLED.dutycycle_RNI554R1Z0Z_8\
        );

    \I__4438\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24671\
        );

    \I__4437\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24666\
        );

    \I__4436\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24666\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__24671\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__24666\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__4433\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24658\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__24658\,
            I => \POWERLED.g1_2_0\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__24655\,
            I => \POWERLED.func_state_RNI3IN21_0Z0Z_1_cascade_\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__24652\,
            I => \N__24649\
        );

    \I__4429\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24643\
        );

    \I__4428\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24643\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__24643\,
            I => \N__24640\
        );

    \I__4426\ : Span4Mux_h
    port map (
            O => \N__24640\,
            I => \N__24637\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__24637\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__24634\,
            I => \N__24630\
        );

    \I__4423\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24625\
        );

    \I__4422\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24625\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__24625\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__24622\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__4419\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24616\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__24616\,
            I => \N__24613\
        );

    \I__4417\ : Span4Mux_h
    port map (
            O => \N__24613\,
            I => \N__24610\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__24610\,
            I => \POWERLED.dutycycle_RNI3IN21Z0Z_6\
        );

    \I__4415\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24604\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__4413\ : Span4Mux_h
    port map (
            O => \N__24601\,
            I => \N__24596\
        );

    \I__4412\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24591\
        );

    \I__4411\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24591\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__24596\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__24591\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6\
        );

    \I__4408\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__24583\,
            I => \POWERLED.N_312\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__24580\,
            I => \N__24569\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__24579\,
            I => \N__24566\
        );

    \I__4404\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24556\
        );

    \I__4403\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24551\
        );

    \I__4402\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24551\
        );

    \I__4401\ : InMux
    port map (
            O => \N__24575\,
            I => \N__24543\
        );

    \I__4400\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24543\
        );

    \I__4399\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24538\
        );

    \I__4398\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24538\
        );

    \I__4397\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24529\
        );

    \I__4396\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24529\
        );

    \I__4395\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24529\
        );

    \I__4394\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24529\
        );

    \I__4393\ : InMux
    port map (
            O => \N__24563\,
            I => \N__24526\
        );

    \I__4392\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24523\
        );

    \I__4391\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24520\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__24560\,
            I => \N__24517\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__24559\,
            I => \N__24514\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__24556\,
            I => \N__24503\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__24551\,
            I => \N__24503\
        );

    \I__4386\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24496\
        );

    \I__4385\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24496\
        );

    \I__4384\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24496\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__24543\,
            I => \N__24493\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__24538\,
            I => \N__24489\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__24529\,
            I => \N__24486\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__24526\,
            I => \N__24479\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__24523\,
            I => \N__24479\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__24520\,
            I => \N__24479\
        );

    \I__4377\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24474\
        );

    \I__4376\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24474\
        );

    \I__4375\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24471\
        );

    \I__4374\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24468\
        );

    \I__4373\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24465\
        );

    \I__4372\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24458\
        );

    \I__4371\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24458\
        );

    \I__4370\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24458\
        );

    \I__4369\ : Span4Mux_s3_v
    port map (
            O => \N__24503\,
            I => \N__24453\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__24496\,
            I => \N__24453\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__24493\,
            I => \N__24450\
        );

    \I__4366\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24447\
        );

    \I__4365\ : Span4Mux_s3_h
    port map (
            O => \N__24489\,
            I => \N__24440\
        );

    \I__4364\ : Span4Mux_s3_h
    port map (
            O => \N__24486\,
            I => \N__24440\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__24479\,
            I => \N__24440\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__24474\,
            I => \POWERLED.func_state\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__24471\,
            I => \POWERLED.func_state\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__24468\,
            I => \POWERLED.func_state\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__24465\,
            I => \POWERLED.func_state\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__24458\,
            I => \POWERLED.func_state\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__24453\,
            I => \POWERLED.func_state\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__24450\,
            I => \POWERLED.func_state\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__24447\,
            I => \POWERLED.func_state\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__24440\,
            I => \POWERLED.func_state\
        );

    \I__4353\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24417\
        );

    \I__4352\ : InMux
    port map (
            O => \N__24420\,
            I => \N__24414\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__24417\,
            I => \N__24411\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24408\
        );

    \I__4349\ : Span4Mux_s3_h
    port map (
            O => \N__24411\,
            I => \N__24405\
        );

    \I__4348\ : Span4Mux_h
    port map (
            O => \N__24408\,
            I => \N__24402\
        );

    \I__4347\ : Span4Mux_v
    port map (
            O => \N__24405\,
            I => \N__24399\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__24402\,
            I => \POWERLED.N_389\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__24399\,
            I => \POWERLED.N_389\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__4343\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24388\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__24388\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__4341\ : InMux
    port map (
            O => \N__24385\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__24382\,
            I => \N__24378\
        );

    \I__4339\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24370\
        );

    \I__4338\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24370\
        );

    \I__4337\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24370\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__24370\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__4335\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24364\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__24364\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__4333\ : InMux
    port map (
            O => \N__24361\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__4332\ : InMux
    port map (
            O => \N__24358\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__4330\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24349\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__24349\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__24346\,
            I => \N__24343\
        );

    \I__4327\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24340\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__24340\,
            I => \N__24337\
        );

    \I__4325\ : Odrv12
    port map (
            O => \N__24337\,
            I => \POWERLED.g0_13_sx\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__24334\,
            I => \POWERLED.un1_clk_100khz_36_and_i_a2_1_sx_cascade_\
        );

    \I__4323\ : IoInMux
    port map (
            O => \N__24331\,
            I => \N__24328\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__24328\,
            I => \N__24319\
        );

    \I__4321\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24316\
        );

    \I__4320\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24310\
        );

    \I__4319\ : InMux
    port map (
            O => \N__24325\,
            I => \N__24310\
        );

    \I__4318\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24305\
        );

    \I__4317\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24305\
        );

    \I__4316\ : InMux
    port map (
            O => \N__24322\,
            I => \N__24302\
        );

    \I__4315\ : Span4Mux_s2_v
    port map (
            O => \N__24319\,
            I => \N__24297\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__24316\,
            I => \N__24297\
        );

    \I__4313\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24294\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__24310\,
            I => \N__24291\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24286\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24283\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__24297\,
            I => \N__24278\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24278\
        );

    \I__4307\ : Span4Mux_v
    port map (
            O => \N__24291\,
            I => \N__24275\
        );

    \I__4306\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24270\
        );

    \I__4305\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24270\
        );

    \I__4304\ : Span4Mux_s3_v
    port map (
            O => \N__24286\,
            I => \N__24265\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__24283\,
            I => \N__24265\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__24278\,
            I => \N__24262\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__24275\,
            I => rsmrstn
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__24270\,
            I => rsmrstn
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__24265\,
            I => rsmrstn
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__24262\,
            I => rsmrstn
        );

    \I__4297\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24242\
        );

    \I__4296\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24242\
        );

    \I__4295\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24233\
        );

    \I__4294\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24233\
        );

    \I__4293\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24233\
        );

    \I__4292\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24233\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__24247\,
            I => \N__24229\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__24242\,
            I => \N__24224\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__24233\,
            I => \N__24221\
        );

    \I__4288\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24216\
        );

    \I__4287\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24216\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__24228\,
            I => \N__24212\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__24227\,
            I => \N__24207\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__24224\,
            I => \N__24204\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__24221\,
            I => \N__24199\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__24216\,
            I => \N__24199\
        );

    \I__4281\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24190\
        );

    \I__4280\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24190\
        );

    \I__4279\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24190\
        );

    \I__4278\ : InMux
    port map (
            O => \N__24210\,
            I => \N__24190\
        );

    \I__4277\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24187\
        );

    \I__4276\ : Span4Mux_v
    port map (
            O => \N__24204\,
            I => \N__24181\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__24199\,
            I => \N__24181\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24176\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__24187\,
            I => \N__24176\
        );

    \I__4272\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24173\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__24181\,
            I => \curr_state_RNIR5QD1_0_0\
        );

    \I__4270\ : Odrv12
    port map (
            O => \N__24176\,
            I => \curr_state_RNIR5QD1_0_0\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__24173\,
            I => \curr_state_RNIR5QD1_0_0\
        );

    \I__4268\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24160\
        );

    \I__4267\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24160\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__24160\,
            I => \POWERLED.g0_1\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__24157\,
            I => \N__24149\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__24156\,
            I => \N__24146\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__24155\,
            I => \N__24140\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__24154\,
            I => \N__24137\
        );

    \I__4261\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24134\
        );

    \I__4260\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24129\
        );

    \I__4259\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24129\
        );

    \I__4258\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24126\
        );

    \I__4257\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24121\
        );

    \I__4256\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24121\
        );

    \I__4255\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24116\
        );

    \I__4254\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24116\
        );

    \I__4253\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24113\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__24134\,
            I => \N__24106\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__24129\,
            I => \N__24106\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__24126\,
            I => \N__24106\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24101\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__24101\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__24113\,
            I => \SUSWARN_N_fast\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__24106\,
            I => \SUSWARN_N_fast\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__24101\,
            I => \SUSWARN_N_fast\
        );

    \I__4244\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24081\
        );

    \I__4243\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24081\
        );

    \I__4242\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24081\
        );

    \I__4241\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24081\
        );

    \I__4240\ : InMux
    port map (
            O => \N__24090\,
            I => \N__24078\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__24081\,
            I => \N__24075\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24070\
        );

    \I__4237\ : Span4Mux_v
    port map (
            O => \N__24075\,
            I => \N__24070\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__24070\,
            I => \N__24067\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__24067\,
            I => \RSMRST_PWRGD_RSMRSTn_fast\
        );

    \I__4234\ : InMux
    port map (
            O => \N__24064\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__4233\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24058\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__24058\,
            I => \N__24055\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__24055\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__4230\ : InMux
    port map (
            O => \N__24052\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__4229\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24046\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__24046\,
            I => \N__24043\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__24043\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__4226\ : InMux
    port map (
            O => \N__24040\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__4225\ : InMux
    port map (
            O => \N__24037\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__24034\,
            I => \N__24030\
        );

    \I__4223\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24022\
        );

    \I__4222\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24022\
        );

    \I__4221\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24022\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__24022\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__4219\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__24016\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__4217\ : InMux
    port map (
            O => \N__24013\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__24010\,
            I => \N__24007\
        );

    \I__4215\ : InMux
    port map (
            O => \N__24007\,
            I => \N__24004\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__24004\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__4213\ : InMux
    port map (
            O => \N__24001\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__4212\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__23995\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__4210\ : InMux
    port map (
            O => \N__23992\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__23989\,
            I => \POWERLED.N_203_i_cascade_\
        );

    \I__4208\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23983\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23978\
        );

    \I__4206\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23973\
        );

    \I__4205\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23973\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__23978\,
            I => \N__23970\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N__23967\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__23970\,
            I => \N__23964\
        );

    \I__4201\ : Span12Mux_s6_h
    port map (
            O => \N__23967\,
            I => \N__23961\
        );

    \I__4200\ : Odrv4
    port map (
            O => \N__23964\,
            I => \POWERLED.func_state_RNI0TA81_0Z0Z_0\
        );

    \I__4199\ : Odrv12
    port map (
            O => \N__23961\,
            I => \POWERLED.func_state_RNI0TA81_0Z0Z_0\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__23956\,
            I => \N__23953\
        );

    \I__4197\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23949\
        );

    \I__4196\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23946\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__23949\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__23946\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23938\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__23938\,
            I => \N__23935\
        );

    \I__4191\ : Odrv12
    port map (
            O => \N__23935\,
            I => \POWERLED.mult1_un131_sum_axb_4_l_fx\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__23932\,
            I => \N__23929\
        );

    \I__4189\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23917\
        );

    \I__4188\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23917\
        );

    \I__4187\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23917\
        );

    \I__4186\ : InMux
    port map (
            O => \N__23926\,
            I => \N__23912\
        );

    \I__4185\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23912\
        );

    \I__4184\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23909\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__23917\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__23912\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__23909\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__23902\,
            I => \N__23899\
        );

    \I__4179\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23896\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__23896\,
            I => \N__23893\
        );

    \I__4177\ : Odrv12
    port map (
            O => \N__23893\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__4176\ : InMux
    port map (
            O => \N__23890\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__4175\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__23881\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__4172\ : InMux
    port map (
            O => \N__23878\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__23875\,
            I => \N__23872\
        );

    \I__4170\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23869\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__23869\,
            I => \N__23866\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__23866\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__4167\ : InMux
    port map (
            O => \N__23863\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__23860\,
            I => \N__23857\
        );

    \I__4165\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23854\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__23854\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__4163\ : InMux
    port map (
            O => \N__23851\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__4162\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23845\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__23845\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__4160\ : InMux
    port map (
            O => \N__23842\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__23839\,
            I => \N__23836\
        );

    \I__4158\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23832\
        );

    \I__4157\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23829\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__23832\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__23829\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__4154\ : InMux
    port map (
            O => \N__23824\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__4153\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23818\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__23818\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__4151\ : InMux
    port map (
            O => \N__23815\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__4150\ : InMux
    port map (
            O => \N__23812\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__23809\,
            I => \POWERLED.mult1_un124_sum_s_8_cascade_\
        );

    \I__4148\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__23803\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__4146\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23797\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__23797\,
            I => \VPP_VDDQ.count_3_15\
        );

    \I__4144\ : InMux
    port map (
            O => \N__23794\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__4143\ : InMux
    port map (
            O => \N__23791\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__4142\ : InMux
    port map (
            O => \N__23788\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__4141\ : InMux
    port map (
            O => \N__23785\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__4140\ : InMux
    port map (
            O => \N__23782\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__4139\ : InMux
    port map (
            O => \N__23779\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__4138\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23773\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__23773\,
            I => \POWERLED.mult1_un131_sum_axb_7_l_fx\
        );

    \I__4136\ : InMux
    port map (
            O => \N__23770\,
            I => \bfn_7_6_0_\
        );

    \I__4135\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23764\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__23764\,
            I => \VPP_VDDQ.curr_state_2_0_1\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__23761\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__4132\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23752\
        );

    \I__4131\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23752\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__23752\,
            I => \VPP_VDDQ.m4_0_a2\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__23749\,
            I => \VPP_VDDQ.m4_0_cascade_\
        );

    \I__4128\ : IoInMux
    port map (
            O => \N__23746\,
            I => \N__23729\
        );

    \I__4127\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23717\
        );

    \I__4126\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23717\
        );

    \I__4125\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23717\
        );

    \I__4124\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23714\
        );

    \I__4123\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23705\
        );

    \I__4122\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23705\
        );

    \I__4121\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23705\
        );

    \I__4120\ : InMux
    port map (
            O => \N__23738\,
            I => \N__23705\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__23737\,
            I => \N__23701\
        );

    \I__4118\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23694\
        );

    \I__4117\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23694\
        );

    \I__4116\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23694\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \N__23691\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__23732\,
            I => \N__23688\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__23729\,
            I => \N__23682\
        );

    \I__4112\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23675\
        );

    \I__4111\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23675\
        );

    \I__4110\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23675\
        );

    \I__4109\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23670\
        );

    \I__4108\ : InMux
    port map (
            O => \N__23724\,
            I => \N__23670\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23651\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__23714\,
            I => \N__23651\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23651\
        );

    \I__4104\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23648\
        );

    \I__4103\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23641\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__23694\,
            I => \N__23634\
        );

    \I__4101\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23627\
        );

    \I__4100\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23627\
        );

    \I__4099\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23627\
        );

    \I__4098\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23619\
        );

    \I__4097\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23619\
        );

    \I__4096\ : IoSpan4Mux
    port map (
            O => \N__23682\,
            I => \N__23616\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__23675\,
            I => \N__23611\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__23670\,
            I => \N__23611\
        );

    \I__4093\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23606\
        );

    \I__4092\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23606\
        );

    \I__4091\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23601\
        );

    \I__4090\ : InMux
    port map (
            O => \N__23666\,
            I => \N__23601\
        );

    \I__4089\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23598\
        );

    \I__4088\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23591\
        );

    \I__4087\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23591\
        );

    \I__4086\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23591\
        );

    \I__4085\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23584\
        );

    \I__4084\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23584\
        );

    \I__4083\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23584\
        );

    \I__4082\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23581\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__23651\,
            I => \N__23576\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__23648\,
            I => \N__23576\
        );

    \I__4079\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23560\
        );

    \I__4078\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23560\
        );

    \I__4077\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23560\
        );

    \I__4076\ : InMux
    port map (
            O => \N__23644\,
            I => \N__23560\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__23641\,
            I => \N__23557\
        );

    \I__4074\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23543\
        );

    \I__4073\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23543\
        );

    \I__4072\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23543\
        );

    \I__4071\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23543\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__23634\,
            I => \N__23538\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__23627\,
            I => \N__23538\
        );

    \I__4068\ : InMux
    port map (
            O => \N__23626\,
            I => \N__23531\
        );

    \I__4067\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23531\
        );

    \I__4066\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23531\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__23619\,
            I => \N__23528\
        );

    \I__4064\ : Span4Mux_s3_h
    port map (
            O => \N__23616\,
            I => \N__23523\
        );

    \I__4063\ : Span4Mux_s1_v
    port map (
            O => \N__23611\,
            I => \N__23523\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__23606\,
            I => \N__23518\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__23601\,
            I => \N__23518\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__23598\,
            I => \N__23513\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__23591\,
            I => \N__23513\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__23584\,
            I => \N__23506\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__23581\,
            I => \N__23506\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__23576\,
            I => \N__23506\
        );

    \I__4055\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23503\
        );

    \I__4054\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23490\
        );

    \I__4053\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23490\
        );

    \I__4052\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23490\
        );

    \I__4051\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23490\
        );

    \I__4050\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23490\
        );

    \I__4049\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23490\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__23560\,
            I => \N__23485\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__23557\,
            I => \N__23485\
        );

    \I__4046\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23480\
        );

    \I__4045\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23480\
        );

    \I__4044\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23473\
        );

    \I__4043\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23473\
        );

    \I__4042\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23473\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__23543\,
            I => \N__23468\
        );

    \I__4040\ : Span4Mux_h
    port map (
            O => \N__23538\,
            I => \N__23468\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23459\
        );

    \I__4038\ : Span4Mux_v
    port map (
            O => \N__23528\,
            I => \N__23459\
        );

    \I__4037\ : Span4Mux_v
    port map (
            O => \N__23523\,
            I => \N__23459\
        );

    \I__4036\ : Span4Mux_v
    port map (
            O => \N__23518\,
            I => \N__23459\
        );

    \I__4035\ : Span4Mux_s3_v
    port map (
            O => \N__23513\,
            I => \N__23454\
        );

    \I__4034\ : Span4Mux_v
    port map (
            O => \N__23506\,
            I => \N__23454\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__23503\,
            I => suswarn_n
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__23490\,
            I => suswarn_n
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__23485\,
            I => suswarn_n
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__23480\,
            I => suswarn_n
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__23473\,
            I => suswarn_n
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__23468\,
            I => suswarn_n
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__23459\,
            I => suswarn_n
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__23454\,
            I => suswarn_n
        );

    \I__4025\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23434\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N__23430\
        );

    \I__4023\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23427\
        );

    \I__4022\ : Span4Mux_h
    port map (
            O => \N__23430\,
            I => \N__23424\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__23427\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__23424\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__23419\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__4018\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23411\
        );

    \I__4017\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23406\
        );

    \I__4016\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23406\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__23411\,
            I => \VPP_VDDQ.N_2877_i\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__23406\,
            I => \VPP_VDDQ.N_2877_i\
        );

    \I__4013\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23394\
        );

    \I__4012\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23394\
        );

    \I__4011\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23391\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__23394\,
            I => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__23391\,
            I => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__23386\,
            I => \VPP_VDDQ.N_2877_i_cascade_\
        );

    \I__4007\ : InMux
    port map (
            O => \N__23383\,
            I => \N__23380\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23375\
        );

    \I__4005\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23370\
        );

    \I__4004\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23370\
        );

    \I__4003\ : Span4Mux_h
    port map (
            O => \N__23375\,
            I => \N__23367\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__23370\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__23367\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__4000\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23359\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__23359\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__3998\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23352\
        );

    \I__3997\ : InMux
    port map (
            O => \N__23355\,
            I => \N__23349\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__23352\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__23349\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__3994\ : InMux
    port map (
            O => \N__23344\,
            I => \DSW_PWRGD.un1_count_1_cry_5\
        );

    \I__3993\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23337\
        );

    \I__3992\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23334\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__23337\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__23334\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__3989\ : InMux
    port map (
            O => \N__23329\,
            I => \DSW_PWRGD.un1_count_1_cry_6\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__23326\,
            I => \N__23322\
        );

    \I__3987\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23319\
        );

    \I__3986\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23316\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__23319\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__23316\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__3983\ : InMux
    port map (
            O => \N__23311\,
            I => \bfn_7_5_0_\
        );

    \I__3982\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23304\
        );

    \I__3981\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23301\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__23304\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__23301\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__3978\ : InMux
    port map (
            O => \N__23296\,
            I => \DSW_PWRGD.un1_count_1_cry_8\
        );

    \I__3977\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23289\
        );

    \I__3976\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23286\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__23289\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__23286\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__3973\ : InMux
    port map (
            O => \N__23281\,
            I => \DSW_PWRGD.un1_count_1_cry_9\
        );

    \I__3972\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23274\
        );

    \I__3971\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23271\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__23274\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__23271\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__3968\ : InMux
    port map (
            O => \N__23266\,
            I => \DSW_PWRGD.un1_count_1_cry_10\
        );

    \I__3967\ : InMux
    port map (
            O => \N__23263\,
            I => \DSW_PWRGD.un1_count_1_cry_11\
        );

    \I__3966\ : InMux
    port map (
            O => \N__23260\,
            I => \DSW_PWRGD.un1_count_1_cry_12\
        );

    \I__3965\ : InMux
    port map (
            O => \N__23257\,
            I => \DSW_PWRGD.un1_count_1_cry_13\
        );

    \I__3964\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23251\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__23251\,
            I => \VPP_VDDQ.count_3_8\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__23248\,
            I => \VPP_VDDQ.countZ0Z_8_cascade_\
        );

    \I__3961\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23242\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__23242\,
            I => \VPP_VDDQ.un13_clk_100khz_11\
        );

    \I__3959\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23235\
        );

    \I__3958\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23232\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__23235\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__23232\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__23227\,
            I => \N__23223\
        );

    \I__3954\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23220\
        );

    \I__3953\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23217\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__23220\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__23217\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__3950\ : InMux
    port map (
            O => \N__23212\,
            I => \DSW_PWRGD.un1_count_1_cry_0\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__23209\,
            I => \N__23205\
        );

    \I__3948\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23202\
        );

    \I__3947\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23199\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__23202\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__23199\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__3944\ : InMux
    port map (
            O => \N__23194\,
            I => \DSW_PWRGD.un1_count_1_cry_1\
        );

    \I__3943\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23187\
        );

    \I__3942\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23184\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__23187\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__23184\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__3939\ : InMux
    port map (
            O => \N__23179\,
            I => \DSW_PWRGD.un1_count_1_cry_2\
        );

    \I__3938\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23172\
        );

    \I__3937\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23169\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__23172\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__23169\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__3934\ : InMux
    port map (
            O => \N__23164\,
            I => \DSW_PWRGD.un1_count_1_cry_3\
        );

    \I__3933\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23157\
        );

    \I__3932\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23154\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__23157\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__23154\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__3929\ : InMux
    port map (
            O => \N__23149\,
            I => \DSW_PWRGD.un1_count_1_cry_4\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__23146\,
            I => \VPP_VDDQ.un13_clk_100khz_9_cascade_\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__23143\,
            I => \VPP_VDDQ.count_RNI_1_10_cascade_\
        );

    \I__3926\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__23137\,
            I => \VPP_VDDQ.count_3_11\
        );

    \I__3924\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23125\
        );

    \I__3923\ : InMux
    port map (
            O => \N__23133\,
            I => \N__23125\
        );

    \I__3922\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23125\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__23125\,
            I => \VPP_VDDQ.N_3013_i\
        );

    \I__3920\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23116\
        );

    \I__3919\ : InMux
    port map (
            O => \N__23121\,
            I => \N__23116\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__23116\,
            I => \VPP_VDDQ.count_3_0\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \VPP_VDDQ.count_en_cascade_\
        );

    \I__3916\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23107\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__23107\,
            I => \VPP_VDDQ.count_3_1\
        );

    \I__3914\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__23101\,
            I => \VPP_VDDQ.count_3_9\
        );

    \I__3912\ : InMux
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__23095\,
            I => \VPP_VDDQ.count_3_6\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__23092\,
            I => \VPP_VDDQ.countZ0Z_6_cascade_\
        );

    \I__3909\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__23086\,
            I => \VPP_VDDQ.count_3_10\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__23083\,
            I => \VPP_VDDQ.count_rst_5_cascade_\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__23080\,
            I => \VPP_VDDQ.N_3013_i_cascade_\
        );

    \I__3905\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__23071\,
            I => \VPP_VDDQ.un13_clk_100khz_8\
        );

    \I__3902\ : InMux
    port map (
            O => \N__23068\,
            I => \POWERLED.un1_dutycycle_94_cry_9\
        );

    \I__3901\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23059\
        );

    \I__3900\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23059\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__23059\,
            I => \POWERLED.dutycycle_rst_6\
        );

    \I__3898\ : InMux
    port map (
            O => \N__23056\,
            I => \POWERLED.un1_dutycycle_94_cry_10_cZ0\
        );

    \I__3897\ : InMux
    port map (
            O => \N__23053\,
            I => \POWERLED.un1_dutycycle_94_cry_11\
        );

    \I__3896\ : InMux
    port map (
            O => \N__23050\,
            I => \POWERLED.un1_dutycycle_94_cry_12\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__23047\,
            I => \N__23038\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__23046\,
            I => \N__23035\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__23045\,
            I => \N__23032\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__23044\,
            I => \N__23028\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__23043\,
            I => \N__23021\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__23042\,
            I => \N__23018\
        );

    \I__3889\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23003\
        );

    \I__3888\ : InMux
    port map (
            O => \N__23038\,
            I => \N__23003\
        );

    \I__3887\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23003\
        );

    \I__3886\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23003\
        );

    \I__3885\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23003\
        );

    \I__3884\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23003\
        );

    \I__3883\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23003\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__23026\,
            I => \N__23000\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__23025\,
            I => \N__22996\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__23024\,
            I => \N__22992\
        );

    \I__3879\ : InMux
    port map (
            O => \N__23021\,
            I => \N__22987\
        );

    \I__3878\ : InMux
    port map (
            O => \N__23018\,
            I => \N__22987\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__23003\,
            I => \N__22984\
        );

    \I__3876\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22973\
        );

    \I__3875\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22973\
        );

    \I__3874\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22973\
        );

    \I__3873\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22973\
        );

    \I__3872\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22973\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__22987\,
            I => \N__22966\
        );

    \I__3870\ : Span4Mux_s1_v
    port map (
            O => \N__22984\,
            I => \N__22966\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22966\
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__22966\,
            I => \POWERLED.N_175_i\
        );

    \I__3867\ : InMux
    port map (
            O => \N__22963\,
            I => \POWERLED.un1_dutycycle_94_cry_13\
        );

    \I__3866\ : InMux
    port map (
            O => \N__22960\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__3865\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22954\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__22954\,
            I => \VPP_VDDQ.count_3_2\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__3862\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__22945\,
            I => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\
        );

    \I__3860\ : InMux
    port map (
            O => \N__22942\,
            I => \POWERLED.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__3859\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__22936\,
            I => \N__22933\
        );

    \I__3857\ : Span4Mux_v
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__22930\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22927\,
            I => \POWERLED.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__3854\ : InMux
    port map (
            O => \N__22924\,
            I => \POWERLED.un1_dutycycle_94_cry_2_cZ0\
        );

    \I__3853\ : InMux
    port map (
            O => \N__22921\,
            I => \POWERLED.un1_dutycycle_94_cry_3\
        );

    \I__3852\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__22915\,
            I => \POWERLED.N_308\
        );

    \I__3850\ : InMux
    port map (
            O => \N__22912\,
            I => \POWERLED.un1_dutycycle_94_cry_4_cZ0\
        );

    \I__3849\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22906\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__22906\,
            I => \POWERLED.N_307\
        );

    \I__3847\ : InMux
    port map (
            O => \N__22903\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3846\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22894\
        );

    \I__3845\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22894\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__22891\,
            I => \N__22888\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__22888\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__3841\ : InMux
    port map (
            O => \N__22885\,
            I => \POWERLED.un1_dutycycle_94_cry_6\
        );

    \I__3840\ : InMux
    port map (
            O => \N__22882\,
            I => \bfn_6_16_0_\
        );

    \I__3839\ : InMux
    port map (
            O => \N__22879\,
            I => \POWERLED.un1_dutycycle_94_cry_8\
        );

    \I__3838\ : InMux
    port map (
            O => \N__22876\,
            I => \N__22873\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__22873\,
            I => \POWERLED.func_state_RNIDUQ02Z0Z_1\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__22870\,
            I => \POWERLED.un1_clk_100khz_51_and_i_m2_0_1_cascade_\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__22867\,
            I => \POWERLED.N_233_N_cascade_\
        );

    \I__3834\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22861\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__22861\,
            I => \POWERLED.N_311\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__22858\,
            I => \POWERLED.dutycycle_eena_13_cascade_\
        );

    \I__3831\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22849\
        );

    \I__3830\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22849\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__22849\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7TZ0Z3\
        );

    \I__3828\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__22843\,
            I => \POWERLED.dutycycle_eena_13\
        );

    \I__3826\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22834\
        );

    \I__3825\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22834\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__22834\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__22831\,
            I => \N__22825\
        );

    \I__3822\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22820\
        );

    \I__3821\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22820\
        );

    \I__3820\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22817\
        );

    \I__3819\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22814\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22811\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__22817\,
            I => \N__22807\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__22814\,
            I => \N__22804\
        );

    \I__3815\ : Span4Mux_s3_v
    port map (
            O => \N__22811\,
            I => \N__22801\
        );

    \I__3814\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22798\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__22807\,
            I => \N__22795\
        );

    \I__3812\ : Odrv12
    port map (
            O => \N__22804\,
            I => \POWERLED.N_388\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__22801\,
            I => \POWERLED.N_388\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__22798\,
            I => \POWERLED.N_388\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__22795\,
            I => \POWERLED.N_388\
        );

    \I__3808\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22783\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__3806\ : Odrv12
    port map (
            O => \N__22780\,
            I => \POWERLED_dutycycle_set_1\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__22777\,
            I => \N__22774\
        );

    \I__3804\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22769\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__22773\,
            I => \N__22766\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__22772\,
            I => \N__22763\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22760\
        );

    \I__3800\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22755\
        );

    \I__3799\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22755\
        );

    \I__3798\ : Span4Mux_s3_v
    port map (
            O => \N__22760\,
            I => \N__22752\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__22755\,
            I => \N__22749\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__22752\,
            I => \POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__22749\,
            I => \POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__3794\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22741\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__22741\,
            I => \N__22731\
        );

    \I__3792\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22726\
        );

    \I__3791\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22726\
        );

    \I__3790\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22723\
        );

    \I__3789\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22713\
        );

    \I__3788\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22713\
        );

    \I__3787\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22713\
        );

    \I__3786\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22713\
        );

    \I__3785\ : Span4Mux_v
    port map (
            O => \N__22731\,
            I => \N__22708\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__22726\,
            I => \N__22708\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__22723\,
            I => \N__22705\
        );

    \I__3782\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22702\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22699\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__22708\,
            I => \N__22696\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__22705\,
            I => \N__22693\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__22702\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3777\ : Odrv12
    port map (
            O => \N__22699\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__22696\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__22693\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__22684\,
            I => \N__22681\
        );

    \I__3773\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22678\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22675\
        );

    \I__3771\ : Odrv12
    port map (
            O => \N__22675\,
            I => \POWERLED.un1_func_state25_6_0_o_N_337_N\
        );

    \I__3770\ : CascadeMux
    port map (
            O => \N__22672\,
            I => \POWERLED.N_31_cascade_\
        );

    \I__3769\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22666\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__22666\,
            I => \POWERLED.g0_i_a6_0\
        );

    \I__3767\ : InMux
    port map (
            O => \N__22663\,
            I => \N__22660\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__22660\,
            I => \POWERLED.N_237\
        );

    \I__3765\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__22651\,
            I => \N__22648\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__22648\,
            I => \POWERLED.un1_clk_100khz_52_and_i_0_1_1\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__22645\,
            I => \POWERLED.N_387_cascade_\
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__22642\,
            I => \N__22635\
        );

    \I__3759\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22626\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__22640\,
            I => \N__22622\
        );

    \I__3757\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22613\
        );

    \I__3756\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22613\
        );

    \I__3755\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22613\
        );

    \I__3754\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22613\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__22633\,
            I => \N__22609\
        );

    \I__3752\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22600\
        );

    \I__3751\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22600\
        );

    \I__3750\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22595\
        );

    \I__3749\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22595\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__22626\,
            I => \N__22592\
        );

    \I__3747\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22589\
        );

    \I__3746\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22586\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22583\
        );

    \I__3744\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22576\
        );

    \I__3743\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22576\
        );

    \I__3742\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22576\
        );

    \I__3741\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22572\
        );

    \I__3740\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22569\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__22605\,
            I => \N__22566\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__22600\,
            I => \N__22558\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__22595\,
            I => \N__22558\
        );

    \I__3736\ : Span4Mux_h
    port map (
            O => \N__22592\,
            I => \N__22555\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__22589\,
            I => \N__22550\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22550\
        );

    \I__3733\ : Span4Mux_v
    port map (
            O => \N__22583\,
            I => \N__22547\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__22576\,
            I => \N__22544\
        );

    \I__3731\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22541\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__22572\,
            I => \N__22536\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__22569\,
            I => \N__22536\
        );

    \I__3728\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22527\
        );

    \I__3727\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22527\
        );

    \I__3726\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22527\
        );

    \I__3725\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22527\
        );

    \I__3724\ : Span4Mux_h
    port map (
            O => \N__22558\,
            I => \N__22524\
        );

    \I__3723\ : Span4Mux_v
    port map (
            O => \N__22555\,
            I => \N__22519\
        );

    \I__3722\ : Span4Mux_v
    port map (
            O => \N__22550\,
            I => \N__22519\
        );

    \I__3721\ : Span4Mux_h
    port map (
            O => \N__22547\,
            I => \N__22512\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__22544\,
            I => \N__22512\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22512\
        );

    \I__3718\ : Span4Mux_h
    port map (
            O => \N__22536\,
            I => \N__22509\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__22527\,
            I => \N__22506\
        );

    \I__3716\ : Span4Mux_v
    port map (
            O => \N__22524\,
            I => \N__22503\
        );

    \I__3715\ : IoSpan4Mux
    port map (
            O => \N__22519\,
            I => \N__22498\
        );

    \I__3714\ : IoSpan4Mux
    port map (
            O => \N__22512\,
            I => \N__22498\
        );

    \I__3713\ : Span4Mux_v
    port map (
            O => \N__22509\,
            I => \N__22493\
        );

    \I__3712\ : Span4Mux_v
    port map (
            O => \N__22506\,
            I => \N__22493\
        );

    \I__3711\ : Span4Mux_h
    port map (
            O => \N__22503\,
            I => \N__22490\
        );

    \I__3710\ : IoSpan4Mux
    port map (
            O => \N__22498\,
            I => \N__22487\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__22493\,
            I => \N__22484\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__22490\,
            I => slp_s3n
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__22487\,
            I => slp_s3n
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__22484\,
            I => slp_s3n
        );

    \I__3705\ : InMux
    port map (
            O => \N__22477\,
            I => \N__22467\
        );

    \I__3704\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22462\
        );

    \I__3703\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22462\
        );

    \I__3702\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22454\
        );

    \I__3701\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22447\
        );

    \I__3700\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22447\
        );

    \I__3699\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22447\
        );

    \I__3698\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22444\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__22467\,
            I => \N__22440\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__22462\,
            I => \N__22437\
        );

    \I__3695\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22426\
        );

    \I__3694\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22426\
        );

    \I__3693\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22426\
        );

    \I__3692\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22426\
        );

    \I__3691\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22426\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22414\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__22447\,
            I => \N__22414\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__22444\,
            I => \N__22414\
        );

    \I__3687\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22411\
        );

    \I__3686\ : Span4Mux_h
    port map (
            O => \N__22440\,
            I => \N__22404\
        );

    \I__3685\ : Span4Mux_s3_h
    port map (
            O => \N__22437\,
            I => \N__22401\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22398\
        );

    \I__3683\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22389\
        );

    \I__3682\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22389\
        );

    \I__3681\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22389\
        );

    \I__3680\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22389\
        );

    \I__3679\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22386\
        );

    \I__3678\ : Span4Mux_h
    port map (
            O => \N__22414\,
            I => \N__22383\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22380\
        );

    \I__3676\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22377\
        );

    \I__3675\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22370\
        );

    \I__3674\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22370\
        );

    \I__3673\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22370\
        );

    \I__3672\ : Span4Mux_v
    port map (
            O => \N__22404\,
            I => \N__22367\
        );

    \I__3671\ : Span4Mux_v
    port map (
            O => \N__22401\,
            I => \N__22362\
        );

    \I__3670\ : Span4Mux_h
    port map (
            O => \N__22398\,
            I => \N__22362\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__22389\,
            I => \N__22357\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22357\
        );

    \I__3667\ : Span4Mux_v
    port map (
            O => \N__22383\,
            I => \N__22352\
        );

    \I__3666\ : Span4Mux_h
    port map (
            O => \N__22380\,
            I => \N__22352\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__22377\,
            I => \N__22347\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22347\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__22367\,
            I => slp_s4n
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__22362\,
            I => slp_s4n
        );

    \I__3661\ : Odrv12
    port map (
            O => \N__22357\,
            I => slp_s4n
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__22352\,
            I => slp_s4n
        );

    \I__3659\ : Odrv12
    port map (
            O => \N__22347\,
            I => slp_s4n
        );

    \I__3658\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22333\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__22333\,
            I => \N__22328\
        );

    \I__3656\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22325\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \N__22320\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__22328\,
            I => \N__22310\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22310\
        );

    \I__3652\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22307\
        );

    \I__3651\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22298\
        );

    \I__3650\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22298\
        );

    \I__3649\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22298\
        );

    \I__3648\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22298\
        );

    \I__3647\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22293\
        );

    \I__3646\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22293\
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__22315\,
            I => \N__22285\
        );

    \I__3644\ : Span4Mux_h
    port map (
            O => \N__22310\,
            I => \N__22275\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22275\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22275\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22275\
        );

    \I__3640\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22270\
        );

    \I__3639\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22270\
        );

    \I__3638\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22263\
        );

    \I__3637\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22263\
        );

    \I__3636\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22263\
        );

    \I__3635\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22258\
        );

    \I__3634\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22258\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__22275\,
            I => \N__22253\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22253\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__22263\,
            I => \N__22250\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__22258\,
            I => \N__22247\
        );

    \I__3629\ : Span4Mux_v
    port map (
            O => \N__22253\,
            I => \N__22244\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__22250\,
            I => \N__22241\
        );

    \I__3627\ : Sp12to4
    port map (
            O => \N__22247\,
            I => \N__22238\
        );

    \I__3626\ : Span4Mux_h
    port map (
            O => \N__22244\,
            I => \N__22233\
        );

    \I__3625\ : Span4Mux_h
    port map (
            O => \N__22241\,
            I => \N__22233\
        );

    \I__3624\ : Span12Mux_v
    port map (
            O => \N__22238\,
            I => \N__22230\
        );

    \I__3623\ : IoSpan4Mux
    port map (
            O => \N__22233\,
            I => \N__22227\
        );

    \I__3622\ : Odrv12
    port map (
            O => \N__22230\,
            I => gpio_fpga_soc_4
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__22227\,
            I => gpio_fpga_soc_4
        );

    \I__3620\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22216\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__22221\,
            I => \N__22213\
        );

    \I__3618\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22207\
        );

    \I__3617\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22207\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22204\
        );

    \I__3615\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22199\
        );

    \I__3614\ : InMux
    port map (
            O => \N__22212\,
            I => \N__22196\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22191\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__22204\,
            I => \N__22191\
        );

    \I__3611\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22186\
        );

    \I__3610\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22186\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__22199\,
            I => \POWERLED.N_372\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__22196\,
            I => \POWERLED.N_372\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__22191\,
            I => \POWERLED.N_372\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__22186\,
            I => \POWERLED.N_372\
        );

    \I__3605\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22171\
        );

    \I__3604\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22171\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__3602\ : Span4Mux_h
    port map (
            O => \N__22168\,
            I => \N__22165\
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__22165\,
            I => \POWERLED_un1_clk_100khz_52_and_i_0\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__22162\,
            I => \COUNTER.N_96_mux_i_i_a8_1_cascade_\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__22159\,
            I => \tmp_1_rep1_RNIC08FV_0_cascade_\
        );

    \I__3598\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22153\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__22153\,
            I => \N__22150\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__22150\,
            I => \POWERLED.dutycycle_RNII69M3Z0Z_5\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__22147\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_6_cascade_\
        );

    \I__3594\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__22141\,
            I => \N_96_mux_i_i_3\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__22138\,
            I => \N_96_mux_i_i_3_cascade_\
        );

    \I__3591\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__22132\,
            I => \COUNTER.N_96_mux_i_i_a8_1\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__22129\,
            I => \N__22125\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__22128\,
            I => \N__22122\
        );

    \I__3587\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22117\
        );

    \I__3586\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22117\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__22117\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3584\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__22111\,
            I => \POWERLED.N_31\
        );

    \I__3582\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22105\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__22105\,
            I => \N__22102\
        );

    \I__3580\ : Span4Mux_h
    port map (
            O => \N__22102\,
            I => \N__22097\
        );

    \I__3579\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22091\
        );

    \I__3578\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22091\
        );

    \I__3577\ : Sp12to4
    port map (
            O => \N__22097\,
            I => \N__22085\
        );

    \I__3576\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22082\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__22091\,
            I => \N__22079\
        );

    \I__3574\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22072\
        );

    \I__3573\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22072\
        );

    \I__3572\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22072\
        );

    \I__3571\ : Odrv12
    port map (
            O => \N__22085\,
            I => \SUSWARN_N_rep1\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__22082\,
            I => \SUSWARN_N_rep1\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__22079\,
            I => \SUSWARN_N_rep1\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__22072\,
            I => \SUSWARN_N_rep1\
        );

    \I__3567\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22058\
        );

    \I__3566\ : InMux
    port map (
            O => \N__22062\,
            I => \N__22053\
        );

    \I__3565\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22053\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22050\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__22053\,
            I => \N_414\
        );

    \I__3562\ : Odrv12
    port map (
            O => \N__22050\,
            I => \N_414\
        );

    \I__3561\ : IoInMux
    port map (
            O => \N__22045\,
            I => \N__22042\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__22042\,
            I => \N__22039\
        );

    \I__3559\ : Span4Mux_s3_v
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__22036\,
            I => \HDA_STRAP.count_enZ0\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__22033\,
            I => \N__22024\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__22032\,
            I => \N__22019\
        );

    \I__3555\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22007\
        );

    \I__3554\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22007\
        );

    \I__3553\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22007\
        );

    \I__3552\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22007\
        );

    \I__3551\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22000\
        );

    \I__3550\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22000\
        );

    \I__3549\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22000\
        );

    \I__3548\ : InMux
    port map (
            O => \N__22022\,
            I => \N__21991\
        );

    \I__3547\ : InMux
    port map (
            O => \N__22019\,
            I => \N__21991\
        );

    \I__3546\ : InMux
    port map (
            O => \N__22018\,
            I => \N__21991\
        );

    \I__3545\ : InMux
    port map (
            O => \N__22017\,
            I => \N__21991\
        );

    \I__3544\ : InMux
    port map (
            O => \N__22016\,
            I => \N__21988\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__22007\,
            I => \N__21985\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__22000\,
            I => \N__21980\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21980\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__21988\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__3539\ : Odrv12
    port map (
            O => \N__21985\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__3538\ : Odrv12
    port map (
            O => \N__21980\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__3537\ : IoInMux
    port map (
            O => \N__21973\,
            I => \N__21970\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21967\
        );

    \I__3535\ : Span4Mux_s3_h
    port map (
            O => \N__21967\,
            I => \N__21964\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__21961\,
            I => v1p8a_en
        );

    \I__3532\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21953\
        );

    \I__3531\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21950\
        );

    \I__3530\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21947\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__21953\,
            I => \N__21939\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__21950\,
            I => \N__21934\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21934\
        );

    \I__3526\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21923\
        );

    \I__3525\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21923\
        );

    \I__3524\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21923\
        );

    \I__3523\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21923\
        );

    \I__3522\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21923\
        );

    \I__3521\ : Span12Mux_s8_h
    port map (
            O => \N__21939\,
            I => \N__21920\
        );

    \I__3520\ : Span4Mux_v
    port map (
            O => \N__21934\,
            I => \N__21917\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__21923\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__3518\ : Odrv12
    port map (
            O => \N__21920\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__21917\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__3516\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21904\
        );

    \I__3515\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21899\
        );

    \I__3514\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21899\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__21907\,
            I => \N__21894\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21889\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21886\
        );

    \I__3510\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21881\
        );

    \I__3509\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21881\
        );

    \I__3508\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21874\
        );

    \I__3507\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21874\
        );

    \I__3506\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21874\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__21889\,
            I => \N__21871\
        );

    \I__3504\ : Span4Mux_s3_h
    port map (
            O => \N__21886\,
            I => \N__21868\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__21881\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__21874\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__21871\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__21868\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21844\
        );

    \I__3498\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21844\
        );

    \I__3497\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21844\
        );

    \I__3496\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21844\
        );

    \I__3495\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21844\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__21844\,
            I => \N__21840\
        );

    \I__3493\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21837\
        );

    \I__3492\ : Span4Mux_v
    port map (
            O => \N__21840\,
            I => \N__21834\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__21837\,
            I => \RSMRSTn_0\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__21834\,
            I => \RSMRSTn_0\
        );

    \I__3489\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21826\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__21826\,
            I => \N__21823\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__21823\,
            I => \N__21818\
        );

    \I__3486\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21813\
        );

    \I__3485\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21813\
        );

    \I__3484\ : Span4Mux_v
    port map (
            O => \N__21818\,
            I => \N__21810\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__21813\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__21810\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3481\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21801\
        );

    \I__3480\ : InMux
    port map (
            O => \N__21804\,
            I => \N__21798\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__21801\,
            I => \N__21795\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__21798\,
            I => \N__21792\
        );

    \I__3477\ : Span12Mux_s5_h
    port map (
            O => \N__21795\,
            I => \N__21787\
        );

    \I__3476\ : Span12Mux_s0_v
    port map (
            O => \N__21792\,
            I => \N__21787\
        );

    \I__3475\ : Odrv12
    port map (
            O => \N__21787\,
            I => \HDA_STRAP.N_2989_i\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__3473\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21775\
        );

    \I__3472\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21775\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__21775\,
            I => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\
        );

    \I__3470\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__21769\,
            I => \POWERLED.count_0_15\
        );

    \I__3468\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21760\
        );

    \I__3467\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21760\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__21760\,
            I => \POWERLED.count_1_7\
        );

    \I__3465\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21754\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__21754\,
            I => \POWERLED.count_0_7\
        );

    \I__3463\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21745\
        );

    \I__3462\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21745\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__21745\,
            I => \POWERLED.count_1_8\
        );

    \I__3460\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21739\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__21739\,
            I => \POWERLED.count_0_8\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__21736\,
            I => \N__21732\
        );

    \I__3457\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21727\
        );

    \I__3456\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21727\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__21727\,
            I => \POWERLED.count_1_9\
        );

    \I__3454\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__21721\,
            I => \POWERLED.count_0_9\
        );

    \I__3452\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__21715\,
            I => \POWERLED.g0_8_sx\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__21712\,
            I => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0_cascade_\
        );

    \I__3449\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21703\
        );

    \I__3448\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21703\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__21703\,
            I => \VPP_VDDQ.delayed_vddq_ok_0\
        );

    \I__3446\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21697\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__21697\,
            I => \N__21694\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__21694\,
            I => \N__21690\
        );

    \I__3443\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21687\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__21690\,
            I => \N__21681\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21678\
        );

    \I__3440\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21671\
        );

    \I__3439\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21671\
        );

    \I__3438\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21671\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__21681\,
            I => \N__21668\
        );

    \I__3436\ : Sp12to4
    port map (
            O => \N__21678\,
            I => \N__21663\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21663\
        );

    \I__3434\ : Sp12to4
    port map (
            O => \N__21668\,
            I => \N__21658\
        );

    \I__3433\ : Span12Mux_v
    port map (
            O => \N__21663\,
            I => \N__21658\
        );

    \I__3432\ : Odrv12
    port map (
            O => \N__21658\,
            I => vddq_ok
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__3430\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21643\
        );

    \I__3429\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21643\
        );

    \I__3428\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21643\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__21643\,
            I => \VPP_VDDQ.N_2897_i\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__3425\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21633\
        );

    \I__3424\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21630\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__21633\,
            I => \VPP_VDDQ.N_297_0\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__21630\,
            I => \VPP_VDDQ.N_297_0\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__21625\,
            I => \POWERLED.un79_clk_100khzlto15_5_cascade_\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__21622\,
            I => \POWERLED.un79_clk_100khzlto15_7_cascade_\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__21619\,
            I => \POWERLED.un79_clk_100khzlt6_cascade_\
        );

    \I__3418\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__21613\,
            I => \POWERLED.un79_clk_100khzlto15_3\
        );

    \I__3416\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__21604\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__3413\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21598\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__21595\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__3410\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__21589\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__3408\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__21583\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__3406\ : InMux
    port map (
            O => \N__21580\,
            I => \bfn_6_7_0_\
        );

    \I__3405\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21574\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__21574\,
            I => \N__21571\
        );

    \I__3403\ : Odrv12
    port map (
            O => \N__21571\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__3401\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21561\
        );

    \I__3400\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21556\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21553\
        );

    \I__3398\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21548\
        );

    \I__3397\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21548\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__21556\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__21553\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__21548\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__21541\,
            I => \DSW_PWRGD.un4_count_11_cascade_\
        );

    \I__3392\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21535\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__21535\,
            I => \DSW_PWRGD.un4_count_10\
        );

    \I__3390\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__21529\,
            I => \DSW_PWRGD.un4_count_8\
        );

    \I__3388\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21523\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__21523\,
            I => \N__21520\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__21520\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__3385\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21514\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__21514\,
            I => \N__21511\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__21511\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__3382\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__21502\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__3379\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21496\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__3377\ : Odrv12
    port map (
            O => \N__21493\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__3376\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21486\
        );

    \I__3375\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21483\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__21486\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__21483\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3372\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21474\
        );

    \I__3371\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21471\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__21474\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__21471\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__21466\,
            I => \N__21462\
        );

    \I__3367\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21459\
        );

    \I__3366\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21456\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__21459\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__21456\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3363\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21447\
        );

    \I__3362\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21444\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__21447\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__21444\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3359\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21435\
        );

    \I__3358\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21432\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__21435\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__21432\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__21427\,
            I => \N__21423\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__21426\,
            I => \N__21419\
        );

    \I__3353\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21416\
        );

    \I__3352\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21411\
        );

    \I__3351\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21411\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__21416\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__21411\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3348\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21401\
        );

    \I__3347\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21396\
        );

    \I__3346\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21396\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__21401\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__21396\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3343\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21388\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__21388\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__3341\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21380\
        );

    \I__3340\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21375\
        );

    \I__3339\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21375\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__21380\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__21375\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3336\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21367\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21364\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__21364\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__3333\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21358\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__21358\,
            I => \N__21353\
        );

    \I__3331\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21348\
        );

    \I__3330\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21348\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__21353\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__21348\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3327\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21338\
        );

    \I__3326\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21335\
        );

    \I__3325\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21332\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__21338\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__21335\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__21332\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3321\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21321\
        );

    \I__3320\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21318\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__21321\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__21318\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3317\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21309\
        );

    \I__3316\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21306\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__21309\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__21306\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__21301\,
            I => \N__21297\
        );

    \I__3312\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21294\
        );

    \I__3311\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21291\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__21294\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__21291\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3308\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21282\
        );

    \I__3307\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21279\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__21282\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__21279\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3304\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21270\
        );

    \I__3303\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21267\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__21270\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__21267\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3300\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21258\
        );

    \I__3299\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21255\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__21258\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__21255\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__21250\,
            I => \N__21246\
        );

    \I__3295\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21243\
        );

    \I__3294\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21240\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__21243\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__21240\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3291\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21231\
        );

    \I__3290\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21228\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__21231\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__21228\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3287\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21220\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__21220\,
            I => \N__21217\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__21217\,
            I => \N__21214\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__21214\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__3283\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21207\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__21210\,
            I => \N__21203\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21200\
        );

    \I__3280\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21195\
        );

    \I__3279\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21195\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__21200\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__21195\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__21190\,
            I => \N__21187\
        );

    \I__3275\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21178\
        );

    \I__3274\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21178\
        );

    \I__3273\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21178\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__21178\,
            I => \HDA_STRAP.N_285\
        );

    \I__3271\ : InMux
    port map (
            O => \N__21175\,
            I => \N__21168\
        );

    \I__3270\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21161\
        );

    \I__3269\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21161\
        );

    \I__3268\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21161\
        );

    \I__3267\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21158\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__21168\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__21161\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__21158\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__21151\,
            I => \HDA_STRAP.N_285_cascade_\
        );

    \I__3262\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21145\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__21145\,
            I => \HDA_STRAP.N_51\
        );

    \I__3260\ : IoInMux
    port map (
            O => \N__21142\,
            I => \N__21139\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__21139\,
            I => \N__21136\
        );

    \I__3258\ : Odrv12
    port map (
            O => \N__21136\,
            I => vccst_pwrgd
        );

    \I__3257\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21130\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21127\
        );

    \I__3255\ : Span4Mux_s2_v
    port map (
            O => \N__21127\,
            I => \N__21124\
        );

    \I__3254\ : Odrv4
    port map (
            O => \N__21124\,
            I => \PCH_PWRGD.delayed_vccin_okZ0\
        );

    \I__3253\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21113\
        );

    \I__3252\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21106\
        );

    \I__3251\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21106\
        );

    \I__3250\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21106\
        );

    \I__3249\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21101\
        );

    \I__3248\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21101\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N_227\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__21106\,
            I => \N_227\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N_227\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__21094\,
            I => \N_227_cascade_\
        );

    \I__3243\ : IoInMux
    port map (
            O => \N__21091\,
            I => \N__21088\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__21088\,
            I => \N__21085\
        );

    \I__3241\ : Span4Mux_s1_h
    port map (
            O => \N__21085\,
            I => \N__21082\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__21082\,
            I => \N__21079\
        );

    \I__3239\ : Sp12to4
    port map (
            O => \N__21079\,
            I => \N__21075\
        );

    \I__3238\ : IoInMux
    port map (
            O => \N__21078\,
            I => \N__21072\
        );

    \I__3237\ : Span12Mux_v
    port map (
            O => \N__21075\,
            I => \N__21067\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__21067\
        );

    \I__3235\ : Odrv12
    port map (
            O => \N__21067\,
            I => pch_pwrok
        );

    \I__3234\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21060\
        );

    \I__3233\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21057\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__21060\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__21057\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3230\ : InMux
    port map (
            O => \N__21052\,
            I => \N__21048\
        );

    \I__3229\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21045\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__21048\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__21045\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__21040\,
            I => \N__21036\
        );

    \I__3225\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21033\
        );

    \I__3224\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21030\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__21033\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__21030\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3221\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21021\
        );

    \I__3220\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21018\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__21021\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__21018\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3217\ : InMux
    port map (
            O => \N__21013\,
            I => \N__21010\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__21010\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__3215\ : InMux
    port map (
            O => \N__21007\,
            I => \N__21004\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__21004\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__21001\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__20998\,
            I => \POWERLED.un1_dutycycle_53_10_0_cascade_\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__20995\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_12_cascade_\
        );

    \I__3210\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20989\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__20989\,
            I => \POWERLED.un1_dutycycle_53_10_2\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__20986\,
            I => \N_414_cascade_\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__20983\,
            I => \N__20980\
        );

    \I__3206\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20977\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__20977\,
            I => \N__20974\
        );

    \I__3204\ : Span4Mux_h
    port map (
            O => \N__20974\,
            I => \N__20971\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__20971\,
            I => gpio_fpga_soc_1
        );

    \I__3202\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20965\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__20965\,
            I => \HDA_STRAP.m6_i_0\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__20962\,
            I => \HDA_STRAP.m6_i_0_cascade_\
        );

    \I__3199\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20956\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__20956\,
            I => \HDA_STRAP.curr_state_3_0\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__20953\,
            I => \HDA_STRAP.N_53_cascade_\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__20950\,
            I => \POWERLED.dutycycle_1_0_0_cascade_\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20944\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__20944\,
            I => \POWERLED.dutycycle_1_0_0\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20937\
        );

    \I__3192\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20934\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20929\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20929\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__20929\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__3188\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20922\
        );

    \I__3187\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20919\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__20922\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__20919\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__20914\,
            I => \N__20911\
        );

    \I__3183\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20904\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__20910\,
            I => \N__20899\
        );

    \I__3181\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20893\
        );

    \I__3180\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20893\
        );

    \I__3179\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20890\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20884\
        );

    \I__3177\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20879\
        );

    \I__3176\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20879\
        );

    \I__3175\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20874\
        );

    \I__3174\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20874\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20867\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__20890\,
            I => \N__20867\
        );

    \I__3171\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20863\
        );

    \I__3170\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20857\
        );

    \I__3169\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20857\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__20884\,
            I => \N__20850\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20850\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__20874\,
            I => \N__20850\
        );

    \I__3165\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20845\
        );

    \I__3164\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20845\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__20867\,
            I => \N__20842\
        );

    \I__3162\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20839\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__20863\,
            I => \N__20836\
        );

    \I__3160\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20833\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__20857\,
            I => \N__20830\
        );

    \I__3158\ : Span4Mux_v
    port map (
            O => \N__20850\,
            I => \N__20827\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20814\
        );

    \I__3156\ : Sp12to4
    port map (
            O => \N__20842\,
            I => \N__20814\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__20839\,
            I => \N__20814\
        );

    \I__3154\ : Span12Mux_s4_h
    port map (
            O => \N__20836\,
            I => \N__20814\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20814\
        );

    \I__3152\ : Span12Mux_s2_v
    port map (
            O => \N__20830\,
            I => \N__20814\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__20827\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3150\ : Odrv12
    port map (
            O => \N__20814\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3149\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20806\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__20806\,
            I => \POWERLED.dutycycle_1_0_1\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__20803\,
            I => \N__20799\
        );

    \I__3146\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20794\
        );

    \I__3145\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20794\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__20794\,
            I => \N__20791\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__20791\,
            I => \POWERLED.dutycycle_eena_0\
        );

    \I__3142\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20782\
        );

    \I__3141\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20782\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__20782\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__20779\,
            I => \POWERLED.dutycycle_1_0_1_cascade_\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__3137\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20770\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__20770\,
            I => \POWERLED.dutycycle_eena_7\
        );

    \I__3135\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20761\
        );

    \I__3134\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20761\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__20761\,
            I => \POWERLED.dutycycleZ1Z_11\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__20758\,
            I => \POWERLED.dutycycle_eena_7_cascade_\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \POWERLED.dutycycleZ0Z_8_cascade_\
        );

    \I__3130\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__20749\,
            I => \POWERLED.N_12\
        );

    \I__3128\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__20743\,
            I => \POWERLED.g0_i_a6_1\
        );

    \I__3126\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20737\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__20737\,
            I => \POWERLED.N_358\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__20734\,
            I => \POWERLED.un1_clk_100khz_42_and_i_a2_3_0_cascade_\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__20731\,
            I => \POWERLED.N_434_N_cascade_\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__20728\,
            I => \N__20721\
        );

    \I__3121\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20716\
        );

    \I__3120\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20713\
        );

    \I__3119\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20708\
        );

    \I__3118\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20708\
        );

    \I__3117\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20701\
        );

    \I__3116\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20701\
        );

    \I__3115\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20701\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20698\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__20713\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__20708\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__20701\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__20698\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__20689\,
            I => \POWERLED.N_372_cascade_\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__20686\,
            I => \POWERLED.N_122_f0_1_cascade_\
        );

    \I__3107\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__20680\,
            I => \POWERLED.N_122_f0_1\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__20677\,
            I => \POWERLED.g0_i_a6_1_1_cascade_\
        );

    \I__3104\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__20671\,
            I => \POWERLED.N_10_0\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__20668\,
            I => \tmp_1_rep1_RNI_cascade_\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__20665\,
            I => \POWERLED.N_358_cascade_\
        );

    \I__3100\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20659\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20656\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__20656\,
            I => \N__20653\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__20653\,
            I => \POWERLED.func_state_1_m2s2_i_0\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \POWERLED.N_344_cascade_\
        );

    \I__3095\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__20644\,
            I => \POWERLED.N_343\
        );

    \I__3093\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__20638\,
            I => \POWERLED.N_79\
        );

    \I__3091\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20629\
        );

    \I__3089\ : Span4Mux_v
    port map (
            O => \N__20629\,
            I => \N__20624\
        );

    \I__3088\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20619\
        );

    \I__3087\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20619\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__20624\,
            I => \POWERLED.func_state_RNI3IN21Z0Z_0\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__20619\,
            I => \POWERLED.func_state_RNI3IN21Z0Z_0\
        );

    \I__3084\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20611\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__20611\,
            I => \POWERLED.N_433\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__20608\,
            I => \POWERLED.N_79_cascade_\
        );

    \I__3081\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20602\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__20602\,
            I => \N__20599\
        );

    \I__3079\ : Span4Mux_v
    port map (
            O => \N__20599\,
            I => \N__20596\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__20596\,
            I => \POWERLED.func_state_1_m2_ns_1_0\
        );

    \I__3077\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20587\
        );

    \I__3076\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20587\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__20587\,
            I => \N__20584\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__20581\,
            I => \POWERLED.func_state_1_m2_0\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__20575\,
            I => \N__20572\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__20572\,
            I => \N__20569\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__20569\,
            I => \POWERLED.un1_func_state25_6_0_2\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__20566\,
            I => \POWERLED.un1_func_state25_6_0_a3_1_cascade_\
        );

    \I__3067\ : CEMux
    port map (
            O => \N__20563\,
            I => \N__20558\
        );

    \I__3066\ : CEMux
    port map (
            O => \N__20562\,
            I => \N__20555\
        );

    \I__3065\ : CEMux
    port map (
            O => \N__20561\,
            I => \N__20552\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__20558\,
            I => \N__20547\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20547\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20542\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__20547\,
            I => \N__20539\
        );

    \I__3060\ : CEMux
    port map (
            O => \N__20546\,
            I => \N__20536\
        );

    \I__3059\ : CEMux
    port map (
            O => \N__20545\,
            I => \N__20528\
        );

    \I__3058\ : Span4Mux_h
    port map (
            O => \N__20542\,
            I => \N__20521\
        );

    \I__3057\ : Span4Mux_h
    port map (
            O => \N__20539\,
            I => \N__20521\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20521\
        );

    \I__3055\ : CEMux
    port map (
            O => \N__20535\,
            I => \N__20515\
        );

    \I__3054\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20502\
        );

    \I__3053\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20502\
        );

    \I__3052\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20502\
        );

    \I__3051\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20502\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20497\
        );

    \I__3049\ : Span4Mux_v
    port map (
            O => \N__20521\,
            I => \N__20494\
        );

    \I__3048\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20487\
        );

    \I__3047\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20487\
        );

    \I__3046\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20487\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20481\
        );

    \I__3044\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20472\
        );

    \I__3043\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20472\
        );

    \I__3042\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20472\
        );

    \I__3041\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20472\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20469\
        );

    \I__3039\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20466\
        );

    \I__3038\ : InMux
    port map (
            O => \N__20500\,
            I => \N__20463\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__20497\,
            I => \N__20456\
        );

    \I__3036\ : Span4Mux_s0_v
    port map (
            O => \N__20494\,
            I => \N__20456\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__20487\,
            I => \N__20456\
        );

    \I__3034\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20449\
        );

    \I__3033\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20449\
        );

    \I__3032\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20449\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__20481\,
            I => \N__20446\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__20472\,
            I => \N__20437\
        );

    \I__3029\ : Span4Mux_s2_h
    port map (
            O => \N__20469\,
            I => \N__20437\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__20466\,
            I => \N__20437\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__20463\,
            I => \N__20437\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__20456\,
            I => \N__20432\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20432\
        );

    \I__3024\ : Span4Mux_s2_h
    port map (
            O => \N__20446\,
            I => \N__20427\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__20437\,
            I => \N__20427\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__20432\,
            I => \POWERLED.dutycycle_RNIH0LB7Z0Z_0\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__20427\,
            I => \POWERLED.dutycycle_RNIH0LB7Z0Z_0\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__20422\,
            I => \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__20419\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__3018\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__20413\,
            I => \N__20410\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__20410\,
            I => \N__20407\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__20407\,
            I => \POWERLED.N_189_i\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__20404\,
            I => \POWERLED.N_189_i_cascade_\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__20401\,
            I => \POWERLED.N_331_N_0_0_cascade_\
        );

    \I__3012\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__20395\,
            I => \POWERLED.g3_1_0_1\
        );

    \I__3010\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__3008\ : Span4Mux_s3_v
    port map (
            O => \N__20386\,
            I => \N__20383\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__20383\,
            I => \POWERLED.g3_1_0\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__20380\,
            I => \POWERLED.func_m1_0_a2Z0Z_0_cascade_\
        );

    \I__3005\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__20374\,
            I => \POWERLED.func_state_1_ss0_i_0_o2_1\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__20371\,
            I => \POWERLED.N_433_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20365\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__20365\,
            I => \POWERLED.func_state_1_m2_ns_1_1\
        );

    \I__3000\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20356\
        );

    \I__2999\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20356\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__20356\,
            I => \POWERLED.func_state_1_m2_1\
        );

    \I__2997\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20350\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__20350\,
            I => \POWERLED.N_345\
        );

    \I__2995\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20336\
        );

    \I__2994\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20336\
        );

    \I__2993\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20336\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__20344\,
            I => \N__20332\
        );

    \I__2991\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20328\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20324\
        );

    \I__2989\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20319\
        );

    \I__2988\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20319\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__20331\,
            I => \N__20314\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20311\
        );

    \I__2985\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20308\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__20324\,
            I => \N__20304\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__20319\,
            I => \N__20301\
        );

    \I__2982\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20294\
        );

    \I__2981\ : InMux
    port map (
            O => \N__20317\,
            I => \N__20294\
        );

    \I__2980\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20294\
        );

    \I__2979\ : Span4Mux_h
    port map (
            O => \N__20311\,
            I => \N__20289\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__20308\,
            I => \N__20289\
        );

    \I__2977\ : InMux
    port map (
            O => \N__20307\,
            I => \N__20286\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__20304\,
            I => \POWERLED.N_164\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__20301\,
            I => \POWERLED.N_164\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__20294\,
            I => \POWERLED.N_164\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__20289\,
            I => \POWERLED.N_164\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__20286\,
            I => \POWERLED.N_164\
        );

    \I__2971\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20271\
        );

    \I__2970\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20268\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__20271\,
            I => \N__20265\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__20268\,
            I => \N__20260\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__20265\,
            I => \N__20260\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__20260\,
            I => \POWERLED.count_1_13\
        );

    \I__2965\ : InMux
    port map (
            O => \N__20257\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__2964\ : InMux
    port map (
            O => \N__20254\,
            I => \POWERLED.un1_count_cry_13\
        );

    \I__2963\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20235\
        );

    \I__2962\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20235\
        );

    \I__2961\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20235\
        );

    \I__2960\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20235\
        );

    \I__2959\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20228\
        );

    \I__2958\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20228\
        );

    \I__2957\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20228\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__20244\,
            I => \N__20216\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20211\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__20228\,
            I => \N__20211\
        );

    \I__2953\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20202\
        );

    \I__2952\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20202\
        );

    \I__2951\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20202\
        );

    \I__2950\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20202\
        );

    \I__2949\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20195\
        );

    \I__2948\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20195\
        );

    \I__2947\ : InMux
    port map (
            O => \N__20221\,
            I => \N__20195\
        );

    \I__2946\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20188\
        );

    \I__2945\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20188\
        );

    \I__2944\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20188\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__20211\,
            I => \N__20185\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20180\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20180\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__20188\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__20185\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__20180\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2937\ : InMux
    port map (
            O => \N__20173\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__2936\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20167\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__20167\,
            I => \N__20163\
        );

    \I__2934\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20160\
        );

    \I__2933\ : Odrv12
    port map (
            O => \N__20163\,
            I => \POWERLED.count_1_14\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__20160\,
            I => \POWERLED.count_1_14\
        );

    \I__2931\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20152\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__20152\,
            I => \N__20149\
        );

    \I__2929\ : Odrv12
    port map (
            O => \N__20149\,
            I => \POWERLED.count_0_14\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__20146\,
            I => \POWERLED.N_8_2_cascade_\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__20143\,
            I => \POWERLED.N_5_0_cascade_\
        );

    \I__2926\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20137\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__20137\,
            I => \POWERLED.g0_5_0\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__20134\,
            I => \N__20130\
        );

    \I__2923\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20127\
        );

    \I__2922\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20124\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__20127\,
            I => \N__20121\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__20124\,
            I => \POWERLED.count_1_4\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__20121\,
            I => \POWERLED.count_1_4\
        );

    \I__2918\ : InMux
    port map (
            O => \N__20116\,
            I => \POWERLED.un1_count_cry_3\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__2916\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20106\
        );

    \I__2915\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20103\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__20106\,
            I => \N__20100\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__20103\,
            I => \POWERLED.count_1_5\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__20100\,
            I => \POWERLED.count_1_5\
        );

    \I__2911\ : InMux
    port map (
            O => \N__20095\,
            I => \POWERLED.un1_count_cry_4\
        );

    \I__2910\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20088\
        );

    \I__2909\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20085\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N__20082\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__20085\,
            I => \POWERLED.count_1_6\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__20082\,
            I => \POWERLED.count_1_6\
        );

    \I__2905\ : InMux
    port map (
            O => \N__20077\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__2904\ : InMux
    port map (
            O => \N__20074\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__2903\ : InMux
    port map (
            O => \N__20071\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__2902\ : InMux
    port map (
            O => \N__20068\,
            I => \bfn_5_9_0_\
        );

    \I__2901\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20059\
        );

    \I__2900\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20059\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__20059\,
            I => \POWERLED.count_1_10\
        );

    \I__2898\ : InMux
    port map (
            O => \N__20056\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__2897\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20050\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__20050\,
            I => \N__20046\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__20049\,
            I => \N__20043\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__20046\,
            I => \N__20040\
        );

    \I__2893\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20037\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__20040\,
            I => \POWERLED.count_1_11\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__20037\,
            I => \POWERLED.count_1_11\
        );

    \I__2890\ : InMux
    port map (
            O => \N__20032\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__2889\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20023\
        );

    \I__2888\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20023\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__20023\,
            I => \POWERLED.count_1_12\
        );

    \I__2886\ : InMux
    port map (
            O => \N__20020\,
            I => \POWERLED.un1_count_cry_11\
        );

    \I__2885\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__20011\,
            I => \N__20008\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__20008\,
            I => \POWERLED.count_0_4\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__20005\,
            I => \N__20001\
        );

    \I__2880\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19995\
        );

    \I__2879\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19995\
        );

    \I__2878\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19992\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__19995\,
            I => \N__19987\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19987\
        );

    \I__2875\ : Span4Mux_h
    port map (
            O => \N__19987\,
            I => \N__19984\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__19984\,
            I => \RSMRST_PWRGD.N_423\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__19981\,
            I => \N__19969\
        );

    \I__2872\ : SRMux
    port map (
            O => \N__19980\,
            I => \N__19962\
        );

    \I__2871\ : SRMux
    port map (
            O => \N__19979\,
            I => \N__19958\
        );

    \I__2870\ : SRMux
    port map (
            O => \N__19978\,
            I => \N__19955\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__19977\,
            I => \N__19952\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__19976\,
            I => \N__19941\
        );

    \I__2867\ : SRMux
    port map (
            O => \N__19975\,
            I => \N__19935\
        );

    \I__2866\ : SRMux
    port map (
            O => \N__19974\,
            I => \N__19932\
        );

    \I__2865\ : SRMux
    port map (
            O => \N__19973\,
            I => \N__19929\
        );

    \I__2864\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19924\
        );

    \I__2863\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19924\
        );

    \I__2862\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19915\
        );

    \I__2861\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19915\
        );

    \I__2860\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19915\
        );

    \I__2859\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19915\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__19962\,
            I => \N__19910\
        );

    \I__2857\ : SRMux
    port map (
            O => \N__19961\,
            I => \N__19907\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19902\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__19955\,
            I => \N__19902\
        );

    \I__2854\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19888\
        );

    \I__2853\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19888\
        );

    \I__2852\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19888\
        );

    \I__2851\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19888\
        );

    \I__2850\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19888\
        );

    \I__2849\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19881\
        );

    \I__2848\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19881\
        );

    \I__2847\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19881\
        );

    \I__2846\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19874\
        );

    \I__2845\ : InMux
    port map (
            O => \N__19941\,
            I => \N__19874\
        );

    \I__2844\ : InMux
    port map (
            O => \N__19940\,
            I => \N__19874\
        );

    \I__2843\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19869\
        );

    \I__2842\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19869\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19866\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__19932\,
            I => \N__19857\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19857\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__19924\,
            I => \N__19857\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19857\
        );

    \I__2836\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19854\
        );

    \I__2835\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19851\
        );

    \I__2834\ : Span4Mux_s1_h
    port map (
            O => \N__19910\,
            I => \N__19846\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19846\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__19902\,
            I => \N__19843\
        );

    \I__2831\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19836\
        );

    \I__2830\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19836\
        );

    \I__2829\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19836\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__19888\,
            I => \N__19833\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__19881\,
            I => \N__19830\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__19874\,
            I => \N__19825\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__19869\,
            I => \N__19825\
        );

    \I__2824\ : Span4Mux_h
    port map (
            O => \N__19866\,
            I => \N__19822\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__19857\,
            I => \N__19817\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19817\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19814\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__19846\,
            I => \N__19805\
        );

    \I__2819\ : Span4Mux_s1_h
    port map (
            O => \N__19843\,
            I => \N__19805\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__19836\,
            I => \N__19805\
        );

    \I__2817\ : Span4Mux_v
    port map (
            O => \N__19833\,
            I => \N__19805\
        );

    \I__2816\ : Span12Mux_s4_h
    port map (
            O => \N__19830\,
            I => \N__19802\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__19825\,
            I => \N__19799\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__19822\,
            I => \N__19794\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__19817\,
            I => \N__19794\
        );

    \I__2812\ : Odrv12
    port map (
            O => \N__19814\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__19805\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2810\ : Odrv12
    port map (
            O => \N__19802\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__19799\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__19794\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2807\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__19777\,
            I => \POWERLED.count_0_13\
        );

    \I__2804\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__19768\,
            I => \POWERLED.count_0_5\
        );

    \I__2801\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__2799\ : Span4Mux_v
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__19756\,
            I => \POWERLED.count_0_6\
        );

    \I__2797\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19749\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__19752\,
            I => \N__19746\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__19749\,
            I => \N__19743\
        );

    \I__2794\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19740\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__19743\,
            I => \POWERLED.count_1_2\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__19740\,
            I => \POWERLED.count_1_2\
        );

    \I__2791\ : InMux
    port map (
            O => \N__19735\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__2790\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19726\
        );

    \I__2789\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19726\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__19726\,
            I => \POWERLED.count_1_3\
        );

    \I__2787\ : InMux
    port map (
            O => \N__19723\,
            I => \POWERLED.un1_count_cry_2\
        );

    \I__2786\ : InMux
    port map (
            O => \N__19720\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__2785\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19711\
        );

    \I__2784\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19711\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__19711\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__19708\,
            I => \N__19705\
        );

    \I__2781\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19699\
        );

    \I__2780\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19699\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__19699\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__19696\,
            I => \N__19692\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__19695\,
            I => \N__19689\
        );

    \I__2776\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19684\
        );

    \I__2775\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19684\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__19684\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2773\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19677\
        );

    \I__2772\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19674\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__19677\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__19674\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__19669\,
            I => \N__19665\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__19668\,
            I => \N__19661\
        );

    \I__2767\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19655\
        );

    \I__2766\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19655\
        );

    \I__2765\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19650\
        );

    \I__2764\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19650\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19647\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__19650\,
            I => \N__19644\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__19647\,
            I => \N__19641\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__19644\,
            I => \N__19638\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__19641\,
            I => \N__19635\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__19638\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__19635\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__19630\,
            I => \N__19626\
        );

    \I__2755\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19621\
        );

    \I__2754\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19621\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__19621\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__2752\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19614\
        );

    \I__2751\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19611\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__19614\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__19611\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2748\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19602\
        );

    \I__2747\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19599\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__19602\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__19599\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__19594\,
            I => \N__19590\
        );

    \I__2743\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19587\
        );

    \I__2742\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19584\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__19587\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__19584\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2739\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19575\
        );

    \I__2738\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19572\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__19575\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__19572\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__19567\,
            I => \VPP_VDDQ.N_2897_i_cascade_\
        );

    \I__2734\ : InMux
    port map (
            O => \N__19564\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__2733\ : InMux
    port map (
            O => \N__19561\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__2732\ : InMux
    port map (
            O => \N__19558\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__2731\ : InMux
    port map (
            O => \N__19555\,
            I => \bfn_5_5_0_\
        );

    \I__2730\ : InMux
    port map (
            O => \N__19552\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__2729\ : InMux
    port map (
            O => \N__19549\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__2728\ : InMux
    port map (
            O => \N__19546\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__2727\ : InMux
    port map (
            O => \N__19543\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__2726\ : InMux
    port map (
            O => \N__19540\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__2725\ : InMux
    port map (
            O => \N__19537\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__2724\ : InMux
    port map (
            O => \N__19534\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__2723\ : InMux
    port map (
            O => \N__19531\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__2722\ : InMux
    port map (
            O => \N__19528\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__2721\ : InMux
    port map (
            O => \N__19525\,
            I => \bfn_5_4_0_\
        );

    \I__2720\ : InMux
    port map (
            O => \N__19522\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__2719\ : InMux
    port map (
            O => \N__19519\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__2718\ : InMux
    port map (
            O => \N__19516\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__2717\ : InMux
    port map (
            O => \N__19513\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__2716\ : InMux
    port map (
            O => \N__19510\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__2715\ : InMux
    port map (
            O => \N__19507\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__2714\ : InMux
    port map (
            O => \N__19504\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__2713\ : InMux
    port map (
            O => \N__19501\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__2712\ : InMux
    port map (
            O => \N__19498\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__2711\ : InMux
    port map (
            O => \N__19495\,
            I => \bfn_5_3_0_\
        );

    \I__2710\ : InMux
    port map (
            O => \N__19492\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__2709\ : InMux
    port map (
            O => \N__19489\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__2708\ : InMux
    port map (
            O => \N__19486\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__2707\ : IoInMux
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19477\
        );

    \I__2705\ : Span4Mux_s0_h
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__19468\,
            I => hda_sdo_atp
        );

    \I__2701\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19462\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__19462\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \HDA_STRAP.curr_state_i_2_cascade_\
        );

    \I__2698\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19453\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__19453\,
            I => \HDA_STRAP.i4_mux\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__19450\,
            I => \N__19447\
        );

    \I__2695\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19438\
        );

    \I__2694\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19438\
        );

    \I__2693\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19438\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__19438\,
            I => \HDA_STRAP.N_208\
        );

    \I__2691\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19426\
        );

    \I__2690\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19426\
        );

    \I__2689\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19426\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__19426\,
            I => \HDA_STRAP.curr_state_i_2\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__19423\,
            I => \HDA_STRAP.N_208_cascade_\
        );

    \I__2686\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19417\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__19417\,
            I => \HDA_STRAP.HDA_SDO_ATP_0\
        );

    \I__2684\ : InMux
    port map (
            O => \N__19414\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__2683\ : InMux
    port map (
            O => \N__19411\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__2682\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__2681\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19402\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__2679\ : Span4Mux_s2_v
    port map (
            O => \N__19399\,
            I => \N__19396\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__19396\,
            I => \POWERLED.count_off_1_6\
        );

    \I__2677\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19390\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__19390\,
            I => \POWERLED.count_off_0_6\
        );

    \I__2675\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19383\
        );

    \I__2674\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19380\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19377\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__19380\,
            I => \N__19374\
        );

    \I__2671\ : Span4Mux_s3_h
    port map (
            O => \N__19377\,
            I => \N__19371\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__19374\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__19371\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2668\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__2667\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19360\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__19360\,
            I => \N__19357\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__19354\,
            I => \POWERLED.count_off_1_7\
        );

    \I__2663\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19348\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__19348\,
            I => \POWERLED.count_off_0_7\
        );

    \I__2661\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19341\
        );

    \I__2660\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19338\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__19341\,
            I => \N__19335\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__19338\,
            I => \N__19332\
        );

    \I__2657\ : Span4Mux_s3_h
    port map (
            O => \N__19335\,
            I => \N__19329\
        );

    \I__2656\ : Odrv12
    port map (
            O => \N__19332\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__19329\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__2654\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__2653\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19318\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__19318\,
            I => \N__19315\
        );

    \I__2651\ : Span4Mux_s2_v
    port map (
            O => \N__19315\,
            I => \N__19312\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__19312\,
            I => \POWERLED.count_off_1_8\
        );

    \I__2649\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__19306\,
            I => \POWERLED.count_off_0_8\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__19303\,
            I => \HDA_STRAP.curr_stateZ0Z_1_cascade_\
        );

    \I__2646\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19297\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__19297\,
            I => \HDA_STRAP.curr_state_2_1\
        );

    \I__2644\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__19291\,
            I => \POWERLED.N_5_1\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__19288\,
            I => \POWERLED.g0_i_a6_0_1_cascade_\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__19285\,
            I => \POWERLED.g2_1_0_0_cascade_\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__19282\,
            I => \POWERLED.dutycycle_en_5_0_0_cascade_\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__19279\,
            I => \POWERLED.dutycycleZ0Z_5_cascade_\
        );

    \I__2638\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19273\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__19273\,
            I => \POWERLED.dutycycle_eena_5_0_N_3_1\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__19270\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_7_cascade_\
        );

    \I__2635\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__19264\,
            I => \POWERLED.g0_i_1\
        );

    \I__2633\ : InMux
    port map (
            O => \N__19261\,
            I => \N__19258\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__19258\,
            I => \POWERLED.dutycycle_en_5_0_0\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \N__19252\
        );

    \I__2630\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19246\
        );

    \I__2629\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19246\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__19246\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__2627\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19239\
        );

    \I__2626\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19236\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__19239\,
            I => \N__19233\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19228\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__19233\,
            I => \N__19228\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__19228\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__19225\,
            I => \N__19221\
        );

    \I__2620\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19216\
        );

    \I__2619\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19216\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__19216\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__2616\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19207\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19204\
        );

    \I__2614\ : Span12Mux_s4_v
    port map (
            O => \N__19204\,
            I => \N__19201\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__19201\,
            I => \POWERLED.N_301\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__19198\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__19195\,
            I => \POWERLED.N_238_cascade_\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__19192\,
            I => \POWERLED.N_118_f0_cascade_\
        );

    \I__2609\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19186\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__19186\,
            I => \POWERLED.dutycycle_RNIS3763Z0Z_2\
        );

    \I__2607\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19177\
        );

    \I__2606\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19177\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__19177\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__2604\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__2603\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19168\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__19168\,
            I => \N__19165\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__19165\,
            I => \POWERLED.N_171\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__19162\,
            I => \POWERLED.dutycycle_RNIS3763Z0Z_2_cascade_\
        );

    \I__2599\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19156\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__19156\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_2\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__19153\,
            I => \POWERLED.dutycycle_cascade_\
        );

    \I__2596\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19143\
        );

    \I__2595\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19143\
        );

    \I__2594\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19140\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__19143\,
            I => \POWERLED.func_state_1_ss0_i_0_a2Z0Z_3\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__19140\,
            I => \POWERLED.func_state_1_ss0_i_0_a2Z0Z_3\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__19135\,
            I => \POWERLED.func_state_cascade_\
        );

    \I__2590\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19129\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__19129\,
            I => \N__19125\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__19128\,
            I => \N__19122\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__19125\,
            I => \N__19119\
        );

    \I__2586\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19116\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__19119\,
            I => \POWERLED.func_state_RNI_4Z0Z_1\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__19116\,
            I => \POWERLED.func_state_RNI_4Z0Z_1\
        );

    \I__2583\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__19102\,
            I => \POWERLED.un1_func_state25_6_0_a2_1\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\
        );

    \I__2578\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__19087\,
            I => vpp_ok
        );

    \I__2574\ : IoInMux
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__2572\ : IoSpan4Mux
    port map (
            O => \N__19078\,
            I => \N__19075\
        );

    \I__2571\ : Span4Mux_s1_v
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__19072\,
            I => vddq_en
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \POWERLED.N_171_cascade_\
        );

    \I__2568\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__2567\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19060\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__19060\,
            I => \N__19057\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__19057\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_oZ0Z3\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__19054\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3_out_cascade_\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__19051\,
            I => \POWERLED.func_state_RNI3IN21Z0Z_0_cascade_\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__19048\,
            I => \POWERLED.func_state_1_m2_ns_1_1_1_cascade_\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \POWERLED.N_2905_i_cascade_\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__19042\,
            I => \POWERLED.N_175_cascade_\
        );

    \I__2559\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19035\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__19038\,
            I => \N__19032\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__19029\
        );

    \I__2556\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19024\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__19029\,
            I => \N__19021\
        );

    \I__2554\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19018\
        );

    \I__2553\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19015\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__19024\,
            I => \N__19012\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__19021\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__19018\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__19015\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__19012\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__2547\ : InMux
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__19000\,
            I => \N__18997\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__18994\,
            I => \POWERLED.count_clk_RNIZ0Z_0\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__18991\,
            I => \N__18988\
        );

    \I__2542\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18985\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__18985\,
            I => \N__18982\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__18982\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0\
        );

    \I__2539\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__18970\,
            I => \POWERLED.count_off_0_2\
        );

    \I__2535\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18964\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18961\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__18961\,
            I => \N__18958\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__18958\,
            I => \N__18954\
        );

    \I__2531\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18951\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__18954\,
            I => \POWERLED.count_off_1_2\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__18951\,
            I => \POWERLED.count_off_1_2\
        );

    \I__2528\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18943\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__18943\,
            I => \N__18939\
        );

    \I__2526\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18936\
        );

    \I__2525\ : Span4Mux_s3_h
    port map (
            O => \N__18939\,
            I => \N__18933\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__18936\,
            I => \N__18930\
        );

    \I__2523\ : Sp12to4
    port map (
            O => \N__18933\,
            I => \N__18925\
        );

    \I__2522\ : Span12Mux_s3_h
    port map (
            O => \N__18930\,
            I => \N__18925\
        );

    \I__2521\ : Odrv12
    port map (
            O => \N__18925\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__2520\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18919\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__18919\,
            I => \N__18916\
        );

    \I__2518\ : Span4Mux_h
    port map (
            O => \N__18916\,
            I => \N__18913\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__18913\,
            I => \POWERLED.count_off_0_3\
        );

    \I__2516\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18907\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18904\
        );

    \I__2514\ : Span4Mux_h
    port map (
            O => \N__18904\,
            I => \N__18901\
        );

    \I__2513\ : Span4Mux_v
    port map (
            O => \N__18901\,
            I => \N__18897\
        );

    \I__2512\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18894\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__18897\,
            I => \POWERLED.count_off_1_3\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__18894\,
            I => \POWERLED.count_off_1_3\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__18889\,
            I => \N__18886\
        );

    \I__2508\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18882\
        );

    \I__2507\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18879\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__18882\,
            I => \N__18876\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__18879\,
            I => \N__18873\
        );

    \I__2504\ : Span4Mux_s3_v
    port map (
            O => \N__18876\,
            I => \N__18870\
        );

    \I__2503\ : Span4Mux_s3_h
    port map (
            O => \N__18873\,
            I => \N__18867\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__18870\,
            I => \N__18864\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__18867\,
            I => \N__18861\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__18864\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__18861\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__18856\,
            I => \N__18853\
        );

    \I__2497\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18850\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__18850\,
            I => \N__18847\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__18844\,
            I => \POWERLED.count_off_0_4\
        );

    \I__2493\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18838\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__18838\,
            I => \N__18835\
        );

    \I__2491\ : Span4Mux_h
    port map (
            O => \N__18835\,
            I => \N__18832\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__18832\,
            I => \N__18828\
        );

    \I__2489\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18825\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__18828\,
            I => \POWERLED.count_off_1_4\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__18825\,
            I => \POWERLED.count_off_1_4\
        );

    \I__2486\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18817\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__18817\,
            I => \N__18813\
        );

    \I__2484\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18810\
        );

    \I__2483\ : Span4Mux_s3_v
    port map (
            O => \N__18813\,
            I => \N__18807\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__18810\,
            I => \N__18804\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__18807\,
            I => \N__18801\
        );

    \I__2480\ : Span12Mux_s7_v
    port map (
            O => \N__18804\,
            I => \N__18798\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__18801\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2478\ : Odrv12
    port map (
            O => \N__18798\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2477\ : IoInMux
    port map (
            O => \N__18793\,
            I => \N__18790\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__2475\ : Span4Mux_s3_h
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__18784\,
            I => vccst_en
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \POWERLED.N_359_cascade_\
        );

    \I__2472\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__18775\,
            I => \POWERLED.count_0_2\
        );

    \I__2470\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18769\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__18769\,
            I => \POWERLED.count_0_11\
        );

    \I__2468\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__18763\,
            I => \POWERLED.count_0_3\
        );

    \I__2466\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18757\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__18757\,
            I => \POWERLED.count_0_12\
        );

    \I__2464\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18751\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__18751\,
            I => \N__18748\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__18748\,
            I => \N__18745\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__18745\,
            I => \POWERLED.curr_state_0_0\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__18742\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__18739\,
            I => \curr_state_RNIR5QD1_0_0_cascade_\
        );

    \I__2458\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18733\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__18733\,
            I => \RSMRST_PWRGD.curr_state_2_0\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__18730\,
            I => \RSMRST_PWRGD.m4_0_0_cascade_\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__18727\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__2454\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18721\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__18721\,
            I => \RSMRST_PWRGD.curr_state_7_1\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__18718\,
            I => \N__18714\
        );

    \I__2451\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18695\
        );

    \I__2450\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18695\
        );

    \I__2449\ : InMux
    port map (
            O => \N__18713\,
            I => \N__18695\
        );

    \I__2448\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18695\
        );

    \I__2447\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18683\
        );

    \I__2446\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18683\
        );

    \I__2445\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18683\
        );

    \I__2444\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18683\
        );

    \I__2443\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18683\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__18706\,
            I => \N__18679\
        );

    \I__2441\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18674\
        );

    \I__2440\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18674\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18670\
        );

    \I__2438\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18667\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__18683\,
            I => \N__18664\
        );

    \I__2436\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18659\
        );

    \I__2435\ : InMux
    port map (
            O => \N__18679\,
            I => \N__18659\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18656\
        );

    \I__2433\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18653\
        );

    \I__2432\ : Odrv12
    port map (
            O => \N__18670\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__18667\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__18664\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__18659\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__18656\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__18653\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2426\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__18637\,
            I => \RSMRST_PWRGD.curr_state_1_1\
        );

    \I__2424\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__18631\,
            I => \POWERLED.count_0_10\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__18628\,
            I => \POWERLED.count_0_sqmuxa_i_cascade_\
        );

    \I__2421\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18622\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__18622\,
            I => \POWERLED.count_0_0\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__18619\,
            I => \POWERLED.count_1_0_cascade_\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__18616\,
            I => \POWERLED.countZ0Z_0_cascade_\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__18613\,
            I => \POWERLED.count_1_1_cascade_\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__18610\,
            I => \POWERLED.countZ0Z_1_cascade_\
        );

    \I__2415\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18604\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__18604\,
            I => \POWERLED.count_0_1\
        );

    \I__2413\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18593\
        );

    \I__2412\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18593\
        );

    \I__2411\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18588\
        );

    \I__2410\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18588\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18583\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__18588\,
            I => \N__18583\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__18583\,
            I => \PCH_PWRGD.curr_state_RNI1IPC1Z0Z_0\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__18580\,
            I => \PCH_PWRGD.N_277_0_cascade_\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__18577\,
            I => \N__18573\
        );

    \I__2404\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18570\
        );

    \I__2403\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18567\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__18570\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__18567\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__18562\,
            I => \N__18557\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__18561\,
            I => \N__18554\
        );

    \I__2398\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18550\
        );

    \I__2397\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18545\
        );

    \I__2396\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18545\
        );

    \I__2395\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18542\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18539\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__18545\,
            I => \PCH_PWRGD.N_2857_i\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__18542\,
            I => \PCH_PWRGD.N_2857_i\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__18539\,
            I => \PCH_PWRGD.N_2857_i\
        );

    \I__2390\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18529\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__18529\,
            I => \PCH_PWRGD.N_413\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__18526\,
            I => \PCH_PWRGD.N_413_cascade_\
        );

    \I__2387\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18517\
        );

    \I__2386\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18517\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18513\
        );

    \I__2384\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18510\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__18513\,
            I => \PCH_PWRGD.N_424\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__18510\,
            I => \PCH_PWRGD.N_424\
        );

    \I__2381\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18493\
        );

    \I__2380\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18493\
        );

    \I__2379\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18493\
        );

    \I__2378\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18493\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__18493\,
            I => \N__18490\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__18490\,
            I => \N__18487\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__18487\,
            I => \N__18484\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__18484\,
            I => vr_ready_vccin
        );

    \I__2373\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18472\
        );

    \I__2372\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18472\
        );

    \I__2371\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18472\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__18469\,
            I => \PCH_PWRGD.N_2859_i\
        );

    \I__2368\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__18463\,
            I => \N__18460\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__18460\,
            I => \PCH_PWRGD.N_278_0\
        );

    \I__2365\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18454\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__18454\,
            I => \N__18450\
        );

    \I__2363\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18447\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__18450\,
            I => \N__18444\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__18447\,
            I => \N__18441\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__18444\,
            I => \RSMRST_PWRGD.count_rst_8\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__18441\,
            I => \RSMRST_PWRGD.count_rst_8\
        );

    \I__2358\ : InMux
    port map (
            O => \N__18436\,
            I => \N__18433\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__18430\,
            I => \N__18427\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__18427\,
            I => \RSMRST_PWRGD.count_4_3\
        );

    \I__2354\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18421\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__18421\,
            I => \N__18417\
        );

    \I__2352\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18414\
        );

    \I__2351\ : Span4Mux_h
    port map (
            O => \N__18417\,
            I => \N__18411\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__18414\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__18411\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__18406\,
            I => \N__18403\
        );

    \I__2347\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18400\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__18400\,
            I => \N__18396\
        );

    \I__2345\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18393\
        );

    \I__2344\ : Odrv12
    port map (
            O => \N__18396\,
            I => \PCH_PWRGD.count_rst_11\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__18393\,
            I => \PCH_PWRGD.count_rst_11\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__18388\,
            I => \N__18380\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__18387\,
            I => \N__18374\
        );

    \I__2340\ : CEMux
    port map (
            O => \N__18386\,
            I => \N__18370\
        );

    \I__2339\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18364\
        );

    \I__2338\ : CEMux
    port map (
            O => \N__18384\,
            I => \N__18361\
        );

    \I__2337\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18352\
        );

    \I__2336\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18352\
        );

    \I__2335\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18352\
        );

    \I__2334\ : CEMux
    port map (
            O => \N__18378\,
            I => \N__18352\
        );

    \I__2333\ : CEMux
    port map (
            O => \N__18377\,
            I => \N__18349\
        );

    \I__2332\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18344\
        );

    \I__2331\ : CEMux
    port map (
            O => \N__18373\,
            I => \N__18344\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18340\
        );

    \I__2329\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18337\
        );

    \I__2328\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18326\
        );

    \I__2327\ : CEMux
    port map (
            O => \N__18367\,
            I => \N__18326\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__18364\,
            I => \N__18323\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18320\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18317\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__18349\,
            I => \N__18312\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__18344\,
            I => \N__18309\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__18343\,
            I => \N__18302\
        );

    \I__2320\ : Span4Mux_s3_h
    port map (
            O => \N__18340\,
            I => \N__18295\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__18337\,
            I => \N__18295\
        );

    \I__2318\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18288\
        );

    \I__2317\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18288\
        );

    \I__2316\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18288\
        );

    \I__2315\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18281\
        );

    \I__2314\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18281\
        );

    \I__2313\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18281\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__18326\,
            I => \N__18278\
        );

    \I__2311\ : Span4Mux_s1_v
    port map (
            O => \N__18323\,
            I => \N__18273\
        );

    \I__2310\ : Span4Mux_h
    port map (
            O => \N__18320\,
            I => \N__18273\
        );

    \I__2309\ : Span4Mux_s2_h
    port map (
            O => \N__18317\,
            I => \N__18270\
        );

    \I__2308\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18265\
        );

    \I__2307\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18265\
        );

    \I__2306\ : Span4Mux_s2_h
    port map (
            O => \N__18312\,
            I => \N__18262\
        );

    \I__2305\ : Span4Mux_s2_v
    port map (
            O => \N__18309\,
            I => \N__18259\
        );

    \I__2304\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18252\
        );

    \I__2303\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18252\
        );

    \I__2302\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18252\
        );

    \I__2301\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18249\
        );

    \I__2300\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18242\
        );

    \I__2299\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18242\
        );

    \I__2298\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18242\
        );

    \I__2297\ : Span4Mux_s2_v
    port map (
            O => \N__18295\,
            I => \N__18239\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__18288\,
            I => \N__18234\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__18281\,
            I => \N__18234\
        );

    \I__2294\ : Odrv12
    port map (
            O => \N__18278\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__18273\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__18270\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__18265\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__18262\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__18259\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__18252\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__18249\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__18242\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__18239\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__18234\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\
        );

    \I__2283\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18207\
        );

    \I__2282\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18203\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__18207\,
            I => \N__18200\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__18206\,
            I => \N__18197\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__18203\,
            I => \N__18194\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__18200\,
            I => \N__18191\
        );

    \I__2277\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18188\
        );

    \I__2276\ : Span4Mux_s1_v
    port map (
            O => \N__18194\,
            I => \N__18185\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__18191\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__18188\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__18185\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__18178\,
            I => \VPP_VDDQ.curr_stateZ0Z_0_cascade_\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__18175\,
            I => \N__18172\
        );

    \I__2270\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18169\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__18169\,
            I => \VPP_VDDQ.curr_state_0_1\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__18166\,
            I => \VPP_VDDQ.curr_stateZ0Z_1_cascade_\
        );

    \I__2267\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18160\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__18160\,
            I => \VPP_VDDQ.curr_state_0_0\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__18157\,
            I => \N__18153\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__18156\,
            I => \N__18150\
        );

    \I__2263\ : InMux
    port map (
            O => \N__18153\,
            I => \N__18147\
        );

    \I__2262\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18144\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__18147\,
            I => \N__18141\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18138\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__2258\ : Odrv12
    port map (
            O => \N__18138\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__18135\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2256\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18127\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__18127\,
            I => \PCH_PWRGD.N_277_0\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__18124\,
            I => \PCH_PWRGD.curr_state_7_0_cascade_\
        );

    \I__2253\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18118\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__18118\,
            I => \PCH_PWRGD.curr_state_1_0\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \PCH_PWRGD.N_2857_i_cascade_\
        );

    \I__2249\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18106\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__18106\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__18103\,
            I => \PCH_PWRGD.curr_state_7_1_cascade_\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__18100\,
            I => \N__18096\
        );

    \I__2245\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18085\
        );

    \I__2244\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18085\
        );

    \I__2243\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18085\
        );

    \I__2242\ : InMux
    port map (
            O => \N__18094\,
            I => \N__18085\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__18085\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__18082\,
            I => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__2239\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18075\
        );

    \I__2238\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18072\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__18075\,
            I => \N__18069\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__18072\,
            I => \N__18066\
        );

    \I__2235\ : Span4Mux_s2_v
    port map (
            O => \N__18069\,
            I => \N__18063\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__18066\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__18063\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__2232\ : SRMux
    port map (
            O => \N__18058\,
            I => \N__18054\
        );

    \I__2231\ : SRMux
    port map (
            O => \N__18057\,
            I => \N__18042\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__18054\,
            I => \N__18038\
        );

    \I__2229\ : SRMux
    port map (
            O => \N__18053\,
            I => \N__18035\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__18052\,
            I => \N__18031\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__18051\,
            I => \N__18018\
        );

    \I__2226\ : SRMux
    port map (
            O => \N__18050\,
            I => \N__18014\
        );

    \I__2225\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18006\
        );

    \I__2224\ : InMux
    port map (
            O => \N__18048\,
            I => \N__17997\
        );

    \I__2223\ : InMux
    port map (
            O => \N__18047\,
            I => \N__17997\
        );

    \I__2222\ : InMux
    port map (
            O => \N__18046\,
            I => \N__17997\
        );

    \I__2221\ : InMux
    port map (
            O => \N__18045\,
            I => \N__17997\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__18042\,
            I => \N__17994\
        );

    \I__2219\ : SRMux
    port map (
            O => \N__18041\,
            I => \N__17991\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__18038\,
            I => \N__17986\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__17986\
        );

    \I__2216\ : InMux
    port map (
            O => \N__18034\,
            I => \N__17977\
        );

    \I__2215\ : InMux
    port map (
            O => \N__18031\,
            I => \N__17977\
        );

    \I__2214\ : InMux
    port map (
            O => \N__18030\,
            I => \N__17977\
        );

    \I__2213\ : InMux
    port map (
            O => \N__18029\,
            I => \N__17977\
        );

    \I__2212\ : InMux
    port map (
            O => \N__18028\,
            I => \N__17972\
        );

    \I__2211\ : InMux
    port map (
            O => \N__18027\,
            I => \N__17972\
        );

    \I__2210\ : InMux
    port map (
            O => \N__18026\,
            I => \N__17965\
        );

    \I__2209\ : InMux
    port map (
            O => \N__18025\,
            I => \N__17965\
        );

    \I__2208\ : InMux
    port map (
            O => \N__18024\,
            I => \N__17965\
        );

    \I__2207\ : InMux
    port map (
            O => \N__18023\,
            I => \N__17958\
        );

    \I__2206\ : InMux
    port map (
            O => \N__18022\,
            I => \N__17958\
        );

    \I__2205\ : InMux
    port map (
            O => \N__18021\,
            I => \N__17958\
        );

    \I__2204\ : InMux
    port map (
            O => \N__18018\,
            I => \N__17953\
        );

    \I__2203\ : InMux
    port map (
            O => \N__18017\,
            I => \N__17953\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__18014\,
            I => \N__17950\
        );

    \I__2201\ : InMux
    port map (
            O => \N__18013\,
            I => \N__17947\
        );

    \I__2200\ : InMux
    port map (
            O => \N__18012\,
            I => \N__17942\
        );

    \I__2199\ : InMux
    port map (
            O => \N__18011\,
            I => \N__17942\
        );

    \I__2198\ : InMux
    port map (
            O => \N__18010\,
            I => \N__17939\
        );

    \I__2197\ : SRMux
    port map (
            O => \N__18009\,
            I => \N__17936\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__18006\,
            I => \N__17933\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__17997\,
            I => \N__17930\
        );

    \I__2194\ : Span4Mux_s2_h
    port map (
            O => \N__17994\,
            I => \N__17924\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__17991\,
            I => \N__17924\
        );

    \I__2192\ : Span4Mux_s1_v
    port map (
            O => \N__17986\,
            I => \N__17919\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__17977\,
            I => \N__17919\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__17972\,
            I => \N__17914\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17914\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__17958\,
            I => \N__17909\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__17953\,
            I => \N__17909\
        );

    \I__2186\ : Span4Mux_s3_h
    port map (
            O => \N__17950\,
            I => \N__17906\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__17947\,
            I => \N__17899\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__17942\,
            I => \N__17899\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__17939\,
            I => \N__17899\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__17936\,
            I => \N__17896\
        );

    \I__2181\ : Span4Mux_s3_h
    port map (
            O => \N__17933\,
            I => \N__17891\
        );

    \I__2180\ : Span4Mux_s3_h
    port map (
            O => \N__17930\,
            I => \N__17891\
        );

    \I__2179\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17888\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__17924\,
            I => \N__17879\
        );

    \I__2177\ : Span4Mux_s2_h
    port map (
            O => \N__17919\,
            I => \N__17879\
        );

    \I__2176\ : Span4Mux_v
    port map (
            O => \N__17914\,
            I => \N__17879\
        );

    \I__2175\ : Span4Mux_s1_v
    port map (
            O => \N__17909\,
            I => \N__17879\
        );

    \I__2174\ : IoSpan4Mux
    port map (
            O => \N__17906\,
            I => \N__17874\
        );

    \I__2173\ : Span4Mux_s3_h
    port map (
            O => \N__17899\,
            I => \N__17874\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__17896\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__17891\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__17888\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__17879\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__17874\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__2167\ : InMux
    port map (
            O => \N__17863\,
            I => \N__17859\
        );

    \I__2166\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17854\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__17859\,
            I => \N__17851\
        );

    \I__2164\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17846\
        );

    \I__2163\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17846\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__17854\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__17851\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__17846\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__2159\ : InMux
    port map (
            O => \N__17839\,
            I => \N__17835\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__17838\,
            I => \N__17832\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__17835\,
            I => \N__17829\
        );

    \I__2156\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17826\
        );

    \I__2155\ : Span4Mux_s2_v
    port map (
            O => \N__17829\,
            I => \N__17823\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__17826\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__17823\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__17818\,
            I => \PCH_PWRGD.count_0_sqmuxa_cascade_\
        );

    \I__2151\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17799\
        );

    \I__2150\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17799\
        );

    \I__2149\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17790\
        );

    \I__2148\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17790\
        );

    \I__2147\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17790\
        );

    \I__2146\ : InMux
    port map (
            O => \N__17810\,
            I => \N__17790\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__17809\,
            I => \N__17787\
        );

    \I__2144\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17770\
        );

    \I__2143\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17770\
        );

    \I__2142\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17770\
        );

    \I__2141\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17770\
        );

    \I__2140\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17770\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__17799\,
            I => \N__17763\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__17790\,
            I => \N__17763\
        );

    \I__2137\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17754\
        );

    \I__2136\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17754\
        );

    \I__2135\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17754\
        );

    \I__2134\ : InMux
    port map (
            O => \N__17784\,
            I => \N__17754\
        );

    \I__2133\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17747\
        );

    \I__2132\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17747\
        );

    \I__2131\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17747\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__17770\,
            I => \N__17744\
        );

    \I__2129\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17739\
        );

    \I__2128\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17739\
        );

    \I__2127\ : Span4Mux_s1_v
    port map (
            O => \N__17763\,
            I => \N__17736\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__17754\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__17747\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__17744\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__17739\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__17736\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__17725\,
            I => \N__17722\
        );

    \I__2120\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17719\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__17719\,
            I => \N__17716\
        );

    \I__2118\ : Span4Mux_s1_v
    port map (
            O => \N__17716\,
            I => \N__17713\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__17713\,
            I => \PCH_PWRGD.count_rst_7\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__17710\,
            I => \POWERLED.count_offZ0Z_9_cascade_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17704\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__17704\,
            I => \POWERLED.un34_clk_100khz_11\
        );

    \I__2113\ : InMux
    port map (
            O => \N__17701\,
            I => \N__17697\
        );

    \I__2112\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17694\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__17697\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__17694\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__2109\ : InMux
    port map (
            O => \N__17689\,
            I => \N__17683\
        );

    \I__2108\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17683\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__17683\,
            I => \POWERLED.count_off_1_10\
        );

    \I__2106\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17677\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__17677\,
            I => \POWERLED.count_off_0_10\
        );

    \I__2104\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17670\
        );

    \I__2103\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17667\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__17670\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__17667\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__2100\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17656\
        );

    \I__2099\ : InMux
    port map (
            O => \N__17661\,
            I => \N__17656\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__17656\,
            I => \POWERLED.count_off_1_11\
        );

    \I__2097\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__17650\,
            I => \POWERLED.count_off_0_11\
        );

    \I__2095\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17644\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__17644\,
            I => \POWERLED.count_off_0_12\
        );

    \I__2093\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17637\
        );

    \I__2092\ : InMux
    port map (
            O => \N__17640\,
            I => \N__17634\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__17637\,
            I => \POWERLED.count_off_1_12\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__17634\,
            I => \POWERLED.count_off_1_12\
        );

    \I__2089\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17625\
        );

    \I__2088\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17622\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__17625\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__17622\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__2085\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17613\
        );

    \I__2084\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17610\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__17613\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__17610\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__17605\,
            I => \N__17602\
        );

    \I__2080\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17598\
        );

    \I__2079\ : InMux
    port map (
            O => \N__17601\,
            I => \N__17595\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__17598\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__17595\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__2076\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17586\
        );

    \I__2075\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17583\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__17586\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__17583\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__17578\,
            I => \POWERLED.count_off_1_1_cascade_\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__17575\,
            I => \POWERLED.count_offZ0Z_1_cascade_\
        );

    \I__2070\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17568\
        );

    \I__2069\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17565\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__17568\,
            I => \N__17562\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__17565\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__17562\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__2065\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17554\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__17554\,
            I => \POWERLED.un34_clk_100khz_10\
        );

    \I__2063\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17548\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__17548\,
            I => \POWERLED.un34_clk_100khz_8\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__17545\,
            I => \POWERLED.un34_clk_100khz_9_cascade_\
        );

    \I__2060\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17535\
        );

    \I__2059\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17535\
        );

    \I__2058\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17532\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__17535\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__17532\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2055\ : InMux
    port map (
            O => \N__17527\,
            I => \N__17524\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__17524\,
            I => \POWERLED.count_off_0_1\
        );

    \I__2053\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17501\
        );

    \I__2052\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17492\
        );

    \I__2051\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17492\
        );

    \I__2050\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17492\
        );

    \I__2049\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17492\
        );

    \I__2048\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17483\
        );

    \I__2047\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17483\
        );

    \I__2046\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17483\
        );

    \I__2045\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17483\
        );

    \I__2044\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17476\
        );

    \I__2043\ : InMux
    port map (
            O => \N__17511\,
            I => \N__17476\
        );

    \I__2042\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17476\
        );

    \I__2041\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17469\
        );

    \I__2040\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17469\
        );

    \I__2039\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17469\
        );

    \I__2038\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17462\
        );

    \I__2037\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17462\
        );

    \I__2036\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17462\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__17501\,
            I => \POWERLED.N_128\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__17492\,
            I => \POWERLED.N_128\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__17483\,
            I => \POWERLED.N_128\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__17476\,
            I => \POWERLED.N_128\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__17469\,
            I => \POWERLED.N_128\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__17462\,
            I => \POWERLED.N_128\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__17449\,
            I => \N__17441\
        );

    \I__2028\ : InMux
    port map (
            O => \N__17448\,
            I => \N__17438\
        );

    \I__2027\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17429\
        );

    \I__2026\ : InMux
    port map (
            O => \N__17446\,
            I => \N__17429\
        );

    \I__2025\ : InMux
    port map (
            O => \N__17445\,
            I => \N__17429\
        );

    \I__2024\ : InMux
    port map (
            O => \N__17444\,
            I => \N__17429\
        );

    \I__2023\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17426\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__17438\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__17429\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__17426\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__2019\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17416\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__17416\,
            I => \POWERLED.count_off_0_0\
        );

    \I__2017\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17410\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__17410\,
            I => \POWERLED.count_off_0_9\
        );

    \I__2015\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17401\
        );

    \I__2014\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17401\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__17401\,
            I => \POWERLED.count_off_1_9\
        );

    \I__2012\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__17395\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__17392\,
            I => \POWERLED.count_off_1_0_cascade_\
        );

    \I__2009\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17386\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__17386\,
            I => \POWERLED.func_state_RNI_3Z0Z_0\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__17383\,
            I => \POWERLED.func_state_RNI_3Z0Z_0_cascade_\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__17380\,
            I => \N__17377\
        );

    \I__2005\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17372\
        );

    \I__2004\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17367\
        );

    \I__2003\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17367\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17364\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17361\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__17364\,
            I => \POWERLED.count_clk_RNI_0Z0Z_1\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__17361\,
            I => \POWERLED.count_clk_RNI_0Z0Z_1\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__17356\,
            I => \POWERLED.N_321_cascade_\
        );

    \I__1997\ : InMux
    port map (
            O => \N__17353\,
            I => \N__17348\
        );

    \I__1996\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17345\
        );

    \I__1995\ : InMux
    port map (
            O => \N__17351\,
            I => \N__17342\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__17348\,
            I => \N__17339\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__17345\,
            I => \N__17334\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__17342\,
            I => \N__17334\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__17339\,
            I => \POWERLED.N_431\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__17334\,
            I => \POWERLED.N_431\
        );

    \I__1989\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17326\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__17326\,
            I => \POWERLED.un1_func_state25_6_0_o_N_336_N\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__17323\,
            I => \POWERLED.un1_func_state25_6_0_0_cascade_\
        );

    \I__1986\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17316\
        );

    \I__1985\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17313\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__17316\,
            I => \N__17309\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__17313\,
            I => \N__17306\
        );

    \I__1982\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17303\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__17309\,
            I => \POWERLED.func_state_RNI_1Z0Z_1\
        );

    \I__1980\ : Odrv12
    port map (
            O => \N__17306\,
            I => \POWERLED.func_state_RNI_1Z0Z_1\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__17303\,
            I => \POWERLED.func_state_RNI_1Z0Z_1\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__17296\,
            I => \N__17292\
        );

    \I__1977\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17289\
        );

    \I__1976\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17286\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17283\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__17286\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__17283\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__1972\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17275\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__17275\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__17272\,
            I => \N__17267\
        );

    \I__1969\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17262\
        );

    \I__1968\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17262\
        );

    \I__1967\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17259\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__17262\,
            I => \N__17256\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17253\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__17256\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__17253\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__17248\,
            I => \POWERLED.count_clkZ0Z_2_cascade_\
        );

    \I__1961\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__1960\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17239\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__17239\,
            I => \N__17235\
        );

    \I__1958\ : InMux
    port map (
            O => \N__17238\,
            I => \N__17232\
        );

    \I__1957\ : Odrv12
    port map (
            O => \N__17235\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__17232\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__1955\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17224\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__17224\,
            I => \POWERLED.N_385\
        );

    \I__1953\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17218\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__17218\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__17215\,
            I => \N__17212\
        );

    \I__1950\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__1949\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17203\
        );

    \I__1948\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17198\
        );

    \I__1947\ : InMux
    port map (
            O => \N__17209\,
            I => \N__17198\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__17206\,
            I => \N__17195\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__17203\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__17198\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__17195\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__17188\,
            I => \POWERLED.N_385_cascade_\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__17185\,
            I => \POWERLED.count_clk_en_0_cascade_\
        );

    \I__1940\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17179\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__17179\,
            I => \N__17176\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__17176\,
            I => \POWERLED.un1_func_state25_4_i_a2_1\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__17173\,
            I => \POWERLED.count_clk_en_2_cascade_\
        );

    \I__1936\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17167\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__17167\,
            I => \N__17164\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__17164\,
            I => \N__17160\
        );

    \I__1933\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17157\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__17160\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__17157\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__1930\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17149\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__17149\,
            I => \N__17146\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__17146\,
            I => \POWERLED.count_clk_0_10\
        );

    \I__1927\ : IoInMux
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__17140\,
            I => \N__17137\
        );

    \I__1925\ : Odrv12
    port map (
            O => \N__17137\,
            I => pwrbtn_led
        );

    \I__1924\ : InMux
    port map (
            O => \N__17134\,
            I => \N__17128\
        );

    \I__1923\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17128\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__17125\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__17122\,
            I => \N__17119\
        );

    \I__1919\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__17116\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__17113\,
            I => \POWERLED.count_clkZ0Z_1_cascade_\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__1915\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17104\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__17104\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__17101\,
            I => \N__17098\
        );

    \I__1912\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17093\
        );

    \I__1911\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17088\
        );

    \I__1910\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17088\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__17093\,
            I => \N__17085\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__17088\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__17085\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__1905\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17072\
        );

    \I__1904\ : InMux
    port map (
            O => \N__17076\,
            I => \N__17067\
        );

    \I__1903\ : InMux
    port map (
            O => \N__17075\,
            I => \N__17067\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__17072\,
            I => \N__17064\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__17067\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__17064\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__17059\,
            I => \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__1897\ : InMux
    port map (
            O => \N__17053\,
            I => \N__17047\
        );

    \I__1896\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17047\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__17047\,
            I => \POWERLED.N_193\
        );

    \I__1894\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17041\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__17041\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__1892\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17032\
        );

    \I__1891\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17032\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__17032\,
            I => \N__17029\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__17029\,
            I => \N__17026\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__17026\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__17023\,
            I => \POWERLED.func_state_RNI_1Z0Z_1_cascade_\
        );

    \I__1886\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17017\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__17017\,
            I => \POWERLED.func_state_1_m2_ns_1_1_0\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__17014\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\
        );

    \I__1883\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17008\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__17008\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_1_0\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__17005\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\
        );

    \I__1880\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__1879\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16996\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16993\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__16993\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__16990\,
            I => \N__16987\
        );

    \I__1875\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16984\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__16984\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__1873\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16975\
        );

    \I__1872\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16975\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__16972\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__16969\,
            I => \N__16966\
        );

    \I__1868\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16963\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__16963\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__1866\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16957\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__16957\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__1864\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16951\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__16951\,
            I => \N__16948\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__16948\,
            I => \N__16945\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__16945\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_4\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__16942\,
            I => \POWERLED.count_clkZ0Z_15_cascade_\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__16939\,
            I => \N__16935\
        );

    \I__1858\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16932\
        );

    \I__1857\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16929\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__16932\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__16929\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__1854\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__1853\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16918\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__16918\,
            I => \N__16915\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__16915\,
            I => \POWERLED.N_178\
        );

    \I__1850\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16906\
        );

    \I__1849\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16906\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__16906\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__1847\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16900\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__16900\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__1845\ : InMux
    port map (
            O => \N__16897\,
            I => \N__16891\
        );

    \I__1844\ : InMux
    port map (
            O => \N__16896\,
            I => \N__16891\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__16891\,
            I => \POWERLED.count_clk_1_14\
        );

    \I__1842\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__16885\,
            I => \POWERLED.count_clk_0_14\
        );

    \I__1840\ : InMux
    port map (
            O => \N__16882\,
            I => \N__16876\
        );

    \I__1839\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16876\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__16876\,
            I => \RSMRST_PWRGD.count_rst_4\
        );

    \I__1837\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16870\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__16870\,
            I => \RSMRST_PWRGD.count_4_15\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__16867\,
            I => \RSMRST_PWRGD.N_240_0_cascade_\
        );

    \I__1834\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16861\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16857\
        );

    \I__1832\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16854\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__16857\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__16854\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1829\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16846\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__16846\,
            I => \N__16842\
        );

    \I__1827\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16839\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__16842\,
            I => \RSMRST_PWRGD.count_4_12\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__16839\,
            I => \RSMRST_PWRGD.count_4_12\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__16834\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0_cascade_\
        );

    \I__1823\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16824\
        );

    \I__1822\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16824\
        );

    \I__1821\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16821\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__16824\,
            I => \RSMRST_PWRGD.count_rst_1\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__16821\,
            I => \RSMRST_PWRGD.count_rst_1\
        );

    \I__1818\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16813\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__16813\,
            I => \RSMRST_PWRGD.un12_clk_100khz_4\
        );

    \I__1816\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16804\
        );

    \I__1815\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16804\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__16804\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__1813\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16798\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__16798\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__16795\,
            I => \N__16792\
        );

    \I__1810\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16788\
        );

    \I__1809\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16785\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__16788\,
            I => \N__16782\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__16785\,
            I => \N__16779\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__16782\,
            I => \RSMRST_PWRGD.un2_count_1_axb_9\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__16779\,
            I => \RSMRST_PWRGD.un2_count_1_axb_9\
        );

    \I__1804\ : InMux
    port map (
            O => \N__16774\,
            I => \N__16768\
        );

    \I__1803\ : InMux
    port map (
            O => \N__16773\,
            I => \N__16768\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__16768\,
            I => \N__16765\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__16765\,
            I => \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1800\ : InMux
    port map (
            O => \N__16762\,
            I => \bfn_2_7_0_\
        );

    \I__1799\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16754\
        );

    \I__1798\ : InMux
    port map (
            O => \N__16758\,
            I => \N__16749\
        );

    \I__1797\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16749\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__16754\,
            I => \N__16746\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__16749\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__16746\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__16741\,
            I => \N__16737\
        );

    \I__1792\ : InMux
    port map (
            O => \N__16740\,
            I => \N__16732\
        );

    \I__1791\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16732\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__16732\,
            I => \N__16729\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__16729\,
            I => \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO\
        );

    \I__1788\ : InMux
    port map (
            O => \N__16726\,
            I => \RSMRST_PWRGD.un2_count_1_cry_9\
        );

    \I__1787\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16719\
        );

    \I__1786\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16716\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__16719\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__16716\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1783\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16705\
        );

    \I__1782\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16705\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__16705\,
            I => \RSMRST_PWRGD.count_rst_0\
        );

    \I__1780\ : InMux
    port map (
            O => \N__16702\,
            I => \RSMRST_PWRGD.un2_count_1_cry_10\
        );

    \I__1779\ : InMux
    port map (
            O => \N__16699\,
            I => \RSMRST_PWRGD.un2_count_1_cry_11\
        );

    \I__1778\ : InMux
    port map (
            O => \N__16696\,
            I => \N__16691\
        );

    \I__1777\ : InMux
    port map (
            O => \N__16695\,
            I => \N__16688\
        );

    \I__1776\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16685\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__16691\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__16688\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__16685\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1772\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16675\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__16675\,
            I => \N__16671\
        );

    \I__1770\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16668\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__16671\,
            I => \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__16668\,
            I => \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\
        );

    \I__1767\ : InMux
    port map (
            O => \N__16663\,
            I => \RSMRST_PWRGD.un2_count_1_cry_12\
        );

    \I__1766\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16657\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__16657\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1764\ : InMux
    port map (
            O => \N__16654\,
            I => \N__16648\
        );

    \I__1763\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16648\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__16648\,
            I => \RSMRST_PWRGD.count_rst_3\
        );

    \I__1761\ : InMux
    port map (
            O => \N__16645\,
            I => \RSMRST_PWRGD.un2_count_1_cry_13\
        );

    \I__1760\ : InMux
    port map (
            O => \N__16642\,
            I => \RSMRST_PWRGD.un2_count_1_cry_14\
        );

    \I__1759\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16636\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__16636\,
            I => \RSMRST_PWRGD.un2_count_1_axb_12\
        );

    \I__1757\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16626\
        );

    \I__1756\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16626\
        );

    \I__1755\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16623\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__16626\,
            I => \RSMRST_PWRGD.un2_count_1_axb_1\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__16623\,
            I => \RSMRST_PWRGD.un2_count_1_axb_1\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__16618\,
            I => \N__16615\
        );

    \I__1751\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16608\
        );

    \I__1750\ : InMux
    port map (
            O => \N__16614\,
            I => \N__16599\
        );

    \I__1749\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16599\
        );

    \I__1748\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16599\
        );

    \I__1747\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16599\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__16608\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__16599\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1744\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16591\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__16591\,
            I => \RSMRST_PWRGD.un2_count_1_axb_2\
        );

    \I__1742\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16579\
        );

    \I__1741\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16579\
        );

    \I__1740\ : InMux
    port map (
            O => \N__16586\,
            I => \N__16579\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__16579\,
            I => \RSMRST_PWRGD.count_rst_7\
        );

    \I__1738\ : InMux
    port map (
            O => \N__16576\,
            I => \RSMRST_PWRGD.un2_count_1_cry_1\
        );

    \I__1737\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16569\
        );

    \I__1736\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16566\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16563\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16560\
        );

    \I__1733\ : Odrv12
    port map (
            O => \N__16563\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__16560\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1731\ : InMux
    port map (
            O => \N__16555\,
            I => \RSMRST_PWRGD.un2_count_1_cry_2\
        );

    \I__1730\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16545\
        );

    \I__1729\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16545\
        );

    \I__1728\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16542\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__16545\,
            I => \RSMRST_PWRGD.un2_count_1_axb_4\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__16542\,
            I => \RSMRST_PWRGD.un2_count_1_axb_4\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__16537\,
            I => \N__16534\
        );

    \I__1724\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16528\
        );

    \I__1723\ : InMux
    port map (
            O => \N__16533\,
            I => \N__16528\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__16528\,
            I => \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1721\ : InMux
    port map (
            O => \N__16525\,
            I => \RSMRST_PWRGD.un2_count_1_cry_3\
        );

    \I__1720\ : InMux
    port map (
            O => \N__16522\,
            I => \N__16519\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__16516\,
            I => \RSMRST_PWRGD.un2_count_1_axb_5\
        );

    \I__1717\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16504\
        );

    \I__1716\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16504\
        );

    \I__1715\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16504\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__16504\,
            I => \N__16501\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__16501\,
            I => \RSMRST_PWRGD.count_rst_10\
        );

    \I__1712\ : InMux
    port map (
            O => \N__16498\,
            I => \RSMRST_PWRGD.un2_count_1_cry_4\
        );

    \I__1711\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16491\
        );

    \I__1710\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16488\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__16491\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__16488\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1707\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16477\
        );

    \I__1706\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16477\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__16477\,
            I => \RSMRST_PWRGD.count_rst_11\
        );

    \I__1704\ : InMux
    port map (
            O => \N__16474\,
            I => \RSMRST_PWRGD.un2_count_1_cry_5\
        );

    \I__1703\ : InMux
    port map (
            O => \N__16471\,
            I => \RSMRST_PWRGD.un2_count_1_cry_6\
        );

    \I__1702\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16463\
        );

    \I__1701\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16460\
        );

    \I__1700\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16457\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__16463\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__16460\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__16457\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1696\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16444\
        );

    \I__1695\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16444\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__16444\,
            I => \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1693\ : InMux
    port map (
            O => \N__16441\,
            I => \RSMRST_PWRGD.un2_count_1_cry_7\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__16438\,
            I => \N__16434\
        );

    \I__1691\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16431\
        );

    \I__1690\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16427\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__16431\,
            I => \N__16424\
        );

    \I__1688\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16421\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__16427\,
            I => \PCH_PWRGD.count_i_0\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__16424\,
            I => \PCH_PWRGD.count_i_0\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__16421\,
            I => \PCH_PWRGD.count_i_0\
        );

    \I__1684\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16410\
        );

    \I__1683\ : InMux
    port map (
            O => \N__16413\,
            I => \N__16407\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__16410\,
            I => \N__16404\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__16407\,
            I => \N__16401\
        );

    \I__1680\ : Span4Mux_s0_v
    port map (
            O => \N__16404\,
            I => \N__16396\
        );

    \I__1679\ : Span4Mux_s1_h
    port map (
            O => \N__16401\,
            I => \N__16396\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__16396\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__16393\,
            I => \RSMRST_PWRGD.count_rst_14_cascade_\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__16390\,
            I => \RSMRST_PWRGD.un2_count_1_axb_9_cascade_\
        );

    \I__1675\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16384\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__16384\,
            I => \RSMRST_PWRGD.count_rst_14\
        );

    \I__1673\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16375\
        );

    \I__1672\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16375\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__16375\,
            I => \RSMRST_PWRGD.count_4_9\
        );

    \I__1670\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16369\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__16369\,
            I => \N__16366\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__16366\,
            I => \RSMRST_PWRGD.un12_clk_100khz_1\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__16363\,
            I => \RSMRST_PWRGD.count_rst_cascade_\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__16360\,
            I => \RSMRST_PWRGD.countZ0Z_10_cascade_\
        );

    \I__1665\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16354\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__16354\,
            I => \RSMRST_PWRGD.count_4_10\
        );

    \I__1663\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16348\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__16348\,
            I => \RSMRST_PWRGD.count_4_13\
        );

    \I__1661\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16339\
        );

    \I__1660\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16339\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__16339\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__16336\,
            I => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0_cascade_\
        );

    \I__1657\ : InMux
    port map (
            O => \N__16333\,
            I => \N__16330\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__16330\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__1655\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16323\
        );

    \I__1654\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16320\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__16323\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__16320\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__16315\,
            I => \PCH_PWRGD.un2_count_1_axb_8_cascade_\
        );

    \I__1650\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16309\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__16309\,
            I => \PCH_PWRGD.count_rst_6\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__16306\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1647\ : InMux
    port map (
            O => \N__16303\,
            I => \N__16300\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__16300\,
            I => \N__16297\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__16297\,
            I => \PCH_PWRGD.un12_clk_100khz_6\
        );

    \I__1644\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16290\
        );

    \I__1643\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16287\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__16290\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__16287\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__16282\,
            I => \N__16279\
        );

    \I__1639\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16273\
        );

    \I__1638\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16273\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__16273\,
            I => \N__16270\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__16270\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1635\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16261\
        );

    \I__1634\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16261\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__16261\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__16258\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__1631\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16250\
        );

    \I__1630\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16245\
        );

    \I__1629\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16245\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__16250\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__16245\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__16240\,
            I => \N__16237\
        );

    \I__1625\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16233\
        );

    \I__1624\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16230\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__16233\,
            I => \N__16227\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__16230\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__16227\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__16222\,
            I => \PCH_PWRGD.countZ0Z_9_cascade_\
        );

    \I__1619\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__16216\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__1617\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__16210\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__1615\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__16204\,
            I => \PCH_PWRGD.count_rst_9\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__16201\,
            I => \N__16197\
        );

    \I__1612\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16194\
        );

    \I__1611\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__16194\,
            I => \PCH_PWRGD.un2_count_1_axb_5\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__16191\,
            I => \PCH_PWRGD.un2_count_1_axb_5\
        );

    \I__1608\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16180\
        );

    \I__1607\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16180\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__16180\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__16177\,
            I => \PCH_PWRGD.un2_count_1_axb_5_cascade_\
        );

    \I__1604\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16168\
        );

    \I__1603\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16168\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__16168\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__1601\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16162\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__16162\,
            I => \N__16159\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__16159\,
            I => \PCH_PWRGD.un12_clk_100khz_1\
        );

    \I__1598\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16153\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__16153\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__1596\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16141\
        );

    \I__1595\ : InMux
    port map (
            O => \N__16149\,
            I => \N__16141\
        );

    \I__1594\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16141\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__16141\,
            I => \N__16138\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__16138\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1591\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16129\
        );

    \I__1590\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16129\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__16129\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__1588\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16120\
        );

    \I__1587\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16120\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__16120\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__1585\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16114\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__16114\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__1583\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16107\
        );

    \I__1582\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16104\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__16107\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__16104\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1579\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16096\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__16096\,
            I => \PCH_PWRGD.count_rst_14\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__16093\,
            I => \PCH_PWRGD.count_rst_14_cascade_\
        );

    \I__1576\ : InMux
    port map (
            O => \N__16090\,
            I => \N__16087\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__16087\,
            I => \N__16084\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__16084\,
            I => \PCH_PWRGD.un2_count_1_axb_0\
        );

    \I__1573\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16075\
        );

    \I__1572\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16075\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__16075\,
            I => \N__16072\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__16072\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__1569\ : InMux
    port map (
            O => \N__16069\,
            I => \N__16066\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__16066\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__16063\,
            I => \PCH_PWRGD.count_rst_9_cascade_\
        );

    \I__1566\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__16057\,
            I => \PCH_PWRGD.un12_clk_100khz_7\
        );

    \I__1564\ : InMux
    port map (
            O => \N__16054\,
            I => \N__16051\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__16051\,
            I => \N__16048\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__16048\,
            I => \PCH_PWRGD.un12_clk_100khz_4\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__16045\,
            I => \PCH_PWRGD.un12_clk_100khz_5_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16039\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__16039\,
            I => \PCH_PWRGD.un12_clk_100khz_0\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__16036\,
            I => \PCH_PWRGD.un12_clk_100khz_13_cascade_\
        );

    \I__1557\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16030\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__16030\,
            I => \PCH_PWRGD.un12_clk_100khz_9\
        );

    \I__1555\ : InMux
    port map (
            O => \N__16027\,
            I => \N__16021\
        );

    \I__1554\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16021\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__16021\,
            I => \N__16018\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__16018\,
            I => \POWERLED.count_off_1_5\
        );

    \I__1551\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16012\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__16012\,
            I => \POWERLED.count_off_0_5\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__16009\,
            I => \N__16006\
        );

    \I__1548\ : InMux
    port map (
            O => \N__16006\,
            I => \N__16000\
        );

    \I__1547\ : InMux
    port map (
            O => \N__16005\,
            I => \N__16000\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__16000\,
            I => \POWERLED.count_off_1_14\
        );

    \I__1545\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15994\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__15994\,
            I => \POWERLED.count_off_0_14\
        );

    \I__1543\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15985\
        );

    \I__1542\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15985\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__15985\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNINZ0Z4153\
        );

    \I__1540\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15979\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__15979\,
            I => \POWERLED.count_off_0_15\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__15976\,
            I => \N__15973\
        );

    \I__1537\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15967\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__15967\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__15964\,
            I => \N__15961\
        );

    \I__1533\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15952\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15952\
        );

    \I__1531\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15952\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__15952\,
            I => \N__15949\
        );

    \I__1529\ : Span4Mux_s1_v
    port map (
            O => \N__15949\,
            I => \N__15946\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__15946\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1527\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15937\
        );

    \I__1526\ : InMux
    port map (
            O => \N__15942\,
            I => \N__15937\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__15937\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__15934\,
            I => \N__15931\
        );

    \I__1523\ : InMux
    port map (
            O => \N__15931\,
            I => \N__15927\
        );

    \I__1522\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15924\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__15927\,
            I => \N__15921\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__15924\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__15921\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1518\ : InMux
    port map (
            O => \N__15916\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__1517\ : InMux
    port map (
            O => \N__15913\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__1516\ : InMux
    port map (
            O => \N__15910\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__1515\ : InMux
    port map (
            O => \N__15907\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__1514\ : InMux
    port map (
            O => \N__15904\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__1513\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15895\
        );

    \I__1512\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15895\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__15895\,
            I => \POWERLED.count_off_1_13\
        );

    \I__1510\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15889\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__15889\,
            I => \POWERLED.count_off_0_13\
        );

    \I__1508\ : InMux
    port map (
            O => \N__15886\,
            I => \POWERLED.un3_count_off_1_cry_1\
        );

    \I__1507\ : InMux
    port map (
            O => \N__15883\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__1506\ : InMux
    port map (
            O => \N__15880\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__1505\ : InMux
    port map (
            O => \N__15877\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__1504\ : InMux
    port map (
            O => \N__15874\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__1503\ : InMux
    port map (
            O => \N__15871\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__1502\ : InMux
    port map (
            O => \N__15868\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__1501\ : InMux
    port map (
            O => \N__15865\,
            I => \bfn_1_15_0_\
        );

    \I__1500\ : InMux
    port map (
            O => \N__15862\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__15859\,
            I => \POWERLED.count_clkZ0Z_13_cascade_\
        );

    \I__1498\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15852\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15849\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__15852\,
            I => \N__15846\
        );

    \I__1495\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15843\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__15846\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__15843\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__15838\,
            I => \N__15835\
        );

    \I__1491\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15831\
        );

    \I__1490\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__15831\,
            I => \N__15825\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__15828\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__15825\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__1486\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15814\
        );

    \I__1485\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15814\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__15814\,
            I => \N__15811\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__15811\,
            I => \POWERLED.count_clk_1_13\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__15808\,
            I => \N__15805\
        );

    \I__1481\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15802\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__15802\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__15799\,
            I => \N__15796\
        );

    \I__1478\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15793\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__15793\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__1476\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15784\
        );

    \I__1475\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15784\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__15784\,
            I => \N__15781\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__15781\,
            I => \POWERLED.count_clk_1_11\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__15778\,
            I => \N__15775\
        );

    \I__1471\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15771\
        );

    \I__1470\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15768\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__15771\,
            I => \N__15765\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__15768\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__15765\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__1466\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15754\
        );

    \I__1465\ : InMux
    port map (
            O => \N__15759\,
            I => \N__15754\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15751\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__15751\,
            I => \POWERLED.count_clk_1_12\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__15748\,
            I => \N__15745\
        );

    \I__1461\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15742\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__15742\,
            I => \POWERLED.count_clk_0_12\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__15739\,
            I => \POWERLED.count_clkZ0Z_5_cascade_\
        );

    \I__1458\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15730\
        );

    \I__1457\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15730\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15727\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__15727\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__15724\,
            I => \N__15721\
        );

    \I__1453\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15718\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__15718\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15711\
        );

    \I__1450\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15708\
        );

    \I__1449\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15705\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__15708\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__15705\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__15700\,
            I => \N__15697\
        );

    \I__1445\ : InMux
    port map (
            O => \N__15697\,
            I => \N__15693\
        );

    \I__1444\ : InMux
    port map (
            O => \N__15696\,
            I => \N__15690\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__15693\,
            I => \N__15687\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__15690\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__15687\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__15682\,
            I => \POWERLED.count_clkZ0Z_9_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__1438\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15673\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__15673\,
            I => \N__15670\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__15670\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__15667\,
            I => \N__15664\
        );

    \I__1434\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15661\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__15661\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__1432\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15652\
        );

    \I__1431\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15652\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__15652\,
            I => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \N__15646\
        );

    \I__1428\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15643\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__15643\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__15640\,
            I => \N__15637\
        );

    \I__1425\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15634\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15631\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__15631\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__1422\ : InMux
    port map (
            O => \N__15628\,
            I => \bfn_1_10_0_\
        );

    \I__1421\ : InMux
    port map (
            O => \N__15625\,
            I => \POWERLED.un1_count_clk_2_cry_9\
        );

    \I__1420\ : InMux
    port map (
            O => \N__15622\,
            I => \POWERLED.un1_count_clk_2_cry_10_cZ0\
        );

    \I__1419\ : InMux
    port map (
            O => \N__15619\,
            I => \POWERLED.un1_count_clk_2_cry_11\
        );

    \I__1418\ : InMux
    port map (
            O => \N__15616\,
            I => \POWERLED.un1_count_clk_2_cry_12\
        );

    \I__1417\ : InMux
    port map (
            O => \N__15613\,
            I => \POWERLED.un1_count_clk_2_cry_13\
        );

    \I__1416\ : InMux
    port map (
            O => \N__15610\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__1415\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15604\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__15604\,
            I => \RSMRST_PWRGD.count_4_11\
        );

    \I__1413\ : InMux
    port map (
            O => \N__15601\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__1412\ : InMux
    port map (
            O => \N__15598\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__1411\ : InMux
    port map (
            O => \N__15595\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__1410\ : InMux
    port map (
            O => \N__15592\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__1409\ : InMux
    port map (
            O => \N__15589\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__1408\ : InMux
    port map (
            O => \N__15586\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15583\,
            I => \POWERLED.un1_count_clk_2_cry_7_cZ0\
        );

    \I__1406\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15577\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__15577\,
            I => \N__15574\
        );

    \I__1404\ : Odrv4
    port map (
            O => \N__15574\,
            I => \RSMRST_PWRGD.un12_clk_100khz_12\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__15571\,
            I => \RSMRST_PWRGD.un12_clk_100khz_11_cascade_\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__15568\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12_cascade_\
        );

    \I__1401\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15562\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__15562\,
            I => \RSMRST_PWRGD.count_4_0\
        );

    \I__1399\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15556\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__15556\,
            I => \RSMRST_PWRGD.count_4_14\
        );

    \I__1397\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15549\
        );

    \I__1396\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15546\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__15549\,
            I => \RSMRST_PWRGD.count_4_5\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__15546\,
            I => \RSMRST_PWRGD.count_4_5\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__15541\,
            I => \RSMRST_PWRGD.countZ0Z_14_cascade_\
        );

    \I__1392\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15535\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__15535\,
            I => \RSMRST_PWRGD.un12_clk_100khz_5\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__15532\,
            I => \RSMRST_PWRGD.countZ0Z_13_cascade_\
        );

    \I__1389\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15526\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__15526\,
            I => \RSMRST_PWRGD.un12_clk_100khz_2\
        );

    \I__1387\ : InMux
    port map (
            O => \N__15523\,
            I => \N__15520\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__15520\,
            I => \RSMRST_PWRGD.count_rst_13\
        );

    \I__1385\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15514\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__15514\,
            I => \RSMRST_PWRGD.count_4_6\
        );

    \I__1383\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15508\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__15508\,
            I => \RSMRST_PWRGD.count_rst_6\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__15505\,
            I => \RSMRST_PWRGD.count_rst_6_cascade_\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__15502\,
            I => \RSMRST_PWRGD.count_rst_5_cascade_\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__15499\,
            I => \RSMRST_PWRGD.countZ0Z_0_cascade_\
        );

    \I__1378\ : InMux
    port map (
            O => \N__15496\,
            I => \N__15492\
        );

    \I__1377\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15489\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__15492\,
            I => \RSMRST_PWRGD.count_4_1\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__15489\,
            I => \RSMRST_PWRGD.count_4_1\
        );

    \I__1374\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15481\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__15481\,
            I => \RSMRST_PWRGD.count_rst_9\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__15478\,
            I => \RSMRST_PWRGD.count_rst_9_cascade_\
        );

    \I__1371\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15472\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__15472\,
            I => \RSMRST_PWRGD.un12_clk_100khz_3\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__15469\,
            I => \RSMRST_PWRGD.un12_clk_100khz_0_cascade_\
        );

    \I__1368\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15460\
        );

    \I__1367\ : InMux
    port map (
            O => \N__15465\,
            I => \N__15460\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__15460\,
            I => \RSMRST_PWRGD.count_4_4\
        );

    \I__1365\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15451\
        );

    \I__1364\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15451\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__15451\,
            I => \RSMRST_PWRGD.count_4_2\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__15448\,
            I => \RSMRST_PWRGD.countZ0Z_8_cascade_\
        );

    \I__1361\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15442\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__15442\,
            I => \RSMRST_PWRGD.count_4_8\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__15439\,
            I => \RSMRST_PWRGD.count_rst_2_cascade_\
        );

    \I__1358\ : InMux
    port map (
            O => \N__15436\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__1357\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15430\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__15430\,
            I => \N__15427\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__15427\,
            I => \N__15422\
        );

    \I__1354\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15417\
        );

    \I__1353\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15417\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__15422\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__15417\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__1350\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15406\
        );

    \I__1349\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15406\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__15406\,
            I => \N__15403\
        );

    \I__1347\ : Span4Mux_s2_v
    port map (
            O => \N__15403\,
            I => \N__15400\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__15400\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1345\ : InMux
    port map (
            O => \N__15397\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__1344\ : InMux
    port map (
            O => \N__15394\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__1343\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15387\
        );

    \I__1342\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15384\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__15387\,
            I => \N__15381\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__15384\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__15381\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1338\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15370\
        );

    \I__1337\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15370\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__15370\,
            I => \N__15367\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__15367\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__1334\ : InMux
    port map (
            O => \N__15364\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__1333\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15357\
        );

    \I__1332\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15354\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__15357\,
            I => \N__15351\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__15354\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__15351\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1328\ : InMux
    port map (
            O => \N__15346\,
            I => \N__15340\
        );

    \I__1327\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15340\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15337\
        );

    \I__1325\ : Odrv12
    port map (
            O => \N__15337\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__1324\ : InMux
    port map (
            O => \N__15334\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__1323\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15328\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__15328\,
            I => \N__15324\
        );

    \I__1321\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15321\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__15324\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__15321\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1318\ : InMux
    port map (
            O => \N__15316\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__1317\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15307\
        );

    \I__1316\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15307\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__15307\,
            I => \N__15304\
        );

    \I__1314\ : Odrv12
    port map (
            O => \N__15304\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__1313\ : InMux
    port map (
            O => \N__15301\,
            I => \PCH_PWRGD.un2_count_1_cry_0\
        );

    \I__1312\ : InMux
    port map (
            O => \N__15298\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__1311\ : InMux
    port map (
            O => \N__15295\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__1310\ : InMux
    port map (
            O => \N__15292\,
            I => \N__15289\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15284\
        );

    \I__1308\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15279\
        );

    \I__1307\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15279\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__15284\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__15279\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__15274\,
            I => \N__15270\
        );

    \I__1303\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15265\
        );

    \I__1302\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15265\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__15265\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1300\ : InMux
    port map (
            O => \N__15262\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__1299\ : InMux
    port map (
            O => \N__15259\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__1298\ : InMux
    port map (
            O => \N__15256\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__1297\ : InMux
    port map (
            O => \N__15253\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__1296\ : InMux
    port map (
            O => \N__15250\,
            I => \bfn_1_4_0_\
        );

    \I__1295\ : InMux
    port map (
            O => \N__15247\,
            I => \PCH_PWRGD.un2_count_1_cry_8\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__15244\,
            I => \PCH_PWRGD.count_rst_3_cascade_\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__15241\,
            I => \PCH_PWRGD.countZ0Z_4_cascade_\
        );

    \I__1292\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15235\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__15235\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__1290\ : InMux
    port map (
            O => \N__15232\,
            I => \N__15229\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__15229\,
            I => \PCH_PWRGD.count_rst_3\
        );

    \I__1288\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15223\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__15223\,
            I => \PCH_PWRGD.count_rst_10\
        );

    \I__1286\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__1285\ : InMux
    port map (
            O => \N__15219\,
            I => \N__15214\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__15214\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__1283\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15208\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__15208\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__1281\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15202\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__15202\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__1279\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15196\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__15196\,
            I => \PCH_PWRGD.count_0_14\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un4_count_1_cry_7_cZ0\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un2_count_1_cry_8\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un2_count_1_cry_16\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.un4_counter_7\,
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_6_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_6_16_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_7_6_0_\
        );

    \HDA_STRAP.count_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22045\,
            GLOBALBUFFEROUTPUT => \HDA_STRAP.count_en_g\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29965\,
            GLOBALBUFFEROUTPUT => \VPP_VDDQ_delayed_vddq_pwrgd_en_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIGIDI3_0_0_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15390\,
            in1 => \N__15360\,
            in2 => \N__16438\,
            in3 => \N__15327\,
            lcout => \PCH_PWRGD.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI2FVK5_15_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18385\,
            in1 => \N__15211\,
            in2 => \_gnd_net_\,
            in3 => \N__15312\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15313\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35092\,
            ce => \N__18377\,
            sr => \N__18050\
        );

    \PCH_PWRGD.count_RNIU8TK5_13_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15376\,
            in1 => \N__15205\,
            in2 => \_gnd_net_\,
            in3 => \N__18333\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15375\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35092\,
            ce => \N__18377\,
            sr => \N__18050\
        );

    \PCH_PWRGD.count_RNI0CUK5_14_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15346\,
            in1 => \N__15199\,
            in2 => \_gnd_net_\,
            in3 => \N__18332\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_14_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15345\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35092\,
            ce => \N__18377\,
            sr => \N__18050\
        );

    \PCH_PWRGD.count_RNIGIDI3_0_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__16099\,
            in1 => \N__16413\,
            in2 => \_gnd_net_\,
            in3 => \N__18331\,
            lcout => \PCH_PWRGD.count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNIORTP1_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__18034\,
            in1 => \N__15412\,
            in2 => \N__17809\,
            in3 => \N__15426\,
            lcout => \PCH_PWRGD.count_rst_3\,
            ltout => \PCH_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQ2RK5_11_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18379\,
            in2 => \N__15244\,
            in3 => \N__15219\,
            lcout => \PCH_PWRGD.un2_count_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIUUIH5_4_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15238\,
            in1 => \N__15226\,
            in2 => \_gnd_net_\,
            in3 => \N__18305\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => \PCH_PWRGD.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__15273\,
            in1 => \N__18030\,
            in2 => \N__15241\,
            in3 => \N__17786\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35259\,
            ce => \N__18378\,
            sr => \N__18009\
        );

    \PCH_PWRGD.count_RNIQ2RK5_0_11_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__15220\,
            in1 => \N__15232\,
            in2 => \N__18388\,
            in3 => \N__16327\,
            lcout => \PCH_PWRGD.un12_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNIA85V1_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__15287\,
            in1 => \N__18029\,
            in2 => \N__15274\,
            in3 => \N__17784\,
            lcout => \PCH_PWRGD.count_rst_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_11_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__17785\,
            in1 => \N__15411\,
            in2 => \N__18052\,
            in3 => \N__15425\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35259\,
            ce => \N__18378\,
            sr => \N__18009\
        );

    \PCH_PWRGD.count_RNISRHH5_0_3_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15288\,
            in1 => \N__18420\,
            in2 => \N__18406\,
            in3 => \N__18383\,
            lcout => \PCH_PWRGD.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_0_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16090\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_0_c_RNI722V1_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18013\,
            in1 => \N__16326\,
            in2 => \_gnd_net_\,
            in3 => \N__15301\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_0\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNI843V1_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__18011\,
            in1 => \_gnd_net_\,
            in2 => \N__15976\,
            in3 => \N__15298\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18211\,
            in2 => \_gnd_net_\,
            in3 => \N__15295\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15292\,
            in2 => \_gnd_net_\,
            in3 => \N__15262\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16200\,
            in2 => \_gnd_net_\,
            in3 => \N__15259\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNICC7V1_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__18012\,
            in1 => \_gnd_net_\,
            in2 => \N__15934\,
            in3 => \N__15256\,
            lcout => \PCH_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17862\,
            in2 => \_gnd_net_\,
            in3 => \N__15253\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16294\,
            in2 => \_gnd_net_\,
            in3 => \N__15250\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16255\,
            in2 => \_gnd_net_\,
            in3 => \N__15247\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIGKBV1_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18046\,
            in1 => \N__16156\,
            in2 => \_gnd_net_\,
            in3 => \N__15436\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15433\,
            in2 => \_gnd_net_\,
            in3 => \N__15397\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNIPTUP1_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18047\,
            in1 => \N__16110\,
            in2 => \_gnd_net_\,
            in3 => \N__15394\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIQVVP1_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18049\,
            in1 => \N__15391\,
            in2 => \_gnd_net_\,
            in3 => \N__15364\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIR11Q1_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18045\,
            in1 => \N__15361\,
            in2 => \_gnd_net_\,
            in3 => \N__15334\,
            lcout => \PCH_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNIS32Q1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__15331\,
            in1 => \N__18048\,
            in2 => \_gnd_net_\,
            in3 => \N__15316\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010011"
        )
    port map (
            in0 => \N__16587\,
            in1 => \N__15457\,
            in2 => \N__28959\,
            in3 => \N__16573\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI8NK06_2_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15456\,
            in1 => \N__28923\,
            in2 => \_gnd_net_\,
            in3 => \N__16586\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNICTM06_4_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28924\,
            in1 => \N__15465\,
            in2 => \_gnd_net_\,
            in3 => \N__15484\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__16551\,
            in1 => \N__16533\,
            in2 => \N__19981\,
            in3 => \N__18704\,
            lcout => \RSMRST_PWRGD.count_rst_9\,
            ltout => \RSMRST_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNICTM06_0_4_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__28928\,
            in1 => \N__15466\,
            in2 => \N__15478\,
            in3 => \N__16467\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un12_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI91BKN_1_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15475\,
            in1 => \N__16372\,
            in2 => \N__15469\,
            in3 => \N__15529\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_4_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__18705\,
            in1 => \N__16552\,
            in2 => \N__16537\,
            in3 => \N__19972\,
            lcout => \RSMRST_PWRGD.count_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35199\,
            ce => \N__28975\,
            sr => \N__19979\
        );

    \RSMRST_PWRGD.count_2_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16588\,
            lcout => \RSMRST_PWRGD.count_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35199\,
            ce => \N__28975\,
            sr => \N__19979\
        );

    \RSMRST_PWRGD.count_RNIK9R06_8_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15445\,
            in1 => \N__28930\,
            in2 => \_gnd_net_\,
            in3 => \N__15523\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => \RSMRST_PWRGD.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_8_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__18682\,
            in1 => \N__16450\,
            in2 => \N__15448\,
            in3 => \N__19944\,
            lcout => \RSMRST_PWRGD.count_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35235\,
            ce => \N__28941\,
            sr => \N__19973\
        );

    \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__18694\,
            in1 => \N__16696\,
            in2 => \N__19976\,
            in3 => \N__16674\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.count_rst_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIC74M5_13_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__28931\,
            in1 => \_gnd_net_\,
            in2 => \N__15439\,
            in3 => \N__16351\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => \RSMRST_PWRGD.countZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__15511\,
            in1 => \N__28932\,
            in2 => \N__15532\,
            in3 => \N__15496\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__16468\,
            in1 => \N__16449\,
            in2 => \N__18706\,
            in3 => \N__19940\,
            lcout => \RSMRST_PWRGD.count_rst_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIG3P06_6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16482\,
            in1 => \N__28929\,
            in2 => \_gnd_net_\,
            in3 => \N__15517\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_6_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16483\,
            lcout => \RSMRST_PWRGD.count_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35235\,
            ce => \N__28941\,
            sr => \N__19973\
        );

    \RSMRST_PWRGD.count_RNIAB7J1_1_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19966\,
            in1 => \N__16611\,
            in2 => \_gnd_net_\,
            in3 => \N__16632\,
            lcout => \RSMRST_PWRGD.count_rst_6\,
            ltout => \RSMRST_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIVV2I5_1_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15495\,
            in2 => \N__15505\,
            in3 => \N__28865\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIAB7J1_0_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19965\,
            in1 => \N__18673\,
            in2 => \_gnd_net_\,
            in3 => \N__16614\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIUU2I5_0_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15565\,
            in2 => \N__15502\,
            in3 => \N__28864\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => \RSMRST_PWRGD.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_1_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19967\,
            in1 => \_gnd_net_\,
            in2 => \N__15499\,
            in3 => \N__16633\,
            lcout => \RSMRST_PWRGD.count_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => \N__28969\,
            sr => \N__19980\
        );

    \RSMRST_PWRGD.count_RNI_11_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16612\,
            in1 => \N__16495\,
            in2 => \N__28774\,
            in3 => \N__16723\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un12_clk_100khz_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI166B31_12_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15580\,
            in1 => \N__16816\,
            in2 => \N__15571\,
            in3 => \N__15538\,
            lcout => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\,
            ltout => \RSMRST_PWRGD.count_RNI166B31Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__16613\,
            in1 => \_gnd_net_\,
            in2 => \N__15568\,
            in3 => \N__19968\,
            lcout => \RSMRST_PWRGD.count_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => \N__28969\,
            sr => \N__19980\
        );

    \RSMRST_PWRGD.count_14_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35282\,
            ce => \N__28970\,
            sr => \N__19974\
        );

    \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16511\,
            in1 => \N__15552\,
            in2 => \_gnd_net_\,
            in3 => \N__28899\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_5_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16513\,
            lcout => \RSMRST_PWRGD.count_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35282\,
            ce => \N__28970\,
            sr => \N__19974\
        );

    \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__28901\,
            in2 => \_gnd_net_\,
            in3 => \N__16653\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => \RSMRST_PWRGD.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__28902\,
            in1 => \N__15553\,
            in2 => \N__15541\,
            in3 => \N__16512\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI812M5_11_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15607\,
            in1 => \N__28900\,
            in2 => \_gnd_net_\,
            in3 => \N__16710\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_11_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35282\,
            ce => \N__28970\,
            sr => \N__19974\
        );

    \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18436\,
            in1 => \N__28898\,
            in2 => \_gnd_net_\,
            in3 => \N__18453\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25667\,
            in2 => \N__19038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25743\,
            in1 => \N__17295\,
            in2 => \_gnd_net_\,
            in3 => \N__15601\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25747\,
            in1 => \N__17238\,
            in2 => \_gnd_net_\,
            in3 => \N__15598\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25744\,
            in1 => \_gnd_net_\,
            in2 => \N__17101\,
            in3 => \N__15595\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25748\,
            in1 => \_gnd_net_\,
            in2 => \N__15700\,
            in3 => \N__15592\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25745\,
            in1 => \_gnd_net_\,
            in2 => \N__17080\,
            in3 => \N__15589\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25749\,
            in1 => \_gnd_net_\,
            in2 => \N__17215\,
            in3 => \N__15586\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25746\,
            in1 => \_gnd_net_\,
            in2 => \N__17272\,
            in3 => \N__15583\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25750\,
            in1 => \_gnd_net_\,
            in2 => \N__15715\,
            in3 => \N__15628\,
            lcout => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25754\,
            in1 => \_gnd_net_\,
            in2 => \N__15855\,
            in3 => \N__15625\,
            lcout => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9\,
            carryout => \POWERLED.un1_count_clk_2_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25751\,
            in1 => \_gnd_net_\,
            in2 => \N__15778\,
            in3 => \N__15622\,
            lcout => \POWERLED.count_clk_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25755\,
            in1 => \_gnd_net_\,
            in2 => \N__15838\,
            in3 => \N__15619\,
            lcout => \POWERLED.count_clk_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11\,
            carryout => \POWERLED.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25752\,
            in1 => \_gnd_net_\,
            in2 => \N__15640\,
            in3 => \N__15616\,
            lcout => \POWERLED.count_clk_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12\,
            carryout => \POWERLED.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25756\,
            in1 => \_gnd_net_\,
            in2 => \N__16939\,
            in3 => \N__15613\,
            lcout => \POWERLED.count_clk_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25753\,
            in1 => \N__16960\,
            in2 => \_gnd_net_\,
            in3 => \N__15610\,
            lcout => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIN1VB_10_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__23742\,
            in1 => \N__17152\,
            in2 => \N__25619\,
            in3 => \N__17163\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI499J_4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23734\,
            in1 => \N__25590\,
            in2 => \N__15667\,
            in3 => \N__15678\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI6CAJ_5_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__25591\,
            in1 => \N__23735\,
            in2 => \N__15724\,
            in3 => \N__15735\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => \POWERLED.count_clkZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_5_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16924\,
            in2 => \N__15739\,
            in3 => \N__15714\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15736\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => \N__25618\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIEOEJ_9_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23736\,
            in1 => \N__25592\,
            in2 => \N__15649\,
            in3 => \N__15657\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => \POWERLED.count_clkZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__16923\,
            in1 => \N__15696\,
            in2 => \N__15682\,
            in3 => \N__19027\,
            lcout => \POWERLED.N_193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15679\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => \N__25618\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15658\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => \N__25618\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => \N__25570\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI4DIB_13_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23745\,
            in1 => \N__25569\,
            in2 => \N__15808\,
            in3 => \N__15819\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => \POWERLED.count_clkZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_10_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15834\,
            in1 => \N__15774\,
            in2 => \N__15859\,
            in3 => \N__15856\,
            lcout => \POWERLED.un2_count_clk_17_0_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2AHB_12_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23744\,
            in1 => \N__25568\,
            in2 => \N__15748\,
            in3 => \N__15759\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15820\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => \N__25570\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI07GB_11_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23743\,
            in1 => \N__25567\,
            in2 => \N__15799\,
            in3 => \N__15789\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => \N__25570\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18957\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => \N__20562\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18900\,
            lcout => \POWERLED.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => \N__20562\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18831\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => \N__20562\,
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17540\,
            in2 => \N__17449\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNI36763_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17519\,
            in1 => \N__18942\,
            in2 => \_gnd_net_\,
            in3 => \N__15886\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNI48863_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17509\,
            in1 => \N__18885\,
            in2 => \_gnd_net_\,
            in3 => \N__15883\,
            lcout => \POWERLED.count_off_1_3\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNI5A963_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17520\,
            in1 => \N__18816\,
            in2 => \_gnd_net_\,
            in3 => \N__15880\,
            lcout => \POWERLED.count_off_1_4\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNI6CA63_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17507\,
            in1 => \N__17572\,
            in2 => \_gnd_net_\,
            in3 => \N__15877\,
            lcout => \POWERLED.count_off_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNI7EB63_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17517\,
            in1 => \N__19243\,
            in2 => \_gnd_net_\,
            in3 => \N__15874\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNI8GC63_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17508\,
            in1 => \N__19387\,
            in2 => \_gnd_net_\,
            in3 => \N__15871\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNI9ID63_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17518\,
            in1 => \N__19345\,
            in2 => \_gnd_net_\,
            in3 => \N__15868\,
            lcout => \POWERLED.count_off_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNIAKE63_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17510\,
            in1 => \N__17398\,
            in2 => \_gnd_net_\,
            in3 => \N__15865\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNIBMF63_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17513\,
            in1 => \N__17700\,
            in2 => \_gnd_net_\,
            in3 => \N__15862\,
            lcout => \POWERLED.count_off_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNIJSS43_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17511\,
            in1 => \N__17673\,
            in2 => \_gnd_net_\,
            in3 => \N__15916\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNIKUT43_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17514\,
            in1 => \N__17628\,
            in2 => \_gnd_net_\,
            in3 => \N__15913\,
            lcout => \POWERLED.count_off_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNIL0V43_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17512\,
            in1 => \N__17601\,
            in2 => \_gnd_net_\,
            in3 => \N__15910\,
            lcout => \POWERLED.count_off_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNIM2053_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17515\,
            in1 => \N__17589\,
            in2 => \_gnd_net_\,
            in3 => \N__15907\,
            lcout => \POWERLED.count_off_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIN4153_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__17616\,
            in1 => \N__17516\,
            in2 => \_gnd_net_\,
            in3 => \N__15904\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNINZ0Z4153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17641\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35340\,
            ce => \N__20563\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILQ6NA_13_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15892\,
            in1 => \N__20532\,
            in2 => \_gnd_net_\,
            in3 => \N__15900\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => \N__20561\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNINMDQA_5_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16015\,
            in1 => \N__20531\,
            in2 => \_gnd_net_\,
            in3 => \N__16026\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => \N__20561\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNINT7NA_14_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15997\,
            in1 => \N__20533\,
            in2 => \_gnd_net_\,
            in3 => \N__16005\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16009\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => \N__20561\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIP09NA_15_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15991\,
            in1 => \N__15982\,
            in2 => \_gnd_net_\,
            in3 => \N__20534\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15990\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => \N__20561\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQOGH5_0_2_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110101"
        )
    port map (
            in0 => \N__15943\,
            in1 => \N__15960\,
            in2 => \N__18387\,
            in3 => \N__15930\,
            lcout => \PCH_PWRGD.un12_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQOGH5_2_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18334\,
            in1 => \_gnd_net_\,
            in2 => \N__15964\,
            in3 => \N__15942\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15959\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35058\,
            ce => \N__18373\,
            sr => \N__18053\
        );

    \PCH_PWRGD.count_RNI25LH5_6_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18335\,
            in1 => \N__16069\,
            in2 => \_gnd_net_\,
            in3 => \N__16081\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI0AK45_0_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16430\,
            in1 => \N__18017\,
            in2 => \_gnd_net_\,
            in3 => \N__17768\,
            lcout => \PCH_PWRGD.count_rst_14\,
            ltout => \PCH_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18336\,
            in1 => \_gnd_net_\,
            in2 => \N__16093\,
            in3 => \N__16414\,
            lcout => \PCH_PWRGD.un2_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35058\,
            ce => \N__18373\,
            sr => \N__18053\
        );

    \PCH_PWRGD.count_3_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__17769\,
            in1 => \N__18078\,
            in2 => \N__18051\,
            in3 => \N__18210\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35058\,
            ce => \N__18373\,
            sr => \N__18053\
        );

    \PCH_PWRGD.count_7_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__17782\,
            in1 => \N__17857\,
            in2 => \N__17838\,
            in3 => \N__18023\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35258\,
            ce => \N__18384\,
            sr => \N__18057\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIBA6V1_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__18021\,
            in1 => \N__17781\,
            in2 => \N__16201\,
            in3 => \N__16185\,
            lcout => \PCH_PWRGD.count_rst_9\,
            ltout => \PCH_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI02KH5_0_5_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__16174\,
            in1 => \N__18308\,
            in2 => \N__16063\,
            in3 => \N__17858\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISBO9M_3_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16060\,
            in1 => \N__16054\,
            in2 => \N__16045\,
            in3 => \N__16303\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNINHV751_2_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16042\,
            in1 => \N__16165\,
            in2 => \N__16036\,
            in3 => \N__16033\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI48MH5_7_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18307\,
            in1 => \_gnd_net_\,
            in2 => \N__17725\,
            in3 => \N__16213\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI02KH5_5_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16173\,
            in1 => \N__16207\,
            in2 => \_gnd_net_\,
            in3 => \N__18306\,
            lcout => \PCH_PWRGD.un2_count_1_axb_5\,
            ltout => \PCH_PWRGD.un2_count_1_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_5_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__18022\,
            in1 => \N__16186\,
            in2 => \N__16177\,
            in3 => \N__17783\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35258\,
            ce => \N__18384\,
            sr => \N__18057\
        );

    \PCH_PWRGD.count_RNIHQ8Q5_0_10_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110001"
        )
    port map (
            in0 => \N__16135\,
            in1 => \N__16111\,
            in2 => \N__18343\,
            in3 => \N__16149\,
            lcout => \PCH_PWRGD.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIHQ8Q5_10_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16150\,
            in1 => \N__16134\,
            in2 => \_gnd_net_\,
            in3 => \N__18300\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_10_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16148\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35197\,
            ce => \N__18386\,
            sr => \N__18041\
        );

    \PCH_PWRGD.count_1_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16344\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35197\,
            ce => \N__18386\,
            sr => \N__18041\
        );

    \PCH_PWRGD.count_12_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16125\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35197\,
            ce => \N__18386\,
            sr => \N__18041\
        );

    \PCH_PWRGD.count_RNIS5SK5_12_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16126\,
            in1 => \N__16117\,
            in2 => \_gnd_net_\,
            in3 => \N__18301\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIJ2LF3_0_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__18010\,
            in1 => \N__18466\,
            in2 => \N__18157\,
            in3 => \N__29971\,
            lcout => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOLFH5_1_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16345\,
            in2 => \N__16336\,
            in3 => \N__16333\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI6BNH5_8_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16266\,
            in1 => \N__16312\,
            in2 => \_gnd_net_\,
            in3 => \N__18315\,
            lcout => \PCH_PWRGD.un2_count_1_axb_8\,
            ltout => \PCH_PWRGD.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNIEG9V1_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16278\,
            in1 => \N__18024\,
            in2 => \N__16315\,
            in3 => \N__17804\,
            lcout => \PCH_PWRGD.count_rst_6\,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI6BNH5_0_8_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__16267\,
            in1 => \N__18316\,
            in2 => \N__16306\,
            in3 => \N__16253\,
            lcout => \PCH_PWRGD.un12_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_8_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16293\,
            in1 => \N__18025\,
            in2 => \N__16282\,
            in3 => \N__17808\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35260\,
            ce => \N__18367\,
            sr => \N__18058\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNIFIAV1_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__17805\,
            in1 => \N__16254\,
            in2 => \N__16240\,
            in3 => \N__18027\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI8EOH5_9_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18368\,
            in2 => \N__16258\,
            in3 => \N__16219\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => \PCH_PWRGD.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_9_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__17806\,
            in1 => \N__16236\,
            in2 => \N__16222\,
            in3 => \N__18028\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35260\,
            ce => \N__18367\,
            sr => \N__18058\
        );

    \PCH_PWRGD.count_0_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16437\,
            in1 => \N__18026\,
            in2 => \_gnd_net_\,
            in3 => \N__17807\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35260\,
            ce => \N__18367\,
            sr => \N__18058\
        );

    \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16773\,
            in1 => \N__19948\,
            in2 => \N__16795\,
            in3 => \N__18707\,
            lcout => \RSMRST_PWRGD.count_rst_14\,
            ltout => \RSMRST_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIMCS06_9_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16380\,
            in2 => \N__16393\,
            in3 => \N__28933\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_9\,
            ltout => \RSMRST_PWRGD.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_9_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16774\,
            in1 => \N__19951\,
            in2 => \N__16390\,
            in3 => \N__18711\,
            lcout => \RSMRST_PWRGD.count_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35198\,
            ce => \N__28965\,
            sr => \N__19978\
        );

    \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__16387\,
            in1 => \N__16381\,
            in2 => \N__28960\,
            in3 => \N__16757\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16758\,
            in1 => \N__19949\,
            in2 => \N__16741\,
            in3 => \N__18708\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.count_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIV86M5_10_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16357\,
            in2 => \N__16363\,
            in3 => \N__28934\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => \RSMRST_PWRGD.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_10_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16740\,
            in1 => \N__19950\,
            in2 => \N__16360\,
            in3 => \N__18710\,
            lcout => \RSMRST_PWRGD.count_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35198\,
            ce => \N__28965\,
            sr => \N__19978\
        );

    \RSMRST_PWRGD.count_13_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__18709\,
            in1 => \N__16695\,
            in2 => \N__19977\,
            in3 => \N__16678\,
            lcout => \RSMRST_PWRGD.count_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35198\,
            ce => \N__28965\,
            sr => \N__19978\
        );

    \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16631\,
            in2 => \N__16618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19938\,
            in1 => \N__16594\,
            in2 => \_gnd_net_\,
            in3 => \N__16576\,
            lcout => \RSMRST_PWRGD.count_rst_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19945\,
            in1 => \N__16572\,
            in2 => \_gnd_net_\,
            in3 => \N__16555\,
            lcout => \RSMRST_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16550\,
            in2 => \_gnd_net_\,
            in3 => \N__16525\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19946\,
            in1 => \N__16522\,
            in2 => \_gnd_net_\,
            in3 => \N__16498\,
            lcout => \RSMRST_PWRGD.count_rst_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19939\,
            in1 => \N__16494\,
            in2 => \_gnd_net_\,
            in3 => \N__16474\,
            lcout => \RSMRST_PWRGD.count_rst_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19947\,
            in1 => \N__28764\,
            in2 => \_gnd_net_\,
            in3 => \N__16471\,
            lcout => \RSMRST_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16466\,
            in2 => \_gnd_net_\,
            in3 => \N__16441\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_7\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16791\,
            in2 => \_gnd_net_\,
            in3 => \N__16762\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16759\,
            in2 => \_gnd_net_\,
            in3 => \N__16726\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19913\,
            in1 => \N__16722\,
            in2 => \_gnd_net_\,
            in3 => \N__16702\,
            lcout => \RSMRST_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19899\,
            in1 => \N__16639\,
            in2 => \_gnd_net_\,
            in3 => \N__16699\,
            lcout => \RSMRST_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16694\,
            in2 => \_gnd_net_\,
            in3 => \N__16663\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19900\,
            in1 => \N__16660\,
            in2 => \_gnd_net_\,
            in3 => \N__16645\,
            lcout => \RSMRST_PWRGD.count_rst_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16864\,
            in1 => \N__19901\,
            in2 => \_gnd_net_\,
            in3 => \N__16642\,
            lcout => \RSMRST_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIA43M5_12_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16849\,
            in1 => \N__28909\,
            in2 => \_gnd_net_\,
            in3 => \N__16829\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_15_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16881\,
            lcout => \RSMRST_PWRGD.count_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35281\,
            ce => \N__28954\,
            sr => \N__19961\
        );

    \RSMRST_PWRGD.count_12_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16830\,
            lcout => \RSMRST_PWRGD.count_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35281\,
            ce => \N__28954\,
            sr => \N__19961\
        );

    \RSMRST_PWRGD.count_RNIGD6M5_15_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16882\,
            in1 => \N__16873\,
            in2 => \_gnd_net_\,
            in3 => \N__28955\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21909\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28045\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_240_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__21957\,
            in1 => \N__19914\,
            in2 => \N__16867\,
            in3 => \N__30999\,
            lcout => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\,
            ltout => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010001"
        )
    port map (
            in0 => \N__16860\,
            in1 => \N__16845\,
            in2 => \N__16834\,
            in3 => \N__16831\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__28044\,
            in1 => \N__21956\,
            in2 => \_gnd_net_\,
            in3 => \N__21908\,
            lcout => \RSMRST_PWRGD.N_423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI268J_3_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25583\,
            in1 => \N__16801\,
            in2 => \N__23732\,
            in3 => \N__16809\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35316\,
            ce => \N__25620\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI6GJB_14_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25584\,
            in1 => \N__16888\,
            in2 => \N__23733\,
            in3 => \N__16896\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8JKB_15_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__16903\,
            in1 => \N__25585\,
            in2 => \N__23737\,
            in3 => \N__16911\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => \POWERLED.count_clkZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_15_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25668\,
            in1 => \N__16954\,
            in2 => \N__16942\,
            in3 => \N__16938\,
            lcout => \POWERLED.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI9LLG_0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__25639\,
            in1 => \N__23687\,
            in2 => \N__18991\,
            in3 => \N__25582\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16912\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35316\,
            ce => \N__25620\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16897\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35316\,
            ce => \N__25620\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5UUJ4_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__20635\,
            in1 => \N__17020\,
            in2 => \N__22831\,
            in3 => \N__22736\,
            lcout => \POWERLED.func_state_1_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__20907\,
            in1 => \N__20345\,
            in2 => \N__24579\,
            in3 => \N__17353\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_1_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22734\,
            in2 => \_gnd_net_\,
            in3 => \N__24564\,
            lcout => \POWERLED.func_state_RNI_1Z0Z_1\,
            ltout => \POWERLED.func_state_RNI_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPS253_0_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__19066\,
            in1 => \N__20908\,
            in2 => \N__17023\,
            in3 => \N__20347\,
            lcout => \POWERLED.func_state_1_m2_ns_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22332\,
            in1 => \N__22735\,
            in2 => \N__17380\,
            in3 => \N__24421\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_0_1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__24565\,
            in1 => \N__20346\,
            in2 => \N__17014\,
            in3 => \N__36146\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1E8A4_0_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17011\,
            in1 => \N__19065\,
            in2 => \N__17005\,
            in3 => \N__17312\,
            lcout => \POWERLED.func_state_RNI1E8A4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_0_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100101011"
        )
    port map (
            in0 => \N__22737\,
            in1 => \N__20909\,
            in2 => \N__24580\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_func_state25_4_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8FBJ_6_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23739\,
            in1 => \N__25587\,
            in2 => \N__16990\,
            in3 => \N__17001\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => \N__25617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNICLDJ_8_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23741\,
            in1 => \N__25589\,
            in2 => \N__16969\,
            in3 => \N__16980\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => \N__25617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAICJ_7_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23740\,
            in1 => \N__25588\,
            in2 => \N__17122\,
            in3 => \N__17133\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => \N__25617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAMLG_1_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__23738\,
            in1 => \N__25586\,
            in2 => \N__17110\,
            in3 => \N__19003\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => \POWERLED.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25760\,
            in2 => \N__17113\,
            in3 => \N__25680\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => \N__25617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17038\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => \N__25579\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_4_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17076\,
            in2 => \_gnd_net_\,
            in3 => \N__17097\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_2_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__17096\,
            in1 => \N__17244\,
            in2 => \N__17296\,
            in3 => \N__17270\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_6_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__17209\,
            in1 => \N__17075\,
            in2 => \N__17059\,
            in3 => \N__17052\,
            lcout => \POWERLED.count_clk_RNIZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_7_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17210\,
            in2 => \N__17056\,
            in3 => \N__17227\,
            lcout => \POWERLED.N_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI037J_2_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__17044\,
            in1 => \N__23704\,
            in2 => \N__25581\,
            in3 => \N__17037\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => \POWERLED.count_clkZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_2_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__17278\,
            in1 => \N__17271\,
            in2 => \N__17248\,
            in3 => \N__17245\,
            lcout => \POWERLED.N_385\,
            ltout => \POWERLED.N_385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_1_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17221\,
            in1 => \N__17211\,
            in2 => \N__17188\,
            in3 => \N__19028\,
            lcout => \POWERLED.count_clk_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIP7PD2_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001010"
        )
    port map (
            in0 => \N__22475\,
            in1 => \N__32918\,
            in2 => \N__29728\,
            in3 => \N__27971\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIFAGK3_0_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__27972\,
            in1 => \N__22336\,
            in2 => \N__17185\,
            in3 => \N__17182\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIH0GD5_1_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__23986\,
            in1 => \N__30992\,
            in2 => \N__17173\,
            in3 => \N__17320\,
            lcout => \POWERLED.count_clk_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_en_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__27973\,
            in1 => \_gnd_net_\,
            in2 => \N__31006\,
            in3 => \N__22476\,
            lcout => \POWERLED.func_state_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17170\,
            lcout => \POWERLED.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => \N__25580\,
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNIEHDM1_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__29107\,
            in1 => \N__29032\,
            in2 => \N__29062\,
            in3 => \N__29125\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNICU6N2_0_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17448\,
            in2 => \_gnd_net_\,
            in3 => \N__17521\,
            lcout => OPEN,
            ltout => \POWERLED.count_off_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIO3ABA_0_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17419\,
            in2 => \N__17392\,
            in3 => \N__20501\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17389\,
            in1 => \N__24327\,
            in2 => \N__22777\,
            in3 => \N__17376\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_336_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_0_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24572\,
            in2 => \_gnd_net_\,
            in3 => \N__20889\,
            lcout => \POWERLED.func_state_RNI_3Z0Z_0\,
            ltout => \POWERLED.func_state_RNI_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIC1SE1_0_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22722\,
            in1 => \N__22828\,
            in2 => \N__17383\,
            in3 => \N__17375\,
            lcout => OPEN,
            ltout => \POWERLED.N_321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICU6N2_1_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__23982\,
            in1 => \N__17352\,
            in2 => \N__17356\,
            in3 => \N__19132\,
            lcout => \POWERLED.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__24573\,
            in1 => \N__23981\,
            in2 => \N__22684\,
            in3 => \N__17351\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__19111\,
            in1 => \N__17329\,
            in2 => \N__17323\,
            in3 => \N__17319\,
            lcout => \POWERLED.un1_func_state25_6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_3_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19344\,
            in1 => \N__19386\,
            in2 => \N__18889\,
            in3 => \N__18820\,
            lcout => \POWERLED.un34_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17617\,
            in1 => \N__17447\,
            in2 => \N__17605\,
            in3 => \N__17590\,
            lcout => \POWERLED.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNICU6N2_1_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__17446\,
            in1 => \N__17542\,
            in2 => \_gnd_net_\,
            in3 => \N__17504\,
            lcout => OPEN,
            ltout => \POWERLED.count_off_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIP4ABA_1_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17527\,
            in2 => \N__17578\,
            in3 => \N__20500\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => \POWERLED.count_offZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18946\,
            in1 => \N__19242\,
            in2 => \N__17575\,
            in3 => \N__17571\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_10_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17557\,
            in1 => \N__17551\,
            in2 => \N__17545\,
            in3 => \N__17707\,
            lcout => \POWERLED.count_off_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__17445\,
            in1 => \N__17541\,
            in2 => \_gnd_net_\,
            in3 => \N__17506\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => \N__20535\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__17505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17444\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => \N__20535\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17407\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35337\,
            ce => \N__20545\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIV2IQA_9_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20511\,
            in1 => \N__17413\,
            in2 => \_gnd_net_\,
            in3 => \N__17406\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => \POWERLED.count_offZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_10_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17674\,
            in1 => \N__17629\,
            in2 => \N__17710\,
            in3 => \N__17701\,
            lcout => \POWERLED.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI8DNOA_10_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20512\,
            in1 => \N__17680\,
            in2 => \_gnd_net_\,
            in3 => \N__17688\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35337\,
            ce => \N__20545\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHK4NA_11_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20513\,
            in1 => \N__17653\,
            in2 => \_gnd_net_\,
            in3 => \N__17661\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17662\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35337\,
            ce => \N__20545\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJN5NA_12_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20514\,
            in1 => \N__17647\,
            in2 => \_gnd_net_\,
            in3 => \N__17640\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__17812\,
            in1 => \N__18095\,
            in2 => \N__18561\,
            in3 => \N__18599\,
            lcout => \PCH_PWRGD.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34991\,
            ce => \N__30948\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__18553\,
            in1 => \N__18522\,
            in2 => \N__18100\,
            in3 => \N__17813\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34991\,
            ce => \N__30948\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__17811\,
            in1 => \N__18598\,
            in2 => \N__18562\,
            in3 => \N__18094\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI02502_0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__23725\,
            in1 => \_gnd_net_\,
            in2 => \N__18124\,
            in3 => \N__18121\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18115\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2857_i\,
            ltout => \PCH_PWRGD.N_2857_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__18099\,
            in1 => \N__18523\,
            in2 => \N__18112\,
            in3 => \N__17810\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.curr_state_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI13502_1_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18109\,
            in2 => \N__18103\,
            in3 => \N__23724\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18082\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2859_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNI964V1_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__18079\,
            in1 => \N__17929\,
            in2 => \N__18206\,
            in3 => \N__17814\,
            lcout => \PCH_PWRGD.count_rst_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18516\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => \PCH_PWRGD.count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNIDE8V1_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__17863\,
            in1 => \N__17839\,
            in2 => \N__17818\,
            in3 => \N__17815\,
            lcout => \PCH_PWRGD.count_rst_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISRHH5_3_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18424\,
            in1 => \N__18399\,
            in2 => \_gnd_net_\,
            in3 => \N__18369\,
            lcout => \PCH_PWRGD.un2_count_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNO_0_1_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18163\,
            in2 => \_gnd_net_\,
            in3 => \N__23728\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__31037\,
            in1 => \N__31065\,
            in2 => \N__18178\,
            in3 => \N__25003\,
            lcout => \VPP_VDDQ.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35083\,
            ce => \N__30945\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI67MK_1_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__25002\,
            in1 => \N__31036\,
            in2 => \N__18175\,
            in3 => \N__23726\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => \VPP_VDDQ.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18166\,
            in3 => \N__31064\,
            lcout => \VPP_VDDQ.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35083\,
            ce => \N__30945\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIJN8A3_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__18600\,
            in1 => \N__18130\,
            in2 => \N__18577\,
            in3 => \N__30996\,
            lcout => \PCH_PWRGD.delayed_vccin_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI1IPC1_0_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18504\,
            in1 => \N__18479\,
            in2 => \N__18156\,
            in3 => \N__27981\,
            lcout => \PCH_PWRGD.curr_state_RNI1IPC1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__21700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31167\,
            lcout => \VPP_VDDQ.N_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI1IPC1_0_0_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__18503\,
            in1 => \N__18532\,
            in2 => \_gnd_net_\,
            in3 => \N__27982\,
            lcout => \PCH_PWRGD.N_277_0\,
            ltout => \PCH_PWRGD.N_277_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__18601\,
            in1 => \N__18576\,
            in2 => \N__18580\,
            in3 => \N__30997\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_0_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18480\,
            in2 => \_gnd_net_\,
            in3 => \N__18560\,
            lcout => \PCH_PWRGD.N_413\,
            ltout => \PCH_PWRGD.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__27983\,
            in1 => \_gnd_net_\,
            in2 => \N__18526\,
            in3 => \N__18502\,
            lcout => \PCH_PWRGD.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI1IPC1_1_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__18505\,
            in1 => \N__18481\,
            in2 => \_gnd_net_\,
            in3 => \N__27980\,
            lcout => \PCH_PWRGD.N_278_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_3_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18457\,
            lcout => \RSMRST_PWRGD.count_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35088\,
            ce => \N__28961\,
            sr => \N__19975\
        );

    \RSMRST_PWRGD.count_7_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28800\,
            lcout => \RSMRST_PWRGD.count_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35088\,
            ce => \N__28961\,
            sr => \N__19975\
        );

    \POWERLED.count_13_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20275\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35093\,
            ce => \N__30944\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_4_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20133\,
            lcout => \POWERLED.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35093\,
            ce => \N__30944\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20113\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35093\,
            ce => \N__30944\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20092\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35093\,
            ce => \N__30944\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20244\,
            in3 => \N__26016\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35122\,
            ce => \N__30947\,
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26805\,
            in2 => \N__25876\,
            in3 => \N__29106\,
            lcout => \POWERLED.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35122\,
            ce => \N__30947\,
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIF5D5_0_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23624\,
            in2 => \N__26817\,
            in3 => \N__25871\,
            lcout => \POWERLED.count_0_sqmuxa_i\,
            ltout => \POWERLED.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_0_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__26018\,
            in1 => \_gnd_net_\,
            in2 => \N__18628\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGAFE_0_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18625\,
            in2 => \N__18619\,
            in3 => \N__23625\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => \POWERLED.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_1_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20220\,
            in2 => \N__18616\,
            in3 => \N__25976\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIHBFE_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18607\,
            in2 => \N__18613\,
            in3 => \N__23626\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => \POWERLED.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__26017\,
            in1 => \_gnd_net_\,
            in2 => \N__18610\,
            in3 => \N__20219\,
            lcout => \POWERLED.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35122\,
            ce => \N__30947\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18640\,
            in1 => \N__18724\,
            in2 => \_gnd_net_\,
            in3 => \N__23556\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28034\,
            in2 => \N__18742\,
            in3 => \N__21942\,
            lcout => \curr_state_RNIR5QD1_0_0\,
            ltout => \curr_state_RNIR5QD1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__21944\,
            in1 => \N__21892\,
            in2 => \N__18739\,
            in3 => \N__18712\,
            lcout => \RSMRST_PWRGD.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => \N__30954\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__24186\,
            in1 => \N__21946\,
            in2 => \N__18718\,
            in3 => \N__21897\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.m4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18736\,
            in2 => \N__18730\,
            in3 => \N__23555\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__18717\,
            in1 => \N__20004\,
            in2 => \N__18727\,
            in3 => \N__21898\,
            lcout => \RSMRST_PWRGD.curr_state_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__21943\,
            in1 => \N__21893\,
            in2 => \N__20005\,
            in3 => \N__18713\,
            lcout => \RSMRST_PWRGD.curr_state_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => \N__30954\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_fast_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28033\,
            in2 => \N__21907\,
            in3 => \N__21945\,
            lcout => \RSMRST_PWRGD_RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => \N__30954\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIKKSP_10_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20065\,
            in1 => \N__18634\,
            in2 => \_gnd_net_\,
            in3 => \N__23637\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20064\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34992\,
            ce => \N__30946\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNITEFN_2_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19753\,
            in1 => \N__18778\,
            in2 => \_gnd_net_\,
            in3 => \N__23638\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19752\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34992\,
            ce => \N__30946\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNITF4O_11_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20053\,
            in1 => \N__18772\,
            in2 => \_gnd_net_\,
            in3 => \N__23639\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20049\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34992\,
            ce => \N__30946\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIVHGN_3_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19732\,
            in1 => \N__18766\,
            in2 => \_gnd_net_\,
            in3 => \N__23640\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19731\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34992\,
            ce => \N__30946\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIVI5O_12_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20029\,
            in1 => \N__18760\,
            in2 => \_gnd_net_\,
            in3 => \N__23669\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20028\,
            lcout => \POWERLED.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35219\,
            ce => \N__30950\,
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI3P6L_0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18754\,
            in1 => \N__23668\,
            in2 => \_gnd_net_\,
            in3 => \N__25837\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19039\,
            in2 => \N__25776\,
            in3 => \N__25675\,
            lcout => \POWERLED.count_clk_RNIZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25769\,
            lcout => \POWERLED.count_clk_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHDAQA_2_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20484\,
            in1 => \N__18979\,
            in2 => \_gnd_net_\,
            in3 => \N__18967\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJGBQA_3_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18922\,
            in1 => \N__18910\,
            in2 => \_gnd_net_\,
            in3 => \N__20485\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILJCQA_4_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__20486\,
            in1 => \_gnd_net_\,
            in2 => \N__18856\,
            in3 => \N__18841\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_0_i_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__21859\,
            in1 => \N__22422\,
            in2 => \N__24227\,
            in3 => \N__23667\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPPHK1_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__22657\,
            in1 => \N__21858\,
            in2 => \N__24228\,
            in3 => \N__24153\,
            lcout => \POWERLED_un1_clk_100khz_52_and_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_2_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22630\,
            in2 => \_gnd_net_\,
            in3 => \N__22424\,
            lcout => OPEN,
            ltout => \POWERLED.N_359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110111"
        )
    port map (
            in0 => \N__24211\,
            in1 => \N__22100\,
            in2 => \N__18781\,
            in3 => \N__21856\,
            lcout => \POWERLED.N_171\,
            ltout => \POWERLED.N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__22632\,
            in1 => \N__22425\,
            in2 => \N__19069\,
            in3 => \N__23666\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_oZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.slp_s3n_signal_i_0_o3_2_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101111111"
        )
    port map (
            in0 => \N__24215\,
            in1 => \N__22631\,
            in2 => \N__24156\,
            in3 => \N__21855\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22629\,
            in2 => \_gnd_net_\,
            in3 => \N__22423\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_0_o3_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110111"
        )
    port map (
            in0 => \N__24210\,
            in1 => \N__22101\,
            in2 => \N__19054\,
            in3 => \N__21857\,
            lcout => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19149\,
            in1 => \N__22222\,
            in2 => \N__20910\,
            in3 => \N__20727\,
            lcout => \POWERLED.func_state_RNI3IN21Z0Z_0\,
            ltout => \POWERLED.func_state_RNI3IN21Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIC1SE1_0_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22810\,
            in2 => \N__19051\,
            in3 => \N__27011\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m2_ns_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIGMCP2_1_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__24513\,
            in1 => \N__30103\,
            in2 => \N__19048\,
            in3 => \N__22739\,
            lcout => \POWERLED.func_state_1_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20898\,
            lcout => \POWERLED.N_2905_i\,
            ltout => \POWERLED.N_2905_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19045\,
            in3 => \N__24492\,
            lcout => \POWERLED.N_175\,
            ltout => \POWERLED.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__22740\,
            in1 => \N__19150\,
            in2 => \N__19042\,
            in3 => \N__27012\,
            lcout => \POWERLED.func_state_1_ss0_i_0_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_1_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__27013\,
            in1 => \_gnd_net_\,
            in2 => \N__19128\,
            in3 => \N__19148\,
            lcout => \POWERLED.N_343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_ss0_i_0_a2_3_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__22421\,
            in1 => \N__22641\,
            in2 => \_gnd_net_\,
            in3 => \N__24322\,
            lcout => \POWERLED.func_state_1_ss0_i_0_a2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNITIO1D_1_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__31153\,
            in1 => \N__19660\,
            in2 => \N__19225\,
            in3 => \N__20361\,
            lcout => \POWERLED.func_state\,
            ltout => \POWERLED.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19135\,
            in3 => \N__22738\,
            lcout => \POWERLED.func_state_RNI_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_1_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__31154\,
            in1 => \N__22607\,
            in2 => \N__22315\,
            in3 => \N__27034\,
            lcout => \POWERLED.un1_func_state25_6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_0_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22284\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIESP71_1_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20307\,
            in1 => \N__22108\,
            in2 => \N__19099\,
            in3 => \N__24512\,
            lcout => \POWERLED.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__19096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31156\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__22606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22410\,
            lcout => \POWERLED.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__20362\,
            in1 => \N__19224\,
            in2 => \N__19668\,
            in3 => \N__31155\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIKUJM1_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__24510\,
            in1 => \N__22612\,
            in2 => \N__19213\,
            in3 => \N__22939\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_0_2\,
            ltout => \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__19183\,
            in1 => \N__19189\,
            in2 => \N__19198\,
            in3 => \N__19174\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35317\,
            ce => 'H',
            sr => \N__32468\
        );

    \POWERLED.dutycycle_RNI_1_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__24509\,
            in1 => \N__27050\,
            in2 => \_gnd_net_\,
            in3 => \N__29345\,
            lcout => OPEN,
            ltout => \POWERLED.N_238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIML1B1_2_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011111"
        )
    port map (
            in0 => \N__22408\,
            in1 => \N__20416\,
            in2 => \N__19195\,
            in3 => \N__27946\,
            lcout => OPEN,
            ltout => \POWERLED.N_118_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIS3763_2_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29941\,
            in2 => \N__19192\,
            in3 => \N__30142\,
            lcout => \POWERLED.dutycycle_RNIS3763Z0Z_2\,
            ltout => \POWERLED.dutycycle_RNIS3763Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI0RNB6_2_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__19182\,
            in1 => \N__19173\,
            in2 => \N__19162\,
            in3 => \N__19159\,
            lcout => \POWERLED.dutycycle\,
            ltout => \POWERLED.dutycycle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5DLR_2_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22407\,
            in2 => \N__19153\,
            in3 => \N__22608\,
            lcout => \POWERLED.g0_13_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_1_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__22409\,
            in1 => \N__24508\,
            in2 => \N__22633\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIAQAN1_0_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__19294\,
            in1 => \N__20327\,
            in2 => \N__20914\,
            in3 => \N__36149\,
            lcout => OPEN,
            ltout => \POWERLED.g0_i_a6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIGGI33_0_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__24323\,
            in1 => \N__19267\,
            in2 => \N__19288\,
            in3 => \N__20746\,
            lcout => OPEN,
            ltout => \POWERLED.g2_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI9EN09_7_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__19276\,
            in1 => \N__29964\,
            in2 => \N__19285\,
            in3 => \N__30141\,
            lcout => \POWERLED.dutycycle_en_5_0_0\,
            ltout => \POWERLED.dutycycle_en_5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIAN5BA_7_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__19251\,
            in1 => \N__32942\,
            in2 => \N__19282\,
            in3 => \N__22899\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => \POWERLED.dutycycleZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJFV14_7_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101110101"
        )
    port map (
            in0 => \N__32943\,
            in1 => \N__24324\,
            in2 => \N__19279\,
            in3 => \N__20392\,
            lcout => \POWERLED.dutycycle_eena_5_0_N_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_7_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37446\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_7\,
            ltout => \POWERLED.dutycycle_RNI_6Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_0_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__20752\,
            in1 => \N__20674\,
            in2 => \N__19270\,
            in3 => \N__36148\,
            lcout => \POWERLED.g0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__19261\,
            in1 => \N__22900\,
            in2 => \N__19255\,
            in3 => \N__32944\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \N__32421\
        );

    \POWERLED.count_off_RNIPPEQA_6_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19408\,
            in1 => \N__19393\,
            in2 => \_gnd_net_\,
            in3 => \N__20518\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19407\,
            lcout => \POWERLED.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => \N__20546\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIRSFQA_7_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19366\,
            in1 => \N__19351\,
            in2 => \_gnd_net_\,
            in3 => \N__20519\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19365\,
            lcout => \POWERLED.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => \N__20546\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNITVGQA_8_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19324\,
            in1 => \N__19309\,
            in2 => \_gnd_net_\,
            in3 => \N__20520\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19323\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => \N__20546\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_1_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__36005\,
            in1 => \N__24607\,
            in2 => \_gnd_net_\,
            in3 => \N__24578\,
            lcout => \POWERLED.func_state_1_m2s2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_1_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36004\,
            lcout => \POWERLED.N_175_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIUGTH4_1_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19300\,
            in1 => \N__21148\,
            in2 => \_gnd_net_\,
            in3 => \N__23662\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => \HDA_STRAP.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101011111010"
        )
    port map (
            in0 => \N__21186\,
            in1 => \N__21175\,
            in2 => \N__19303\,
            in3 => \N__21119\,
            lcout => \HDA_STRAP.curr_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34850\,
            ce => \N__30942\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110101010"
        )
    port map (
            in0 => \N__19420\,
            in1 => \N__19435\,
            in2 => \N__19450\,
            in3 => \N__23664\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000101"
        )
    port map (
            in0 => \N__19433\,
            in1 => \N__19446\,
            in2 => \N__21190\,
            in3 => \N__21120\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34850\,
            ce => \N__30942\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIVHTH4_2_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__19465\,
            in1 => \N__19456\,
            in2 => \_gnd_net_\,
            in3 => \N__23663\,
            lcout => \HDA_STRAP.curr_state_i_2\,
            ltout => \HDA_STRAP.curr_state_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__21185\,
            in1 => \N__19445\,
            in2 => \N__19459\,
            in3 => \N__21118\,
            lcout => \HDA_STRAP.i4_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNI_0_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21171\,
            in2 => \_gnd_net_\,
            in3 => \N__21805\,
            lcout => \HDA_STRAP.N_208\,
            ltout => \HDA_STRAP.N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__19434\,
            in1 => \_gnd_net_\,
            in2 => \N__19423\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.HDA_SDO_ATP_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34850\,
            ce => \N__30942\,
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21406\,
            in2 => \N__21568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21342\,
            in2 => \_gnd_net_\,
            in3 => \N__19414\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21211\,
            in2 => \_gnd_net_\,
            in3 => \N__19411\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21361\,
            in2 => \_gnd_net_\,
            in3 => \N__19510\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21385\,
            in2 => \_gnd_net_\,
            in3 => \N__19507\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21427\,
            in3 => \N__19504\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21439\,
            in2 => \_gnd_net_\,
            in3 => \N__19501\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__35018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21451\,
            in2 => \_gnd_net_\,
            in3 => \N__19498\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__35018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21478\,
            in2 => \_gnd_net_\,
            in3 => \N__19495\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21465\,
            in2 => \_gnd_net_\,
            in3 => \N__19492\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21490\,
            in2 => \_gnd_net_\,
            in3 => \N__19489\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21025\,
            in2 => \_gnd_net_\,
            in3 => \N__19486\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21052\,
            in2 => \_gnd_net_\,
            in3 => \N__19537\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21039\,
            in2 => \_gnd_net_\,
            in3 => \N__19534\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21064\,
            in2 => \_gnd_net_\,
            in3 => \N__19531\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21286\,
            in2 => \_gnd_net_\,
            in3 => \N__19528\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__35046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21300\,
            in2 => \_gnd_net_\,
            in3 => \N__19525\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21313\,
            in2 => \_gnd_net_\,
            in3 => \N__19522\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21325\,
            in2 => \_gnd_net_\,
            in3 => \N__19519\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21249\,
            in2 => \_gnd_net_\,
            in3 => \N__19516\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21235\,
            in2 => \_gnd_net_\,
            in3 => \N__19513\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21262\,
            in2 => \_gnd_net_\,
            in3 => \N__19564\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21274\,
            in2 => \_gnd_net_\,
            in3 => \N__19561\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19681\,
            in2 => \_gnd_net_\,
            in3 => \N__19558\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__35084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19708\,
            in3 => \N__19555\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19696\,
            in3 => \N__19552\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19717\,
            in2 => \_gnd_net_\,
            in3 => \N__19549\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19579\,
            in2 => \_gnd_net_\,
            in3 => \N__19546\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19606\,
            in2 => \_gnd_net_\,
            in3 => \N__19543\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19593\,
            in2 => \_gnd_net_\,
            in3 => \N__19540\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19618\,
            in2 => \_gnd_net_\,
            in3 => \N__19720\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19716\,
            in1 => \N__19704\,
            in2 => \N__19695\,
            in3 => \N__19680\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHPASE_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__31151\,
            in1 => \N__19664\,
            in2 => \N__19630\,
            in3 => \N__20592\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__20593\,
            in1 => \N__19629\,
            in2 => \N__19669\,
            in3 => \N__31152\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19617\,
            in1 => \N__19605\,
            in2 => \N__19594\,
            in3 => \N__19578\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23383\,
            lcout => \VPP_VDDQ.N_2897_i\,
            ltout => \VPP_VDDQ.N_2897_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__21693\,
            in1 => \_gnd_net_\,
            in2 => \N__19567\,
            in3 => \N__23437\,
            lcout => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22016\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23575\,
            lcout => suswarn_n,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35176\,
            ce => \N__34443\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI1LHN_4_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__23570\,
            in1 => \_gnd_net_\,
            in2 => \N__20134\,
            in3 => \N__20017\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20000\,
            in2 => \_gnd_net_\,
            in3 => \N__23569\,
            lcout => \RSMRST_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI1M6O_13_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23571\,
            in1 => \N__19783\,
            in2 => \_gnd_net_\,
            in3 => \N__20274\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI3OIN_5_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19774\,
            in1 => \N__23572\,
            in2 => \_gnd_net_\,
            in3 => \N__20109\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI3P7O_14_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23573\,
            in1 => \N__20155\,
            in2 => \_gnd_net_\,
            in3 => \N__20170\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI5RJN_6_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19765\,
            in1 => \N__23574\,
            in2 => \_gnd_net_\,
            in3 => \N__20091\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26022\,
            in2 => \N__25983\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20226\,
            in1 => \N__25934\,
            in2 => \_gnd_net_\,
            in3 => \N__19735\,
            lcout => \POWERLED.count_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20245\,
            in1 => \N__26396\,
            in2 => \_gnd_net_\,
            in3 => \N__19723\,
            lcout => \POWERLED.count_1_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2\,
            carryout => \POWERLED.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNID629_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20224\,
            in1 => \N__26357\,
            in2 => \_gnd_net_\,
            in3 => \N__20116\,
            lcout => \POWERLED.count_1_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3\,
            carryout => \POWERLED.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20246\,
            in1 => \N__26319\,
            in2 => \_gnd_net_\,
            in3 => \N__20095\,
            lcout => \POWERLED.count_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20225\,
            in1 => \N__26282\,
            in2 => \_gnd_net_\,
            in3 => \N__20077\,
            lcout => \POWERLED.count_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20247\,
            in1 => \N__26241\,
            in2 => \_gnd_net_\,
            in3 => \N__20074\,
            lcout => \POWERLED.count_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20227\,
            in1 => \N__26202\,
            in2 => \_gnd_net_\,
            in3 => \N__20071\,
            lcout => \POWERLED.count_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20223\,
            in1 => \N__26157\,
            in2 => \_gnd_net_\,
            in3 => \N__20068\,
            lcout => \POWERLED.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20248\,
            in1 => \_gnd_net_\,
            in2 => \N__26637\,
            in3 => \N__20056\,
            lcout => \POWERLED.count_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20222\,
            in1 => \_gnd_net_\,
            in2 => \N__26604\,
            in3 => \N__20032\,
            lcout => \POWERLED.count_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20249\,
            in1 => \N__26558\,
            in2 => \_gnd_net_\,
            in3 => \N__20020\,
            lcout => \POWERLED.count_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20221\,
            in1 => \N__26525\,
            in2 => \_gnd_net_\,
            in3 => \N__20257\,
            lcout => \POWERLED.count_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20250\,
            in1 => \N__26493\,
            in2 => \_gnd_net_\,
            in3 => \N__20254\,
            lcout => \POWERLED.count_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__20251\,
            in2 => \_gnd_net_\,
            in3 => \N__20173\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20166\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35218\,
            ce => \N__30951\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5QAN_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000101"
        )
    port map (
            in0 => \N__24550\,
            in1 => \N__22289\,
            in2 => \N__36147\,
            in3 => \N__22634\,
            lcout => \POWERLED.g3_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6RAN_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__22290\,
            in1 => \N__22471\,
            in2 => \_gnd_net_\,
            in3 => \N__24548\,
            lcout => OPEN,
            ltout => \POWERLED.N_8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIECGS1_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__22292\,
            in1 => \N__20335\,
            in2 => \N__20146\,
            in3 => \N__20902\,
            lcout => \POWERLED.g0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3NQD_1_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__22470\,
            in1 => \N__24549\,
            in2 => \_gnd_net_\,
            in3 => \N__36112\,
            lcout => OPEN,
            ltout => \POWERLED.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJP5O2_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22639\,
            in2 => \N__20143\,
            in3 => \N__20140\,
            lcout => \POWERLED.g0_8_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20903\,
            in1 => \N__22472\,
            in2 => \N__22642\,
            in3 => \N__22291\,
            lcout => OPEN,
            ltout => \POWERLED.N_331_N_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIIO5O2_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110011"
        )
    port map (
            in0 => \N__22473\,
            in1 => \N__22638\,
            in2 => \N__20401\,
            in3 => \N__20398\,
            lcout => \POWERLED.g3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__22288\,
            in1 => \N__24315\,
            in2 => \N__20344\,
            in3 => \N__22096\,
            lcout => \POWERLED.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_m1_0_a2_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22316\,
            in1 => \N__24252\,
            in2 => \N__24154\,
            in3 => \N__20343\,
            lcout => \POWERLED.func_m1_0_a2Z0Z_0\,
            ltout => \POWERLED.func_m1_0_a2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPUCL3_0_1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__20353\,
            in1 => \_gnd_net_\,
            in2 => \N__20380\,
            in3 => \N__20377\,
            lcout => \POWERLED.N_433\,
            ltout => \POWERLED.N_433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2K64A_1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011011111"
        )
    port map (
            in0 => \N__20641\,
            in1 => \N__20627\,
            in2 => \N__20371\,
            in3 => \N__20368\,
            lcout => \POWERLED.func_state_1_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIIN481_1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__23661\,
            in1 => \N__20318\,
            in2 => \N__24560\,
            in3 => \N__24326\,
            lcout => \POWERLED.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_m1_0_a2_0_iso_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__24253\,
            in2 => \N__20331\,
            in3 => \N__23659\,
            lcout => \POWERLED.func_m1_0_a2_0_isoZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIIN481_0_1_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23660\,
            in1 => \N__20317\,
            in2 => \N__24559\,
            in3 => \N__24325\,
            lcout => OPEN,
            ltout => \POWERLED.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPUCL3_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30093\,
            in1 => \N__20662\,
            in2 => \N__20650\,
            in3 => \N__20647\,
            lcout => \POWERLED.N_79\,
            ltout => \POWERLED.N_79_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNINROUB_0_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001001111"
        )
    port map (
            in0 => \N__20628\,
            in1 => \N__20614\,
            in2 => \N__20608\,
            in3 => \N__20605\,
            lcout => \POWERLED.func_state_1_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__35994\,
            in1 => \N__26969\,
            in2 => \_gnd_net_\,
            in3 => \N__22219\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIH0LB7_0_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__29932\,
            in2 => \N__20566\,
            in3 => \N__20724\,
            lcout => \POWERLED.dutycycle_RNIH0LB7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI0TA81_0_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001111"
        )
    port map (
            in0 => \N__20725\,
            in1 => \N__26970\,
            in2 => \N__31828\,
            in3 => \N__22220\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3F2B2_1_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35995\,
            in2 => \N__20422\,
            in3 => \N__24619\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPHPH3_1_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22324\,
            in2 => \N__20419\,
            in3 => \N__27932\,
            lcout => \POWERLED.N_189_i\,
            ltout => \POWERLED.N_189_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIML1B1_1_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110001"
        )
    port map (
            in0 => \N__27933\,
            in1 => \N__22477\,
            in2 => \N__20404\,
            in3 => \N__24420\,
            lcout => \POWERLED.N_122_f0_1\,
            ltout => \POWERLED.N_122_f0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNID9PI3_0_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__30092\,
            in1 => \N__27934\,
            in2 => \N__20686\,
            in3 => \N__35657\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNID9PI3_1_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110010"
        )
    port map (
            in0 => \N__27935\,
            in1 => \N__20683\,
            in2 => \N__30133\,
            in3 => \N__32097\,
            lcout => \POWERLED.dutycycle_eena_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_1_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__27051\,
            in1 => \N__32073\,
            in2 => \_gnd_net_\,
            in3 => \N__22203\,
            lcout => OPEN,
            ltout => \POWERLED.g0_i_a6_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__36757\,
            in1 => \N__35656\,
            in2 => \N__20677\,
            in3 => \N__30241\,
            lcout => \POWERLED.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__30242\,
            in1 => \N__32074\,
            in2 => \N__29383\,
            in3 => \N__36702\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_rep1_RNI_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30240\,
            lcout => \tmp_1_rep1_RNI\,
            ltout => \tmp_1_rep1_RNI_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_0_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__36756\,
            in1 => \N__35655\,
            in2 => \N__20668\,
            in3 => \N__32072\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_6_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27185\,
            in1 => \N__27053\,
            in2 => \N__36789\,
            in3 => \N__30243\,
            lcout => \POWERLED.N_358\,
            ltout => \POWERLED.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__20866\,
            in1 => \N__20726\,
            in2 => \N__20665\,
            in3 => \N__22202\,
            lcout => \POWERLED.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__30250\,
            in1 => \N__24511\,
            in2 => \_gnd_net_\,
            in3 => \N__27052\,
            lcout => \POWERLED.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22212\,
            in1 => \N__20862\,
            in2 => \_gnd_net_\,
            in3 => \N__20719\,
            lcout => \POWERLED.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_1_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__22443\,
            in1 => \N__24562\,
            in2 => \N__22640\,
            in3 => \N__22669\,
            lcout => \POWERLED.g0_i_a6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__32672\,
            in1 => \_gnd_net_\,
            in2 => \N__27139\,
            in3 => \N__37141\,
            lcout => \POWERLED.N_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__20740\,
            in1 => \N__20873\,
            in2 => \N__20728\,
            in3 => \N__27135\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_42_and_i_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3IN21_2_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__31818\,
            in1 => \N__32941\,
            in2 => \N__20734\,
            in3 => \N__29336\,
            lcout => OPEN,
            ltout => \POWERLED.N_434_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGV14_12_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011111111"
        )
    port map (
            in0 => \N__37142\,
            in1 => \N__32671\,
            in2 => \N__20731\,
            in3 => \N__27248\,
            lcout => \POWERLED.N_235_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_2_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32163\,
            in3 => \N__29335\,
            lcout => \POWERLED.N_372\,
            ltout => \POWERLED.N_372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_0_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20720\,
            in1 => \N__22575\,
            in2 => \N__20689\,
            in3 => \N__20872\,
            lcout => \POWERLED.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0TA81_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__24577\,
            in1 => \N__20888\,
            in2 => \N__35683\,
            in3 => \N__26978\,
            lcout => \POWERLED.dutycycle_1_0_0\,
            ltout => \POWERLED.dutycycle_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITOAI5_0_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__20925\,
            in1 => \N__20940\,
            in2 => \N__20950\,
            in3 => \N__29956\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__20926\,
            in1 => \N__20947\,
            in2 => \N__29970\,
            in3 => \N__20941\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \N__32476\
        );

    \POWERLED.dutycycle_1_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__20809\,
            in1 => \N__20788\,
            in2 => \N__20803\,
            in3 => \N__29961\,
            lcout => \POWERLED.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \N__32476\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001101"
        )
    port map (
            in0 => \N__24576\,
            in1 => \N__26977\,
            in2 => \N__22951\,
            in3 => \N__20887\,
            lcout => \POWERLED.dutycycle_1_0_1\,
            ltout => \POWERLED.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI149J5_1_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__20802\,
            in1 => \N__20787\,
            in2 => \N__20779\,
            in3 => \N__29957\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__23065\,
            in1 => \N__29963\,
            in2 => \N__20776\,
            in3 => \N__20767\,
            lcout => \POWERLED.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \N__32440\
        );

    \POWERLED.dutycycle_RNI778D2_11_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__32952\,
            in1 => \N__32651\,
            in2 => \N__30175\,
            in3 => \N__30021\,
            lcout => \POWERLED.dutycycle_eena_7\,
            ltout => \POWERLED.dutycycle_eena_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI01PN4_11_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__23064\,
            in1 => \N__20766\,
            in2 => \N__20758\,
            in3 => \N__29962\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => \POWERLED.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20755\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_11\,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_11_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31945\,
            in2 => \N__21001\,
            in3 => \N__37144\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__37227\,
            in1 => \N__36438\,
            in2 => \N__20998\,
            in3 => \N__37146\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_12_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20995\,
            in3 => \N__20992\,
            lcout => \POWERLED.un1_dutycycle_53_axb_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011011111110"
        )
    port map (
            in0 => \N__37143\,
            in1 => \N__36437\,
            in2 => \N__37261\,
            in3 => \N__32194\,
            lcout => \POWERLED.un1_dutycycle_53_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21804\,
            lcout => \N_414\,
            ltout => \N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20968\,
            in2 => \N__20986\,
            in3 => \N__34198\,
            lcout => \HDA_STRAP.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34990\,
            ce => \N__30949\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010011101"
        )
    port map (
            in0 => \N__21172\,
            in1 => \N__21821\,
            in2 => \N__20983\,
            in3 => \N__21117\,
            lcout => \HDA_STRAP.m6_i_0\,
            ltout => \HDA_STRAP.m6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m6_i_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34196\,
            in2 => \N__20962\,
            in3 => \N__22061\,
            lcout => OPEN,
            ltout => \HDA_STRAP.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNITJDR4_0_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20959\,
            in2 => \N__20953\,
            in3 => \N__23665\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34197\,
            in2 => \_gnd_net_\,
            in3 => \N__22062\,
            lcout => \HDA_STRAP.N_285\,
            ltout => \HDA_STRAP.N_285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m8_i_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__21174\,
            in1 => \N__21822\,
            in2 => \N__21151\,
            in3 => \N__21116\,
            lcout => \HDA_STRAP.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNI9A8D5_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__21577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21121\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21133\,
            in2 => \_gnd_net_\,
            in3 => \N__27991\,
            lcout => \N_227\,
            ltout => \N_227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_0_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21094\,
            in3 => \_gnd_net_\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21063\,
            in1 => \N__21051\,
            in2 => \N__21040\,
            in3 => \N__21024\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__21013\,
            in1 => \N__21422\,
            in2 => \_gnd_net_\,
            in3 => \N__22031\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22028\,
            in1 => \N__21405\,
            in2 => \_gnd_net_\,
            in3 => \N__21564\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__21007\,
            in1 => \N__21343\,
            in2 => \_gnd_net_\,
            in3 => \N__22029\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21489\,
            in1 => \N__21477\,
            in2 => \N__21466\,
            in3 => \N__21450\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21438\,
            in1 => \N__21383\,
            in2 => \N__21426\,
            in3 => \N__21404\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__21384\,
            in1 => \N__21391\,
            in2 => \_gnd_net_\,
            in3 => \N__22030\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22023\,
            in1 => \N__21370\,
            in2 => \_gnd_net_\,
            in3 => \N__21357\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21356\,
            in1 => \N__21341\,
            in2 => \N__21210\,
            in3 => \N__21559\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21324\,
            in1 => \N__21312\,
            in2 => \N__21301\,
            in3 => \N__21285\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21273\,
            in1 => \N__21261\,
            in2 => \N__21250\,
            in3 => \N__21234\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__21206\,
            in1 => \N__21223\,
            in2 => \_gnd_net_\,
            in3 => \N__22027\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__21560\,
            in1 => \_gnd_net_\,
            in2 => \N__22033\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIBCB91_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23292\,
            in1 => \N__23238\,
            in2 => \N__23326\,
            in3 => \N__23277\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.un4_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIB8TE4_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21538\,
            in1 => \N__25258\,
            in2 => \N__21541\,
            in3 => \N__21532\,
            lcout => \DSW_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIH71P_2_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23160\,
            in1 => \N__23190\,
            in2 => \N__23209\,
            in3 => \N__23340\,
            lcout => \DSW_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIKA1P_1_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23355\,
            in1 => \N__23175\,
            in2 => \N__23227\,
            in3 => \N__23307\,
            lcout => \DSW_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21517\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21508\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21499\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21610\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21601\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21592\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21586\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER.un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_THRU_LUT4_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21580\,
            lcout => \COUNTER.un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__31004\,
            in1 => \N__23399\,
            in2 => \N__21640\,
            in3 => \N__21709\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__23553\,
            in1 => \N__26818\,
            in2 => \_gnd_net_\,
            in3 => \N__25858\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21686\,
            in1 => \N__23414\,
            in2 => \N__21655\,
            in3 => \N__23552\,
            lcout => \VPP_VDDQ.count_2_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23433\,
            in1 => \N__21651\,
            in2 => \_gnd_net_\,
            in3 => \N__21685\,
            lcout => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__31003\,
            in1 => \N__21708\,
            in2 => \N__21712\,
            in3 => \N__21636\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__23415\,
            in1 => \N__21684\,
            in2 => \_gnd_net_\,
            in3 => \N__21650\,
            lcout => \VPP_VDDQ.N_297_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIHU1M_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26819\,
            in1 => \N__23554\,
            in2 => \N__25870\,
            in3 => \N__31001\,
            lcout => \POWERLED.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26600\,
            in1 => \N__26529\,
            in2 => \N__26572\,
            in3 => \N__26633\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_15_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26456\,
            in2 => \N__21625\,
            in3 => \N__26489\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_8_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26201\,
            in1 => \N__26156\,
            in2 => \N__21622\,
            in3 => \N__21616\,
            lcout => \POWERLED.count_RNIZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_2_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25935\,
            in1 => \N__26358\,
            in2 => \_gnd_net_\,
            in3 => \N__26403\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_5_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__26283\,
            in1 => \N__26240\,
            in2 => \N__21619\,
            in3 => \N__26315\,
            lcout => \POWERLED.un79_clk_100khzlto15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI5S8O_15_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21772\,
            in1 => \N__23644\,
            in2 => \_gnd_net_\,
            in3 => \N__21780\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21784\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35177\,
            ce => \N__30952\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI7UKN_7_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21766\,
            in1 => \N__21757\,
            in2 => \_gnd_net_\,
            in3 => \N__23645\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21765\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35177\,
            ce => \N__30952\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI91MN_8_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21751\,
            in1 => \N__21742\,
            in2 => \_gnd_net_\,
            in3 => \N__23646\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21750\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35177\,
            ce => \N__30952\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIB4NN_9_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21724\,
            in1 => \N__23647\,
            in2 => \_gnd_net_\,
            in3 => \N__21735\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21736\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35177\,
            ce => \N__30952\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHU7V2_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110101"
        )
    port map (
            in0 => \N__24090\,
            in1 => \N__24232\,
            in2 => \N__24157\,
            in3 => \N__21718\,
            lcout => \POWERLED.func_state_RNIHU7V2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_0_o3_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101111111111"
        )
    port map (
            in0 => \N__22089\,
            in1 => \N__21843\,
            in2 => \N__24247\,
            in3 => \N__22474\,
            lcout => \VCCST_EN_i_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_fast_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__24152\,
            in1 => \N__22022\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SUSWARN_N_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_rep1_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__22090\,
            in1 => \_gnd_net_\,
            in2 => \N__22032\,
            in3 => \_gnd_net_\,
            lcout => \SUSWARN_N_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_rep1_RNI2PKG_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22088\,
            in2 => \_gnd_net_\,
            in3 => \N__22017\,
            lcout => \VPP_VDDQ_delayed_vddq_pwrgd_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_en_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22063\,
            in2 => \_gnd_net_\,
            in3 => \N__30998\,
            lcout => \HDA_STRAP.count_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNIBJDJ_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23658\,
            in2 => \_gnd_net_\,
            in3 => \N__22018\,
            lcout => \un4_counter_7_c_RNIBJDJ\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25152\,
            lcout => v1p8a_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21958\,
            in1 => \N__28043\,
            in2 => \_gnd_net_\,
            in3 => \N__21910\,
            lcout => \RSMRSTn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35277\,
            ce => \N__30955\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNI_1_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21829\,
            lcout => \HDA_STRAP.N_2989_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29168\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNII69M3_5_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__29933\,
            in1 => \N__22176\,
            in2 => \N__22129\,
            in3 => \N__30070\,
            lcout => \POWERLED.dutycycle_RNII69M3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_rep1_RNILDD26_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__22177\,
            in1 => \N__22786\,
            in2 => \_gnd_net_\,
            in3 => \N__29934\,
            lcout => \COUNTER.N_96_mux_i_i_a8_1\,
            ltout => \COUNTER.N_96_mux_i_i_a8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_rep1_RNIC08FV_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__26749\,
            in1 => \N__22144\,
            in2 => \N__22162\,
            in3 => \N__26736\,
            lcout => \tmp_1_rep1_RNIC08FV_0\,
            ltout => \tmp_1_rep1_RNIC08FV_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_6_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__26901\,
            in1 => \_gnd_net_\,
            in2 => \N__22159\,
            in3 => \N__31906\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_6Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2T1A8_5_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__22156\,
            in1 => \N__22114\,
            in2 => \N__22147\,
            in3 => \N__26884\,
            lcout => \N_96_mux_i_i_3\,
            ltout => \N_96_mux_i_i_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__26737\,
            in1 => \N__26748\,
            in2 => \N__22138\,
            in3 => \N__22135\,
            lcout => \POWERLED.dutycycleZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35001\,
            ce => 'H',
            sr => \N__32390\
        );

    \POWERLED.dutycycle_RNIAI9E2_5_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30069\,
            in2 => \N__22128\,
            in3 => \N__27967\,
            lcout => \POWERLED.N_31\,
            ltout => \POWERLED.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIAI9E2_0_5_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000001111"
        )
    port map (
            in0 => \N__26900\,
            in1 => \_gnd_net_\,
            in2 => \N__22672\,
            in3 => \N__31905\,
            lcout => \POWERLED.N_96_mux_i_i_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001011"
        )
    port map (
            in0 => \N__36133\,
            in1 => \N__36037\,
            in2 => \N__32005\,
            in3 => \N__31827\,
            lcout => \POWERLED.g2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI34G9_6_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36132\,
            lcout => \POWERLED.g0_i_a6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_2_1_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__22663\,
            in1 => \N__22460\,
            in2 => \N__22605\,
            in3 => \N__22323\,
            lcout => \POWERLED.un1_clk_100khz_52_and_i_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_1_1_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__22565\,
            in2 => \N__22331\,
            in3 => \N__24575\,
            lcout => OPEN,
            ltout => \POWERLED.N_387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDUQ02_1_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__36134\,
            in1 => \N__22461\,
            in2 => \N__22645\,
            in3 => \N__22625\,
            lcout => \POWERLED.func_state_RNIDUQ02Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__22458\,
            in1 => \N__22564\,
            in2 => \_gnd_net_\,
            in3 => \N__24574\,
            lcout => \POWERLED.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_0_0_6_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__22563\,
            in1 => \N__22457\,
            in2 => \_gnd_net_\,
            in3 => \N__22319\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_6_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27184\,
            in1 => \N__30239\,
            in2 => \N__22221\,
            in3 => \N__36755\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7T3_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__36030\,
            in1 => \N__22909\,
            in2 => \N__30171\,
            in3 => \N__22830\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7TZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILF063_6_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110000"
        )
    port map (
            in0 => \N__22876\,
            in1 => \N__36028\,
            in2 => \N__22772\,
            in3 => \N__36787\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_m2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM6QF4_6_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101101010"
        )
    port map (
            in0 => \N__36788\,
            in1 => \N__24290\,
            in2 => \N__22870\,
            in3 => \N__24812\,
            lcout => OPEN,
            ltout => \POWERLED.N_233_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQOL27_6_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__24586\,
            in1 => \N__30146\,
            in2 => \N__22867\,
            in3 => \N__22864\,
            lcout => \POWERLED.dutycycle_eena_13\,
            ltout => \POWERLED.dutycycle_eena_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBE4NB_6_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__22855\,
            in1 => \N__22839\,
            in2 => \N__22858\,
            in3 => \N__29911\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__22840\,
            in1 => \N__22854\,
            in2 => \N__29955\,
            in3 => \N__22846\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35243\,
            ce => 'H',
            sr => \N__32472\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIQQ6T3_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__36029\,
            in1 => \N__22918\,
            in2 => \N__30170\,
            in3 => \N__22829\,
            lcout => \POWERLED_dutycycle_set_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__24289\,
            in1 => \N__36027\,
            in2 => \N__22773\,
            in3 => \N__22744\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_337_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_0_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35654\,
            in3 => \N__32067\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32068\,
            in2 => \N__23043\,
            in3 => \N__22942\,
            lcout => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29369\,
            in2 => \N__23024\,
            in3 => \N__22927\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22995\,
            in2 => \N__37004\,
            in3 => \N__22924\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36701\,
            in2 => \N__23025\,
            in3 => \N__22921\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32908\,
            in1 => \N__22999\,
            in2 => \N__30272\,
            in3 => \N__22912\,
            lcout => \POWERLED.N_308\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIB6R31_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32940\,
            in1 => \N__36786\,
            in2 => \N__23026\,
            in3 => \N__22903\,
            lcout => \POWERLED.N_307\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37510\,
            in2 => \N__23042\,
            in3 => \N__22885\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37335\,
            in2 => \N__23047\,
            in3 => \N__22882\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\,
            ltout => OPEN,
            carryin => \bfn_6_16_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23041\,
            in2 => \N__37251\,
            in3 => \N__22879\,
            lcout => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36419\,
            in2 => \N__23046\,
            in3 => \N__23068\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32919\,
            in1 => \N__23027\,
            in2 => \N__31980\,
            in3 => \N__23056\,
            lcout => \POWERLED.dutycycle_rst_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32953\,
            in1 => \N__37121\,
            in2 => \N__23044\,
            in3 => \N__23053\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23031\,
            in2 => \N__32749\,
            in3 => \N__23050\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32323\,
            in2 => \N__23045\,
            in3 => \N__22963\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__30395\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__22960\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_6_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25048\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34586\,
            ce => \N__27559\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI7AQ41_2_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24831\,
            in1 => \N__22957\,
            in2 => \_gnd_net_\,
            in3 => \N__27526\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24832\,
            lcout => \VPP_VDDQ.count_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34586\,
            ce => \N__27559\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFMU41_6_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23098\,
            in1 => \N__27529\,
            in2 => \_gnd_net_\,
            in3 => \N__25047\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => \VPP_VDDQ.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_10_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24921\,
            in1 => \N__25371\,
            in2 => \N__23092\,
            in3 => \N__24844\,
            lcout => \VPP_VDDQ.un13_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIUHA31_10_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24907\,
            in1 => \N__23089\,
            in2 => \_gnd_net_\,
            in3 => \N__27527\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_10_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24906\,
            lcout => \VPP_VDDQ.count_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34586\,
            ce => \N__27559\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI95OO_12_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__27325\,
            in2 => \_gnd_net_\,
            in3 => \N__27528\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_0_c_RNO_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__24993\,
            in1 => \N__23132\,
            in2 => \N__27525\,
            in3 => \N__23122\,
            lcout => \VPP_VDDQ.un4_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_0_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24992\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI513Q_0_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23121\,
            in2 => \N__23083\,
            in3 => \N__27484\,
            lcout => \VPP_VDDQ.N_3013_i\,
            ltout => \VPP_VDDQ.N_3013_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_15_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27577\,
            in1 => \N__27415\,
            in2 => \N__23080\,
            in3 => \N__25344\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un13_clk_100khz_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_0_10_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__23077\,
            in1 => \N__24715\,
            in2 => \N__23146\,
            in3 => \N__23245\,
            lcout => \VPP_VDDQ.count_RNI_1_10\,
            ltout => \VPP_VDDQ.count_RNI_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI72NO_11_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__25384\,
            in1 => \N__23140\,
            in2 => \N__23143\,
            in3 => \N__27489\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_11_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25383\,
            lcout => \VPP_VDDQ.count_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34812\,
            ce => \N__27488\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24995\,
            lcout => \VPP_VDDQ.count_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34812\,
            ce => \N__27488\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_8_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25014\,
            lcout => \VPP_VDDQ.count_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => \N__27519\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNILV151_9_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__24934\,
            in2 => \_gnd_net_\,
            in3 => \N__27521\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_1_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24856\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => \N__27519\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI2PKG_1_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31046\,
            in2 => \_gnd_net_\,
            in3 => \N__29943\,
            lcout => \VPP_VDDQ.count_en\,
            ltout => \VPP_VDDQ.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI57P41_1_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24855\,
            in2 => \N__23113\,
            in3 => \N__23110\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_9_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24933\,
            lcout => \VPP_VDDQ.count_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => \N__27519\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIJS051_8_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27520\,
            in1 => \N__23254\,
            in2 => \_gnd_net_\,
            in3 => \N__25015\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => \VPP_VDDQ.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_11_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24945\,
            in1 => \N__25395\,
            in2 => \N__23248\,
            in3 => \N__24868\,
            lcout => \VPP_VDDQ.un13_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27844\,
            in1 => \N__23239\,
            in2 => \N__25438\,
            in3 => \N__25437\,
            lcout => \DSW_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_0\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27840\,
            in1 => \N__23226\,
            in2 => \_gnd_net_\,
            in3 => \N__23212\,
            lcout => \DSW_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_0\,
            carryout => \DSW_PWRGD.un1_count_1_cry_1\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_2_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27845\,
            in1 => \N__23208\,
            in2 => \_gnd_net_\,
            in3 => \N__23194\,
            lcout => \DSW_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_1\,
            carryout => \DSW_PWRGD.un1_count_1_cry_2\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_3_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27841\,
            in1 => \N__23191\,
            in2 => \_gnd_net_\,
            in3 => \N__23179\,
            lcout => \DSW_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_2\,
            carryout => \DSW_PWRGD.un1_count_1_cry_3\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_4_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27846\,
            in1 => \N__23176\,
            in2 => \_gnd_net_\,
            in3 => \N__23164\,
            lcout => \DSW_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_3\,
            carryout => \DSW_PWRGD.un1_count_1_cry_4\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_5_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27842\,
            in1 => \N__23161\,
            in2 => \_gnd_net_\,
            in3 => \N__23149\,
            lcout => \DSW_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_4\,
            carryout => \DSW_PWRGD.un1_count_1_cry_5\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_6_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27847\,
            in1 => \N__23356\,
            in2 => \_gnd_net_\,
            in3 => \N__23344\,
            lcout => \DSW_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_5\,
            carryout => \DSW_PWRGD.un1_count_1_cry_6\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_7_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27843\,
            in1 => \N__23341\,
            in2 => \_gnd_net_\,
            in3 => \N__23329\,
            lcout => \DSW_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_6\,
            carryout => \DSW_PWRGD.un1_count_1_cry_7\,
            clk => \N__34819\,
            ce => 'H',
            sr => \N__27744\
        );

    \DSW_PWRGD.count_8_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27839\,
            in1 => \N__23325\,
            in2 => \_gnd_net_\,
            in3 => \N__23311\,
            lcout => \DSW_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_8\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.count_9_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27835\,
            in1 => \N__23308\,
            in2 => \_gnd_net_\,
            in3 => \N__23296\,
            lcout => \DSW_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_8\,
            carryout => \DSW_PWRGD.un1_count_1_cry_9\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.count_10_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27836\,
            in1 => \N__23293\,
            in2 => \_gnd_net_\,
            in3 => \N__23281\,
            lcout => \DSW_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_9\,
            carryout => \DSW_PWRGD.un1_count_1_cry_10\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.count_11_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27833\,
            in1 => \N__23278\,
            in2 => \_gnd_net_\,
            in3 => \N__23266\,
            lcout => \DSW_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_10\,
            carryout => \DSW_PWRGD.un1_count_1_cry_11\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.count_12_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27837\,
            in1 => \N__25270\,
            in2 => \_gnd_net_\,
            in3 => \N__23263\,
            lcout => \DSW_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_11\,
            carryout => \DSW_PWRGD.un1_count_1_cry_12\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.count_13_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27834\,
            in1 => \N__25309\,
            in2 => \_gnd_net_\,
            in3 => \N__23260\,
            lcout => \DSW_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_12\,
            carryout => \DSW_PWRGD.un1_count_1_cry_13\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.count_14_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27838\,
            in1 => \N__25284\,
            in2 => \_gnd_net_\,
            in3 => \N__23257\,
            lcout => \DSW_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_13\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14\,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__27737\
        );

    \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31666\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_14\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_15_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25297\,
            in2 => \_gnd_net_\,
            in3 => \N__23770\,
            lcout => \DSW_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34820\,
            ce => \N__25786\,
            sr => \N__27745\
        );

    \VPP_VDDQ.curr_state_2_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__23758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27642\,
            lcout => \VPP_VDDQ.curr_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34821\,
            ce => \N__30943\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__23686\,
            in1 => \N__23757\,
            in2 => \N__27646\,
            in3 => \N__23767\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23761\,
            in3 => \N__33074\,
            lcout => \VPP_VDDQ.m4_0_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__23379\,
            in1 => \N__23401\,
            in2 => \N__33079\,
            in3 => \N__23416\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23362\,
            in2 => \N__23749\,
            in3 => \N__23685\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23419\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_2877_i\,
            ltout => \VPP_VDDQ.N_2877_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__23400\,
            in1 => \N__33075\,
            in2 => \N__23386\,
            in3 => \N__23378\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34821\,
            ce => \N__30943\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29431\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23806\,
            in2 => \N__26080\,
            in3 => \N__23794\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23941\,
            in2 => \N__23956\,
            in3 => \N__23791\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23928\,
            in2 => \N__23860\,
            in3 => \N__23788\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23848\,
            in2 => \N__23932\,
            in3 => \N__23785\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__26059\,
            in1 => \N__23776\,
            in2 => \N__23839\,
            in3 => \N__23782\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23779\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23927\,
            in2 => \_gnd_net_\,
            in3 => \N__23835\,
            lcout => \POWERLED.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29302\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26431\,
            in2 => \N__26097\,
            in3 => \N__23863\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26093\,
            in2 => \N__23902\,
            in3 => \N__23851\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23887\,
            in2 => \N__26132\,
            in3 => \N__23842\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26126\,
            in2 => \N__23875\,
            in3 => \N__23824\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23924\,
            in1 => \N__24061\,
            in2 => \N__26098\,
            in3 => \N__23815\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24049\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23812\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => \POWERLED.mult1_un124_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23809\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFERO_15_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27561\,
            in1 => \N__23800\,
            in2 => \_gnd_net_\,
            in3 => \N__25323\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_15_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35131\,
            ce => \N__27560\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_6_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31819\,
            lcout => \POWERLED.N_203_i\,
            ltout => \POWERLED.N_203_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23989\,
            in3 => \N__36031\,
            lcout => \POWERLED.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0TA81_0_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26976\,
            in2 => \_gnd_net_\,
            in3 => \N__27056\,
            lcout => \POWERLED.func_state_RNI0TA81_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23926\,
            lcout => \POWERLED.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29248\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24029\,
            in2 => \N__24355\,
            in3 => \N__23890\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24019\,
            in2 => \N__24034\,
            in3 => \N__23878\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26709\,
            in2 => \N__24010\,
            in3 => \N__24064\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23998\,
            in2 => \N__26713\,
            in3 => \N__24052\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__26114\,
            in1 => \N__24033\,
            in2 => \N__24394\,
            in3 => \N__24040\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24037\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26708\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29211\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24377\,
            in2 => \N__26725\,
            in3 => \N__24013\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28687\,
            in2 => \N__24382\,
            in3 => \N__24001\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29169\,
            in2 => \N__28672\,
            in3 => \N__23992\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28654\,
            in2 => \N__29173\,
            in3 => \N__24385\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__26706\,
            in1 => \N__24381\,
            in2 => \N__28639\,
            in3 => \N__24361\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24358\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29212\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3IN21_0_2_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__24248\,
            in1 => \N__24145\,
            in2 => \N__24346\,
            in3 => \N__24094\,
            lcout => \POWERLED.g1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__24166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36131\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_36_and_i_a2_1_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_2_1_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__24250\,
            in1 => \N__24144\,
            in2 => \N__24334\,
            in3 => \N__24093\,
            lcout => \POWERLED.N_332_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24092\,
            in1 => \N__24143\,
            in2 => \_gnd_net_\,
            in3 => \N__24251\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_0_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__24249\,
            in1 => \N__24165\,
            in2 => \N__24155\,
            in3 => \N__24091\,
            lcout => \POWERLED.func_state_RNI3IN21_0Z0Z_1\,
            ltout => \POWERLED.func_state_RNI3IN21_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI64F52_0_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__24661\,
            in2 => \N__24655\,
            in3 => \N__27070\,
            lcout => \POWERLED.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__32179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32122\,
            lcout => \POWERLED.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31594\,
            lcout => \POWERLED.mult1_un96_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32854\,
            in1 => \N__24633\,
            in2 => \N__24652\,
            in3 => \N__27286\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35242\,
            ce => 'H',
            sr => \N__32459\
        );

    \POWERLED.dutycycle_RNIN84N7_14_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__27285\,
            in1 => \N__24648\,
            in2 => \N__24634\,
            in3 => \N__32853\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_15_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__30387\,
            in1 => \_gnd_net_\,
            in2 => \N__24622\,
            in3 => \N__32607\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3IN21_6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__26935\,
            in1 => \N__26671\,
            in2 => \_gnd_net_\,
            in3 => \N__24599\,
            lcout => \POWERLED.dutycycle_RNI3IN21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIU6GQ_1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__24600\,
            in1 => \N__27055\,
            in2 => \N__31168\,
            in3 => \N__24563\,
            lcout => \POWERLED.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27054\,
            in2 => \_gnd_net_\,
            in3 => \N__24561\,
            lcout => \POWERLED.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQU4T5_4_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__32503\,
            in2 => \N__27256\,
            in3 => \N__24700\,
            lcout => \POWERLED.dutycycle_en_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI554R1_8_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110011"
        )
    port map (
            in0 => \N__24709\,
            in1 => \N__24676\,
            in2 => \N__32938\,
            in3 => \N__29949\,
            lcout => \POWERLED.dutycycle_RNI554R1Z0Z_8\,
            ltout => \POWERLED.dutycycle_RNI554R1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJC6E7_8_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000001111"
        )
    port map (
            in0 => \N__30153\,
            in1 => \N__24674\,
            in2 => \N__24703\,
            in3 => \N__24691\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI778D2_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__32901\,
            in1 => \N__30154\,
            in2 => \N__32542\,
            in3 => \N__36160\,
            lcout => \POWERLED.func_state_RNI778D2Z0Z_1\,
            ltout => \POWERLED.func_state_RNI778D2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQU4T5_3_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__27245\,
            in1 => \N__29942\,
            in2 => \N__24694\,
            in3 => \N__31606\,
            lcout => \POWERLED.dutycycle_RNIQU4T5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGV14_8_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101011111"
        )
    port map (
            in0 => \N__32541\,
            in1 => \N__37336\,
            in2 => \N__24820\,
            in3 => \N__27241\,
            lcout => \POWERLED.dutycycle_RNIKGV14Z0Z_8\,
            ltout => \POWERLED.dutycycle_RNIKGV14Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011101111"
        )
    port map (
            in0 => \N__30155\,
            in1 => \N__24675\,
            in2 => \N__24685\,
            in3 => \N__24682\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35152\,
            ce => 'H',
            sr => \N__32431\
        );

    \POWERLED.dutycycle_4_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__29580\,
            in1 => \N__29559\,
            in2 => \N__32939\,
            in3 => \N__29544\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35152\,
            ce => 'H',
            sr => \N__32431\
        );

    \POWERLED.dutycycle_9_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__24793\,
            in1 => \N__24759\,
            in2 => \N__24784\,
            in3 => \N__30174\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35311\,
            ce => 'H',
            sr => \N__32471\
        );

    \POWERLED.dutycycle_RNIKGV14_9_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101111"
        )
    port map (
            in0 => \N__29739\,
            in1 => \N__37207\,
            in2 => \N__24819\,
            in3 => \N__27246\,
            lcout => \POWERLED.N_116_f0\,
            ltout => \POWERLED.N_116_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMG7E7_9_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__24779\,
            in1 => \N__24760\,
            in2 => \N__24787\,
            in3 => \N__30173\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI785R1_9_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32890\,
            in1 => \N__24780\,
            in2 => \N__24769\,
            in3 => \N__29950\,
            lcout => \POWERLED.dutycycle_e_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8BF97_10_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__24738\,
            in1 => \N__24745\,
            in2 => \N__24727\,
            in3 => \N__32889\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => \POWERLED.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGV14_10_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__32891\,
            in1 => \N__27247\,
            in2 => \N__24751\,
            in3 => \N__36161\,
            lcout => OPEN,
            ltout => \POWERLED.N_157_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQU4T5_10_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__29732\,
            in1 => \N__29947\,
            in2 => \N__24748\,
            in3 => \N__30172\,
            lcout => \POWERLED.dutycycle_en_4\,
            ltout => \POWERLED.dutycycle_en_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__32892\,
            in1 => \N__24739\,
            in2 => \N__24730\,
            in3 => \N__24726\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35311\,
            ce => 'H',
            sr => \N__32471\
        );

    \VPP_VDDQ.count_RNI_3_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25078\,
            in1 => \N__25036\,
            in2 => \N__25129\,
            in3 => \N__25102\,
            lcout => \VPP_VDDQ.un13_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI9DR41_3_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24892\,
            in1 => \N__27530\,
            in2 => \_gnd_net_\,
            in3 => \N__25113\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34597\,
            ce => \N__27558\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIBGS41_4_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24886\,
            in1 => \N__27531\,
            in2 => \_gnd_net_\,
            in3 => \N__25089\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_4_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34597\,
            ce => \N__27558\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIDJT41_5_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25065\,
            in1 => \N__24880\,
            in2 => \_gnd_net_\,
            in3 => \N__27532\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_5_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25066\,
            lcout => \VPP_VDDQ.count_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34597\,
            ce => \N__27558\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIHPV41_7_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27304\,
            in1 => \N__27533\,
            in2 => \_gnd_net_\,
            in3 => \N__27316\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_0_c_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24874\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \VPP_VDDQ.un4_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_0_c_RNIV4MA_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24867\,
            in2 => \_gnd_net_\,
            in3 => \N__24847\,
            lcout => \VPP_VDDQ.count_rst_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24843\,
            in2 => \_gnd_net_\,
            in3 => \N__24823\,
            lcout => \VPP_VDDQ.count_rst_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_1\,
            carryout => \VPP_VDDQ.un4_count_1_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__24996\,
            in1 => \N__25125\,
            in2 => \_gnd_net_\,
            in3 => \N__25105\,
            lcout => \VPP_VDDQ.count_rst_8\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_2_cZ0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__24999\,
            in1 => \N__25101\,
            in2 => \_gnd_net_\,
            in3 => \N__25081\,
            lcout => \VPP_VDDQ.count_rst_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_3_cZ0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__24997\,
            in1 => \N__25077\,
            in2 => \_gnd_net_\,
            in3 => \N__25057\,
            lcout => \VPP_VDDQ.count_rst_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_4_cZ0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25054\,
            in2 => \_gnd_net_\,
            in3 => \N__25039\,
            lcout => \VPP_VDDQ.count_rst_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_5\,
            carryout => \VPP_VDDQ.un4_count_1_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__24998\,
            in1 => \N__25035\,
            in2 => \_gnd_net_\,
            in3 => \N__25024\,
            lcout => \VPP_VDDQ.count_rst_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_6_cZ0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25001\,
            in1 => \N__25021\,
            in2 => \_gnd_net_\,
            in3 => \N__25006\,
            lcout => \VPP_VDDQ.count_rst_13\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \VPP_VDDQ.un4_count_1_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25000\,
            in1 => \N__24946\,
            in2 => \_gnd_net_\,
            in3 => \N__24925\,
            lcout => \VPP_VDDQ.count_rst_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_8_cZ0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24922\,
            in2 => \_gnd_net_\,
            in3 => \N__24895\,
            lcout => \VPP_VDDQ.count_rst\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_9\,
            carryout => \VPP_VDDQ.un4_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6C_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25396\,
            in2 => \_gnd_net_\,
            in3 => \N__25375\,
            lcout => \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6CZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_10\,
            carryout => \VPP_VDDQ.un4_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25372\,
            in2 => \_gnd_net_\,
            in3 => \N__25357\,
            lcout => \VPP_VDDQ.count_rst_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_11\,
            carryout => \VPP_VDDQ.un4_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27573\,
            in2 => \_gnd_net_\,
            in3 => \N__25354\,
            lcout => \VPP_VDDQ.count_rst_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_12\,
            carryout => \VPP_VDDQ.un4_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27414\,
            in3 => \N__25351\,
            lcout => \VPP_VDDQ.count_rst_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_13\,
            carryout => \VPP_VDDQ.un4_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25348\,
            in2 => \_gnd_net_\,
            in3 => \N__25327\,
            lcout => \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25308\,
            in1 => \N__25296\,
            in2 => \N__25285\,
            in3 => \N__25269\,
            lcout => \DSW_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNILLF15_0_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__28175\,
            in1 => \N__28206\,
            in2 => \N__25462\,
            in3 => \N__28152\,
            lcout => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25232\,
            in1 => \N__25204\,
            in2 => \N__25195\,
            in3 => \N__25156\,
            lcout => \N_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_7_1_0__m3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25460\,
            in1 => \N__28203\,
            in2 => \_gnd_net_\,
            in3 => \N__28153\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.i3_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010101010"
        )
    port map (
            in0 => \N__28154\,
            in1 => \N__28178\,
            in2 => \N__25465\,
            in3 => \N__27829\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_7_1_0__m5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__28177\,
            in1 => \N__28204\,
            in2 => \_gnd_net_\,
            in3 => \N__25461\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_1_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__28155\,
            in1 => \N__28179\,
            in2 => \N__25441\,
            in3 => \N__27830\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNIADII_0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__28176\,
            in1 => \N__28205\,
            in2 => \_gnd_net_\,
            in3 => \N__28151\,
            lcout => \DSW_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29467\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25475\,
            in2 => \N__28495\,
            in3 => \N__25423\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2_c\,
            carryout => \POWERLED.mult1_un138_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25420\,
            in2 => \N__25480\,
            in3 => \N__25411\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3_c\,
            carryout => \POWERLED.mult1_un138_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25408\,
            in2 => \N__26071\,
            in3 => \N__25399\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4_c\,
            carryout => \POWERLED.mult1_un138_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26070\,
            in2 => \N__25828\,
            in3 => \N__25816\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5_c\,
            carryout => \POWERLED.mult1_un138_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28272\,
            in1 => \N__25479\,
            in2 => \N__25813\,
            in3 => \N__25801\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6_c\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25789\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNO_0_15_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27828\,
            in2 => \_gnd_net_\,
            in3 => \N__27727\,
            lcout => \DSW_PWRGD.N_22_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25777\,
            in2 => \_gnd_net_\,
            in3 => \N__25684\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35108\,
            ce => \N__25624\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26061\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29488\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28442\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35700\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28516\,
            in1 => \N__25889\,
            in2 => \N__25906\,
            in3 => \_gnd_net_\,
            lcout => \G_2898\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28357\,
            in2 => \N__25894\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28342\,
            in2 => \N__28522\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28520\,
            in2 => \N__28597\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25893\,
            in2 => \N__28579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__28540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25879\,
            lcout => \POWERLED.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28447\,
            lcout => \POWERLED.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__25875\,
            in1 => \N__26820\,
            in2 => \_gnd_net_\,
            in3 => \N__29092\,
            lcout => \POWERLED.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26134\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29298\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28521\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26060\,
            lcout => \POWERLED.mult1_un131_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25993\,
            in2 => \N__26038\,
            in3 => \N__26026\,
            lcout => \POWERLED.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25987\,
            in1 => \N__25945\,
            in2 => \N__25957\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6108_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25912\,
            in2 => \N__28705\,
            in3 => \N__25939\,
            lcout => \POWERLED.N_6109_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26380\,
            in2 => \N__26419\,
            in3 => \N__26407\,
            lcout => \POWERLED.N_6110_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26341\,
            in2 => \N__26374\,
            in3 => \N__26365\,
            lcout => \POWERLED.N_6111_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26296\,
            in2 => \N__26335\,
            in3 => \N__26323\,
            lcout => \POWERLED.N_6112_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26290\,
            in1 => \N__26254\,
            in2 => \N__26266\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6113_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26248\,
            in1 => \N__26215\,
            in2 => \N__26224\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6114_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26209\,
            in1 => \N__26185\,
            in2 => \N__26686\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6115_i\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26140\,
            in2 => \N__26179\,
            in3 => \N__26164\,
            lcout => \POWERLED.N_6116_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26611\,
            in2 => \N__26650\,
            in3 => \N__26638\,
            lcout => \POWERLED.N_6117_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26605\,
            in1 => \N__26578\,
            in2 => \N__28747\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6118_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26568\,
            in1 => \N__26536\,
            in2 => \N__28480\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6119_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26530\,
            in1 => \N__26503\,
            in2 => \N__26770\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6120_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__26470\,
            in2 => \N__35491\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6121_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26464\,
            in1 => \N__26440\,
            in2 => \N__36196\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6122_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26434\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29241\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI2PKG_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31002\,
            in2 => \_gnd_net_\,
            in3 => \N__26821\,
            lcout => \POWERLED.g0_i_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35404\,
            lcout => \POWERLED.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJ2678_5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000011001"
        )
    port map (
            in0 => \N__31903\,
            in1 => \N__26758\,
            in2 => \N__26914\,
            in3 => \N__26658\,
            lcout => \N_96_mux_i_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2JIR8_6_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100101111"
        )
    port map (
            in0 => \N__26659\,
            in1 => \N__31904\,
            in2 => \N__27987\,
            in3 => \N__26872\,
            lcout => \N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_2_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32909\,
            lcout => \POWERLED.count_off_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI61QD3_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26863\,
            in1 => \N__26670\,
            in2 => \_gnd_net_\,
            in3 => \N__27076\,
            lcout => \POWERLED.un1_dutycycle_172_m4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110101111"
        )
    port map (
            in0 => \N__27153\,
            in1 => \N__27067\,
            in2 => \N__26855\,
            in3 => \N__29391\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3F2B2_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010100000"
        )
    port map (
            in0 => \N__26979\,
            in1 => \N__32910\,
            in2 => \N__27079\,
            in3 => \N__27154\,
            lcout => \POWERLED.un1_dutycycle_172_m1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_1_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__32911\,
            in1 => \N__26849\,
            in2 => \_gnd_net_\,
            in3 => \N__27069\,
            lcout => OPEN,
            ltout => \POWERLED.N_134_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3F2B2_0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__26980\,
            in1 => \N__26931\,
            in2 => \N__26917\,
            in3 => \N__30276\,
            lcout => \POWERLED.un1_dutycycle_172_m0\,
            ltout => \POWERLED.un1_dutycycle_172_m0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9JHG4_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__30277\,
            in1 => \N__26905\,
            in2 => \N__26887\,
            in3 => \N__26883\,
            lcout => \POWERLED.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_6_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__36823\,
            in1 => \_gnd_net_\,
            in2 => \N__27190\,
            in3 => \N__32172\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_6_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26857\,
            in2 => \N__26866\,
            in3 => \N__36151\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__26856\,
            in1 => \N__36649\,
            in2 => \_gnd_net_\,
            in3 => \N__32109\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__29392\,
            in1 => \N__36982\,
            in2 => \N__26824\,
            in3 => \N__36822\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__36983\,
            in1 => \N__36650\,
            in2 => \_gnd_net_\,
            in3 => \N__36530\,
            lcout => \POWERLED.N_361\,
            ltout => \POWERLED.N_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_3_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27186\,
            in2 => \N__27157\,
            in3 => \N__36150\,
            lcout => \POWERLED.dutycycle_RNI_9Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__37260\,
            in1 => \N__27145\,
            in2 => \N__32248\,
            in3 => \N__30386\,
            lcout => \POWERLED.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__27088\,
            in1 => \N__32872\,
            in2 => \N__27115\,
            in3 => \N__27099\,
            lcout => \POWERLED.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \N__32470\
        );

    \POWERLED.dutycycle_RNI_4_7_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__36977\,
            in1 => \_gnd_net_\,
            in2 => \N__37515\,
            in3 => \N__36654\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__36854\,
            in1 => \N__36973\,
            in2 => \_gnd_net_\,
            in3 => \N__32078\,
            lcout => \POWERLED.d_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__32079\,
            in1 => \N__36651\,
            in2 => \N__37002\,
            in3 => \N__36855\,
            lcout => OPEN,
            ltout => \POWERLED.un1_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_3_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__29262\,
            in1 => \N__27124\,
            in2 => \N__27118\,
            in3 => \N__30273\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJRE77_3_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32871\,
            in1 => \N__27111\,
            in2 => \N__27100\,
            in3 => \N__27087\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => \POWERLED.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_7_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__36652\,
            in1 => \_gnd_net_\,
            in2 => \N__27292\,
            in3 => \N__37501\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_8_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__30274\,
            in1 => \N__36653\,
            in2 => \N__27289\,
            in3 => \N__37334\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQU4T5_14_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__29946\,
            in1 => \N__30168\,
            in2 => \N__27268\,
            in3 => \N__29731\,
            lcout => \POWERLED.dutycycle_en_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGV14_13_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__32724\,
            in1 => \N__27257\,
            in2 => \N__36180\,
            in3 => \N__32894\,
            lcout => OPEN,
            ltout => \POWERLED.N_156_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQU4T5_13_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__29945\,
            in1 => \N__30167\,
            in2 => \N__27271\,
            in3 => \N__29730\,
            lcout => \POWERLED.dutycycle_en_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGV14_14_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__32319\,
            in1 => \N__27258\,
            in2 => \N__36181\,
            in3 => \N__32895\,
            lcout => \POWERLED.N_158_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIPB5N7_15_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32896\,
            in1 => \N__27354\,
            in2 => \N__27376\,
            in3 => \N__27196\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => \POWERLED.dutycycleZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGV14_15_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__32897\,
            in1 => \N__27259\,
            in2 => \N__27202\,
            in3 => \N__36176\,
            lcout => OPEN,
            ltout => \POWERLED.N_161_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQU4T5_15_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__29740\,
            in1 => \N__30166\,
            in2 => \N__27199\,
            in3 => \N__29944\,
            lcout => \POWERLED.dutycycle_en_12\,
            ltout => \POWERLED.dutycycle_en_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__27375\,
            in1 => \N__27355\,
            in2 => \N__27358\,
            in3 => \N__32893\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35254\,
            ce => 'H',
            sr => \N__32466\
        );

    \VPP_VDDQ.count_12_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27342\,
            lcout => \VPP_VDDQ.count_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34895\,
            ce => \N__27562\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_13_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27592\,
            lcout => \VPP_VDDQ.count_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34895\,
            ce => \N__27562\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_14_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27430\,
            lcout => \VPP_VDDQ.count_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34895\,
            ce => \N__27562\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_7_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27315\,
            lcout => \VPP_VDDQ.count_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34895\,
            ce => \N__27562\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI4AD02_15_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30742\,
            in1 => \N__27298\,
            in2 => \_gnd_net_\,
            in3 => \N__33361\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30741\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35075\,
            ce => \N__33362\,
            sr => \N__33579\
        );

    \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27396\,
            in1 => \N__30653\,
            in2 => \_gnd_net_\,
            in3 => \N__33360\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35075\,
            ce => \N__33362\,
            sr => \N__33579\
        );

    \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27604\,
            in1 => \N__30684\,
            in2 => \_gnd_net_\,
            in3 => \N__33359\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35075\,
            ce => \N__33362\,
            sr => \N__33579\
        );

    \VPP_VDDQ.count_RNIB8PO_13_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27598\,
            in1 => \N__27591\,
            in2 => \_gnd_net_\,
            in3 => \N__27554\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIDBQO_14_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27553\,
            in1 => \N__27436\,
            in2 => \_gnd_net_\,
            in3 => \N__27429\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__27685\,
            in1 => \N__33333\,
            in2 => \N__30727\,
            in3 => \N__30514\,
            lcout => \VPP_VDDQ.un29_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI27C02_14_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33330\,
            in1 => \N__27675\,
            in2 => \_gnd_net_\,
            in3 => \N__30782\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__27397\,
            in1 => \N__33332\,
            in2 => \N__30661\,
            in3 => \N__30627\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un29_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPT4L7_10_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27652\,
            in1 => \N__27667\,
            in2 => \N__27385\,
            in3 => \N__27382\,
            lcout => \VPP_VDDQ.un29_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34945\,
            ce => \N__33384\,
            sr => \N__33602\
        );

    \VPP_VDDQ.count_2_12_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30513\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34945\,
            ce => \N__33384\,
            sr => \N__33602\
        );

    \VPP_VDDQ.count_2_RNIU0A02_12_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27684\,
            in1 => \N__33329\,
            in2 => \_gnd_net_\,
            in3 => \N__30512\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI27C02_0_14_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010011"
        )
    port map (
            in0 => \N__33331\,
            in1 => \N__30756\,
            in2 => \N__30787\,
            in3 => \N__27676\,
            lcout => \VPP_VDDQ.un29_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIASDQ1_9_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33527\,
            in1 => \N__30612\,
            in2 => \N__27661\,
            in3 => \N__33327\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__30613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33578\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35079\,
            ce => \N__33355\,
            sr => \N__33576\
        );

    \VPP_VDDQ.count_2_11_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30544\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35079\,
            ce => \N__33355\,
            sr => \N__33576\
        );

    \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010001"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__27613\,
            in2 => \N__33387\,
            in3 => \N__30583\,
            lcout => \VPP_VDDQ.un29_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__27641\,
            in1 => \N__33526\,
            in2 => \_gnd_net_\,
            in3 => \N__31000\,
            lcout => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27612\,
            in2 => \N__27616\,
            in3 => \N__30581\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35079\,
            ce => \N__33355\,
            sr => \N__33576\
        );

    \DSW_PWRGD.DSW_PWROK_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__28132\,
            in1 => \N__28213\,
            in2 => \N__28068\,
            in3 => \N__27832\,
            lcout => dsw_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.DSW_PWROK_RNO_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28180\,
            in2 => \_gnd_net_\,
            in3 => \N__28156\,
            lcout => \DSW_PWRGD.curr_state10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28126\,
            in1 => \N__28114\,
            in2 => \N__28102\,
            in3 => \N__28064\,
            lcout => OPEN,
            ltout => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__28012\,
            in1 => \_gnd_net_\,
            in2 => \N__27994\,
            in3 => \N__27988\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNI09TK5_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27853\,
            in2 => \_gnd_net_\,
            in3 => \N__27831\,
            lcout => \un4_counter_7_c_RNI09TK5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIST802_11_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__33328\,
            in1 => \N__30543\,
            in2 => \N__27706\,
            in3 => \N__33575\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29484\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28247\,
            in2 => \N__27697\,
            in3 => \N__27688\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28333\,
            in2 => \N__28252\,
            in3 => \N__28327\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28274\,
            in2 => \N__28324\,
            in3 => \N__28315\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28312\,
            in2 => \N__28281\,
            in3 => \N__28306\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28437\,
            in1 => \N__28251\,
            in2 => \N__28303\,
            in3 => \N__28294\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28291\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28285\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28273\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29394\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28406\,
            in2 => \N__28237\,
            in3 => \N__28225\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28222\,
            in2 => \N__28411\,
            in3 => \N__28216\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28438\,
            in2 => \N__28465\,
            in3 => \N__28456\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28453\,
            in2 => \N__28446\,
            in3 => \N__28414\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28723\,
            in1 => \N__28410\,
            in2 => \N__28396\,
            in3 => \N__28387\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28378\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => \POWERLED.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28375\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32131\,
            in2 => \_gnd_net_\,
            in3 => \N__36690\,
            lcout => \POWERLED.g0_7_1\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28559\,
            in2 => \N__28372\,
            in3 => \N__28351\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28348\,
            in2 => \N__28564\,
            in3 => \N__28336\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28724\,
            in2 => \N__28606\,
            in3 => \N__28588\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28585\,
            in2 => \N__28731\,
            in3 => \N__28567\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28515\,
            in1 => \N__28563\,
            in2 => \N__28549\,
            in3 => \N__28534\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28525\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34383\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34312\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31558\,
            lcout => \POWERLED.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31428\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28732\,
            lcout => \POWERLED.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29197\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29135\,
            in2 => \N__28696\,
            in3 => \N__28675\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31396\,
            in2 => \N__29140\,
            in3 => \N__28657\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31378\,
            in2 => \N__31593\,
            in3 => \N__28642\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31588\,
            in2 => \N__31357\,
            in3 => \N__28624\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29151\,
            in1 => \N__29139\,
            in2 => \N__31336\,
            in3 => \N__28609\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29176\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__29022\,
            in1 => \N__29118\,
            in2 => \N__29096\,
            in3 => \N__29055\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35228\,
            ce => 'H',
            sr => \N__29011\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29639\,
            in2 => \N__29617\,
            in3 => \N__29760\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__29761\,
            in1 => \_gnd_net_\,
            in2 => \N__29644\,
            in3 => \N__29616\,
            lcout => \POWERLED.mult1_un40_sum_i_5\,
            ltout => \POWERLED.mult1_un40_sum_i_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28996\,
            in3 => \N__31684\,
            lcout => \POWERLED.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__31496\,
            in1 => \N__31497\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29638\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNII6Q06_7_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28993\,
            in1 => \N__28971\,
            in2 => \_gnd_net_\,
            in3 => \N__28804\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35684\,
            in2 => \N__37015\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35685\,
            in2 => \N__29656\,
            in3 => \N__29449\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29387\,
            in2 => \N__29446\,
            in3 => \N__29410\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29407\,
            in2 => \N__29395\,
            in3 => \N__29281\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29278\,
            in2 => \N__29266\,
            in3 => \N__29230\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30265\,
            in2 => \N__29227\,
            in3 => \N__29200\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30266\,
            in2 => \N__30187\,
            in3 => \N__29182\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36469\,
            in2 => \N__29593\,
            in3 => \N__29179\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31984\,
            in2 => \N__32215\,
            in3 => \N__29530\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37145\,
            in2 => \N__37039\,
            in3 => \N__29527\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32750\,
            in2 => \N__32491\,
            in3 => \N__29524\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32325\,
            in2 => \N__31930\,
            in3 => \N__29521\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30388\,
            in2 => \N__30340\,
            in3 => \N__29518\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32751\,
            in2 => \N__29665\,
            in3 => \N__29515\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32326\,
            in2 => \N__30325\,
            in3 => \N__29512\,
            lcout => \POWERLED.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30396\,
            in2 => \N__29509\,
            in3 => \N__29494\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30397\,
            in2 => \N__29749\,
            in3 => \N__29491\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29764\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32312\,
            in2 => \_gnd_net_\,
            in3 => \N__32608\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29729\,
            lcout => \POWERLED.func_state_RNI_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_13_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \N__32748\,
            in1 => \N__35899\,
            in2 => \N__32230\,
            in3 => \N__29677\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36655\,
            in1 => \N__35699\,
            in2 => \_gnd_net_\,
            in3 => \N__32123\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29643\,
            in3 => \N__29612\,
            lcout => \POWERLED.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_9_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__36878\,
            in1 => \N__30286\,
            in2 => \_gnd_net_\,
            in3 => \N__37280\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_7_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__37509\,
            in1 => \N__36880\,
            in2 => \N__29596\,
            in3 => \N__36462\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILUF77_4_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__29581\,
            in1 => \N__32937\,
            in2 => \N__29566\,
            in3 => \N__29545\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_9_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110101000"
        )
    port map (
            in0 => \N__37278\,
            in1 => \N__36877\,
            in2 => \N__30292\,
            in3 => \N__36561\,
            lcout => OPEN,
            ltout => \POWERLED.g0_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__37360\,
            in1 => \N__36456\,
            in2 => \N__30289\,
            in3 => \N__37279\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_7_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010111"
        )
    port map (
            in0 => \N__36647\,
            in1 => \N__36978\,
            in2 => \N__37516\,
            in3 => \N__37358\,
            lcout => \POWERLED.un1_dutycycle_53_25_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_7_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001000"
        )
    port map (
            in0 => \N__37359\,
            in1 => \N__36648\,
            in2 => \N__37003\,
            in3 => \N__37508\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_9_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__37281\,
            in1 => \N__36879\,
            in2 => \N__30280\,
            in3 => \N__30275\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__29995\,
            in1 => \N__30001\,
            in2 => \N__29969\,
            in3 => \N__29983\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \N__32467\
        );

    \POWERLED.dutycycle_RNI778D2_12_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101111"
        )
    port map (
            in0 => \N__37110\,
            in1 => \N__30169\,
            in2 => \N__32951\,
            in3 => \N__30022\,
            lcout => \POWERLED.dutycycle_eena_9\,
            ltout => \POWERLED.dutycycle_eena_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI24QN4_12_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__29994\,
            in1 => \N__29982\,
            in2 => \N__29974\,
            in3 => \N__29951\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => \POWERLED.dutycycleZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30412\,
            in3 => \N__30373\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111010010"
        )
    port map (
            in0 => \N__31976\,
            in1 => \N__30409\,
            in2 => \N__30403\,
            in3 => \N__36339\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30400\,
            in3 => \N__30374\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010011010"
        )
    port map (
            in0 => \N__32335\,
            in1 => \N__32679\,
            in2 => \N__37150\,
            in3 => \N__36340\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30328\,
            in3 => \N__32324\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__33405\,
            in1 => \N__30313\,
            in2 => \N__30451\,
            in3 => \N__30301\,
            lcout => \VPP_VDDQ.un29_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__30462\,
            in1 => \N__33049\,
            in2 => \N__30481\,
            in3 => \N__33559\,
            lcout => \VPP_VDDQ.count_2_rst_6\,
            ltout => \VPP_VDDQ.count_2_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS66Q1_2_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30300\,
            in2 => \N__30307\,
            in3 => \N__33385\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_2\,
            ltout => \VPP_VDDQ.un1_count_2_1_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__30463\,
            in1 => \N__33054\,
            in2 => \N__30304\,
            in3 => \N__33563\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35215\,
            ce => \N__33404\,
            sr => \N__33547\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__33560\,
            in1 => \N__30429\,
            in2 => \N__33065\,
            in3 => \N__30450\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU97Q1_3_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33386\,
            in1 => \_gnd_net_\,
            in2 => \N__30493\,
            in3 => \N__30487\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => \VPP_VDDQ.count_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__33561\,
            in1 => \N__30430\,
            in2 => \N__30490\,
            in3 => \N__33060\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35215\,
            ce => \N__33404\,
            sr => \N__33547\
        );

    \VPP_VDDQ.count_2_0_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33681\,
            in1 => \N__33053\,
            in2 => \_gnd_net_\,
            in3 => \N__33562\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35215\,
            ce => \N__33404\,
            sr => \N__33547\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33697\,
            in2 => \N__33680\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30480\,
            in3 => \N__30454\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30446\,
            in2 => \_gnd_net_\,
            in3 => \N__30421\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33569\,
            in1 => \N__33216\,
            in2 => \_gnd_net_\,
            in3 => \N__30418\,
            lcout => \VPP_VDDQ.count_2_rst_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33142\,
            in2 => \_gnd_net_\,
            in3 => \N__30415\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33570\,
            in1 => \N__33102\,
            in2 => \_gnd_net_\,
            in3 => \N__30673\,
            lcout => \VPP_VDDQ.count_2_rst_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33606\,
            in1 => \N__30670\,
            in2 => \_gnd_net_\,
            in3 => \N__30637\,
            lcout => \VPP_VDDQ.count_2_rst_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32568\,
            in3 => \N__30634\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30631\,
            in2 => \_gnd_net_\,
            in3 => \N__30598\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33571\,
            in1 => \N__30595\,
            in2 => \_gnd_net_\,
            in3 => \N__30565\,
            lcout => \VPP_VDDQ.count_2_rst_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30562\,
            in2 => \_gnd_net_\,
            in3 => \N__30526\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33572\,
            in1 => \N__30523\,
            in2 => \_gnd_net_\,
            in3 => \N__30499\,
            lcout => \VPP_VDDQ.count_2_rst_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30720\,
            in2 => \_gnd_net_\,
            in3 => \N__30496\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33573\,
            in1 => \N__30796\,
            in2 => \_gnd_net_\,
            in3 => \N__30766\,
            lcout => \VPP_VDDQ.count_2_rst_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__30763\,
            in1 => \N__33574\,
            in2 => \_gnd_net_\,
            in3 => \N__30745\,
            lcout => \VPP_VDDQ.count_2_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI04B02_13_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33383\,
            in1 => \N__33551\,
            in2 => \N__33625\,
            in3 => \N__33636\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI_0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34158\,
            in2 => \_gnd_net_\,
            in3 => \N__33838\,
            lcout => OPEN,
            ltout => \HDA_STRAP.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNINQ6P_0_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30697\,
            in2 => \N__30709\,
            in3 => \N__34515\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => \HDA_STRAP.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI68FK1_1_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33202\,
            in1 => \N__33919\,
            in2 => \N__30706\,
            in3 => \N__30802\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un25_clk_100khz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI6OA47_8_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30817\,
            in1 => \N__30691\,
            in2 => \N__30703\,
            in3 => \N__31207\,
            lcout => \HDA_STRAP.count_RNI6OA47Z0Z_8\,
            ltout => \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30700\,
            in3 => \N__33837\,
            lcout => \HDA_STRAP.count_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35010\,
            ce => \N__34448\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNILLET_0_8_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__33940\,
            in1 => \N__34517\,
            in2 => \N__30847\,
            in3 => \N__33975\,
            lcout => \HDA_STRAP.un25_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35010\,
            ce => \N__34448\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNILLET_8_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30843\,
            in1 => \N__34516\,
            in2 => \_gnd_net_\,
            in3 => \N__33974\,
            lcout => \HDA_STRAP.un2_count_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34015\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35121\,
            ce => \N__34447\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35121\,
            ce => \N__34447\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDB8R_15_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34512\,
            in1 => \N__30828\,
            in2 => \_gnd_net_\,
            in3 => \N__34241\,
            lcout => \HDA_STRAP.un2_count_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIHFCT_6_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30835\,
            in1 => \N__34511\,
            in2 => \_gnd_net_\,
            in3 => \N__34014\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => \HDA_STRAP.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDB8R_0_15_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__34514\,
            in1 => \N__30829\,
            in2 => \N__30820\,
            in3 => \N__34242\,
            lcout => \HDA_STRAP.un25_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIEC8R_16_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30811\,
            in1 => \N__34214\,
            in2 => \_gnd_net_\,
            in3 => \N__34513\,
            lcout => \HDA_STRAP.un2_count_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34215\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35121\,
            ce => \N__34447\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIEC8R_0_16_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__30810\,
            in1 => \N__34510\,
            in2 => \N__34219\,
            in3 => \N__34102\,
            lcout => \HDA_STRAP.un25_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33883\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35159\,
            ce => \N__34446\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35159\,
            ce => \N__34446\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNINOFT_9_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34531\,
            in1 => \N__30858\,
            in2 => \_gnd_net_\,
            in3 => \N__33953\,
            lcout => \HDA_STRAP.un2_count_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB0VU_12_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30865\,
            in1 => \N__33882\,
            in2 => \_gnd_net_\,
            in3 => \N__34533\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => \HDA_STRAP.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNINOFT_0_9_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__34534\,
            in1 => \N__30859\,
            in2 => \N__30850\,
            in3 => \N__33954\,
            lcout => \HDA_STRAP.un25_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIFCBT_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__34530\,
            in2 => \_gnd_net_\,
            in3 => \N__33716\,
            lcout => \HDA_STRAP.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35159\,
            ce => \N__34446\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI0THV_10_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34030\,
            in1 => \N__34041\,
            in2 => \_gnd_net_\,
            in3 => \N__34532\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB69T_0_3_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__34524\,
            in1 => \N__31177\,
            in2 => \N__33766\,
            in3 => \N__33744\,
            lcout => \HDA_STRAP.un25_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33765\,
            lcout => \HDA_STRAP.count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35227\,
            ce => \N__34444\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIFCBT_0_5_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__34525\,
            in1 => \N__33999\,
            in2 => \N__31240\,
            in3 => \N__33721\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un25_clk_100khz_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIUE4N3_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31198\,
            in1 => \N__31225\,
            in2 => \N__31219\,
            in3 => \N__31216\,
            lcout => \HDA_STRAP.un25_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNID30V_0_13_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__34526\,
            in1 => \N__34266\,
            in2 => \N__31192\,
            in3 => \N__33864\,
            lcout => \HDA_STRAP.un25_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35227\,
            ce => \N__34444\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNID30V_13_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34523\,
            in1 => \N__31188\,
            in2 => \_gnd_net_\,
            in3 => \N__33863\,
            lcout => \HDA_STRAP.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB69T_3_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31176\,
            in1 => \N__33761\,
            in2 => \_gnd_net_\,
            in3 => \N__34522\,
            lcout => \HDA_STRAP.un2_count_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111011101"
        )
    port map (
            in0 => \N__31166\,
            in1 => \N__31012\,
            in2 => \N__31051\,
            in3 => \N__31005\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31078\,
            in2 => \_gnd_net_\,
            in3 => \N__31047\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35160\,
            ce => \N__30953\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNID9AT_4_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34072\,
            in1 => \N__34527\,
            in2 => \_gnd_net_\,
            in3 => \N__34086\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIF61V_14_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34529\,
            in1 => \N__35347\,
            in2 => \_gnd_net_\,
            in3 => \N__35361\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIJIDT_7_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34065\,
            in1 => \N__34051\,
            in2 => \_gnd_net_\,
            in3 => \N__34528\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31291\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31442\,
            in2 => \N__31270\,
            in3 => \N__31255\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34366\,
            in2 => \N__31447\,
            in3 => \N__31252\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34304\,
            in2 => \N__34357\,
            in3 => \N__31249\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34345\,
            in2 => \N__34311\,
            in3 => \N__31246\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31548\,
            in1 => \N__31446\,
            in2 => \N__34336\,
            in3 => \N__31243\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31450\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34303\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31524\,
            in2 => \N__31411\,
            in3 => \N__31387\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31384\,
            in2 => \N__31528\,
            in3 => \N__31369\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31550\,
            in2 => \N__31366\,
            in3 => \N__31345\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31342\,
            in2 => \N__31557\,
            in3 => \N__31324\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31574\,
            in1 => \N__31523\,
            in2 => \N__31321\,
            in3 => \N__31303\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31294\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31549\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36307\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31855\,
            in3 => \N__31513\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31633\,
            in2 => \N__31615\,
            in3 => \N__31510\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31662\,
            in2 => \N__31726\,
            in3 => \N__31507\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31658\,
            in2 => \N__31699\,
            in3 => \N__31504\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35555\,
            in1 => \N__31501\,
            in2 => \N__31480\,
            in3 => \N__31468\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31680\,
            in2 => \N__31465\,
            in3 => \N__31453\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => \POWERLED.mult1_un54_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31762\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31879\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31759\,
            in3 => \N__31744\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31741\,
            in3 => \N__31717\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31654\,
            in2 => \N__31714\,
            in3 => \N__31690\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31687\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__31631\,
            in1 => \N__31632\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37005\,
            lcout => \POWERLED.un1_clk_100khz_43_and_i_0_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__32121\,
            in1 => \N__35693\,
            in2 => \_gnd_net_\,
            in3 => \N__32177\,
            lcout => OPEN,
            ltout => \POWERLED.m21_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_6_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011111"
        )
    port map (
            in0 => \N__36870\,
            in1 => \N__35947\,
            in2 => \N__31909\,
            in3 => \N__31830\,
            lcout => \POWERLED.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31875\,
            lcout => \POWERLED.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__36871\,
            in1 => \N__31843\,
            in2 => \N__35701\,
            in3 => \N__31831\,
            lcout => \POWERLED.g0_10_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_0_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35692\,
            in2 => \_gnd_net_\,
            in3 => \N__32176\,
            lcout => OPEN,
            ltout => \POWERLED.g2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_1_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__36869\,
            in1 => \N__31829\,
            in2 => \N__31765\,
            in3 => \N__32120\,
            lcout => \POWERLED.g0_10_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_8_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110001"
        )
    port map (
            in0 => \N__36846\,
            in1 => \N__36699\,
            in2 => \N__36551\,
            in3 => \N__37365\,
            lcout => \POWERLED.un1_dutycycle_53_10_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36465\,
            in2 => \_gnd_net_\,
            in3 => \N__37147\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_4_a1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_8_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36848\,
            in1 => \N__36700\,
            in2 => \N__32233\,
            in3 => \N__37369\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_7_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011111110"
        )
    port map (
            in0 => \N__32200\,
            in1 => \N__36847\,
            in2 => \N__37397\,
            in3 => \N__37492\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_9_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \N__31975\,
            in1 => \N__36907\,
            in2 => \N__32218\,
            in3 => \N__37021\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110111"
        )
    port map (
            in0 => \N__36698\,
            in1 => \N__37255\,
            in2 => \N__37396\,
            in3 => \N__37008\,
            lcout => \POWERLED.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_7_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37511\,
            in3 => \N__37361\,
            lcout => \POWERLED.un1_dutycycle_53_4_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__36865\,
            in1 => \N__32178\,
            in2 => \N__32130\,
            in3 => \N__35698\,
            lcout => \POWERLED.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_10_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101000"
        )
    port map (
            in0 => \N__37276\,
            in1 => \N__31915\,
            in2 => \N__36472\,
            in3 => \N__37400\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__36461\,
            in1 => \N__32322\,
            in2 => \N__31987\,
            in3 => \N__31974\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_9_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001001010"
        )
    port map (
            in0 => \N__36556\,
            in1 => \N__36867\,
            in2 => \N__37292\,
            in3 => \N__36683\,
            lcout => \POWERLED.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32531\,
            in2 => \_gnd_net_\,
            in3 => \N__36659\,
            lcout => \POWERLED.un1_clk_100khz_40_and_i_0_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_8_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__36660\,
            in1 => \N__32673\,
            in2 => \N__36562\,
            in3 => \N__37398\,
            lcout => \POWERLED.un1_dutycycle_53_49_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_9_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__36682\,
            in1 => \N__37271\,
            in2 => \_gnd_net_\,
            in3 => \N__36555\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_6Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_8_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__37275\,
            in1 => \N__36868\,
            in2 => \N__32494\,
            in3 => \N__37399\,
            lcout => \POWERLED.un1_dutycycle_53_34_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36460\,
            in1 => \N__37277\,
            in2 => \N__32752\,
            in3 => \N__36886\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_9_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__36866\,
            in1 => \N__37222\,
            in2 => \N__32680\,
            in3 => \N__36559\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32992\,
            in1 => \N__32980\,
            in2 => \N__32968\,
            in3 => \N__32933\,
            lcout => \POWERLED.dutycycleZ1Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \N__32469\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32320\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32711\,
            lcout => \POWERLED.un1_dutycycle_53_axb_14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_13_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32712\,
            in1 => \N__32321\,
            in2 => \N__37415\,
            in3 => \N__36464\,
            lcout => \POWERLED.un2_count_clk_17_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_8_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010101"
        )
    port map (
            in0 => \N__32677\,
            in1 => \N__36560\,
            in2 => \N__36706\,
            in3 => \N__37401\,
            lcout => \POWERLED.un1_dutycycle_53_2_1_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIL53N7_13_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32991\,
            in1 => \N__32979\,
            in2 => \N__32967\,
            in3 => \N__32932\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => \POWERLED.dutycycleZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__36463\,
            in1 => \N__32678\,
            in2 => \N__32620\,
            in3 => \N__37125\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_9_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__37223\,
            in1 => \N__32617\,
            in2 => \N__32611\,
            in3 => \N__36352\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33231\,
            lcout => \VPP_VDDQ.count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35080\,
            ce => \N__33403\,
            sr => \N__33615\
        );

    \VPP_VDDQ.count_2_8_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__32564\,
            in1 => \N__33616\,
            in2 => \N__33066\,
            in3 => \N__32590\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35080\,
            ce => \N__33403\,
            sr => \N__33615\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__32589\,
            in1 => \N__33055\,
            in2 => \N__32569\,
            in3 => \N__33604\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32578\,
            in2 => \N__32572\,
            in3 => \N__33388\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => \VPP_VDDQ.count_2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__33118\,
            in1 => \N__33151\,
            in2 => \N__32545\,
            in3 => \N__33391\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un29_clk_100khz_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINKK9B_2_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33175\,
            in1 => \N__33169\,
            in2 => \N__33157\,
            in3 => \N__33085\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => \VPP_VDDQ.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__33130\,
            in1 => \N__33141\,
            in2 => \N__33154\,
            in3 => \N__33603\,
            lcout => \VPP_VDDQ.count_2_rst_3\,
            ltout => \VPP_VDDQ.count_2_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33117\,
            in2 => \N__33145\,
            in3 => \N__33389\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_5\,
            ltout => \VPP_VDDQ.un1_count_2_1_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__33129\,
            in1 => \N__33056\,
            in2 => \N__33121\,
            in3 => \N__33605\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35120\,
            ce => \N__33390\,
            sr => \N__33601\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33109\,
            in1 => \N__33217\,
            in2 => \N__33682\,
            in3 => \N__33695\,
            lcout => \VPP_VDDQ.un29_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINUSC_0_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33679\,
            in1 => \N__33064\,
            in2 => \_gnd_net_\,
            in3 => \N__33549\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIC4UI1_0_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33007\,
            in2 => \N__32998\,
            in3 => \N__33380\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINUSC_1_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__33696\,
            in1 => \_gnd_net_\,
            in2 => \N__32995\,
            in3 => \N__33548\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID5UI1_1_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33643\,
            in2 => \N__33700\,
            in3 => \N__33382\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => \VPP_VDDQ.count_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33675\,
            in2 => \N__33646\,
            in3 => \N__33600\,
            lcout => \VPP_VDDQ.count_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35082\,
            ce => \N__33406\,
            sr => \N__33599\
        );

    \VPP_VDDQ.count_2_13_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33637\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35082\,
            ce => \N__33406\,
            sr => \N__33599\
        );

    \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__33381\,
            in1 => \N__33241\,
            in2 => \N__33232\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI938T_2_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34519\,
            in1 => \_gnd_net_\,
            in2 => \N__33790\,
            in3 => \N__33850\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => \HDA_STRAP.countZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIOR6P_0_1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__33196\,
            in1 => \N__33184\,
            in2 => \N__33205\,
            in3 => \N__34521\,
            lcout => \HDA_STRAP.un25_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI_1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33810\,
            in1 => \N__33834\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_RNIZ0Z_1\,
            ltout => \HDA_STRAP.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIOR6P_1_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33183\,
            in2 => \N__33190\,
            in3 => \N__34518\,
            lcout => \HDA_STRAP.un2_count_1_axb_1\,
            ltout => \HDA_STRAP.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33835\,
            in2 => \N__33187\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35017\,
            ce => \N__34449\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33789\,
            lcout => \HDA_STRAP.count_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35017\,
            ce => \N__34449\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI9TTU_11_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34520\,
            in1 => \N__33844\,
            in2 => \_gnd_net_\,
            in3 => \N__33903\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35017\,
            ce => \N__34449\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_1_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33836\,
            in2 => \N__33814\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \HDA_STRAP.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33796\,
            in2 => \_gnd_net_\,
            in3 => \N__33778\,
            lcout => \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_1\,
            carryout => \HDA_STRAP.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33775\,
            in2 => \_gnd_net_\,
            in3 => \N__33748\,
            lcout => \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_2\,
            carryout => \HDA_STRAP.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33745\,
            in2 => \_gnd_net_\,
            in3 => \N__33730\,
            lcout => \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_3\,
            carryout => \HDA_STRAP.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33727\,
            in2 => \_gnd_net_\,
            in3 => \N__33703\,
            lcout => \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_4\,
            carryout => \HDA_STRAP.un2_count_1_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34159\,
            in1 => \N__34021\,
            in2 => \_gnd_net_\,
            in3 => \N__34006\,
            lcout => \HDA_STRAP.count_1_6\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_5_cZ0\,
            carryout => \HDA_STRAP.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34003\,
            in2 => \_gnd_net_\,
            in3 => \N__33985\,
            lcout => \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_6\,
            carryout => \HDA_STRAP.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34160\,
            in1 => \N__33982\,
            in2 => \_gnd_net_\,
            in3 => \N__33964\,
            lcout => \HDA_STRAP.count_1_8\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_7\,
            carryout => \HDA_STRAP.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33961\,
            in2 => \_gnd_net_\,
            in3 => \N__33943\,
            lcout => \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \HDA_STRAP.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__34185\,
            in1 => \_gnd_net_\,
            in2 => \N__33939\,
            in3 => \N__33922\,
            lcout => \HDA_STRAP.count_1_10\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_9\,
            carryout => \HDA_STRAP.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34187\,
            in1 => \N__33918\,
            in2 => \_gnd_net_\,
            in3 => \N__33892\,
            lcout => \HDA_STRAP.count_1_11\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_10\,
            carryout => \HDA_STRAP.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33889\,
            in2 => \_gnd_net_\,
            in3 => \N__33874\,
            lcout => \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_11\,
            carryout => \HDA_STRAP.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33871\,
            in2 => \_gnd_net_\,
            in3 => \N__33853\,
            lcout => \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_12\,
            carryout => \HDA_STRAP.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34267\,
            in2 => \_gnd_net_\,
            in3 => \N__34252\,
            lcout => \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_13\,
            carryout => \HDA_STRAP.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34249\,
            in2 => \_gnd_net_\,
            in3 => \N__34231\,
            lcout => \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_14\,
            carryout => \HDA_STRAP.un2_count_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__34186\,
            in1 => \_gnd_net_\,
            in2 => \N__34228\,
            in3 => \N__34201\,
            lcout => \HDA_STRAP.count_1_16\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_15\,
            carryout => \HDA_STRAP.un2_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34101\,
            in1 => \N__34188\,
            in2 => \_gnd_net_\,
            in3 => \N__34135\,
            lcout => \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNILF4V_17_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34128\,
            in1 => \N__34114\,
            in2 => \_gnd_net_\,
            in3 => \N__34509\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34087\,
            lcout => \HDA_STRAP.count_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35151\,
            ce => \N__34445\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34066\,
            lcout => \HDA_STRAP.count_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35151\,
            ce => \N__34445\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34045\,
            lcout => \HDA_STRAP.count_1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35151\,
            ce => \N__34445\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35362\,
            lcout => \HDA_STRAP.count_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35151\,
            ce => \N__34445\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34387\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34277\,
            in2 => \N__35920\,
            in3 => \N__34360\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35458\,
            in2 => \N__34282\,
            in3 => \N__34348\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35393\,
            in2 => \N__35449\,
            in3 => \N__34339\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35437\,
            in2 => \N__35400\,
            in3 => \N__34327\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34302\,
            in1 => \N__34281\,
            in2 => \N__35428\,
            in3 => \N__34318\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34315\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35392\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35941\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35732\,
            in2 => \N__35371\,
            in3 => \N__35452\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35890\,
            in2 => \N__35737\,
            in3 => \N__35440\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35872\,
            in2 => \N__35767\,
            in3 => \N__35431\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35766\,
            in2 => \N__35854\,
            in3 => \N__35419\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35391\,
            in1 => \N__35736\,
            in2 => \N__35830\,
            in3 => \N__35410\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35788\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35407\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35476\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36274\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36283\,
            in2 => \N__35523\,
            in3 => \N__35584\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35519\,
            in2 => \N__35581\,
            in3 => \N__35572\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35569\,
            in2 => \N__35560\,
            in3 => \N__35563\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35559\,
            in2 => \N__35542\,
            in3 => \N__35533\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36225\,
            in1 => \N__35530\,
            in2 => \N__35524\,
            in3 => \N__35506\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35503\,
            in3 => \N__35494\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35757\,
            lcout => \POWERLED.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35475\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35807\,
            in2 => \N__36253\,
            in3 => \N__35881\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35878\,
            in2 => \N__35812\,
            in3 => \N__35863\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35860\,
            in2 => \N__36236\,
            in3 => \N__35839\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35836\,
            in2 => \N__36237\,
            in3 => \N__35815\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35756\,
            in1 => \N__35811\,
            in2 => \N__35797\,
            in3 => \N__35779\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35770\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => \POWERLED.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35740\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__37006\,
            in1 => \N__36177\,
            in2 => \N__35719\,
            in3 => \N__35697\,
            lcout => \POWERLED.g3_1_3_0\,
            ltout => \POWERLED.g3_1_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110010"
        )
    port map (
            in0 => \N__36044\,
            in1 => \N__36179\,
            in2 => \N__36325\,
            in3 => \N__36322\,
            lcout => \POWERLED.N_3034_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36303\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36273\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36235\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011100"
        )
    port map (
            in0 => \N__36178\,
            in1 => \N__36052\,
            in2 => \N__36046\,
            in3 => \N__35953\,
            lcout => \POWERLED.N_3034_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35937\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36471\,
            in2 => \N__35908\,
            in3 => \N__37148\,
            lcout => \POWERLED.un1_dutycycle_53_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_8_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36692\,
            in2 => \_gnd_net_\,
            in3 => \N__37412\,
            lcout => \POWERLED.un1_dutycycle_53_4_a0_1\,
            ltout => \POWERLED.un1_dutycycle_53_4_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_9_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110111"
        )
    port map (
            in0 => \N__36916\,
            in1 => \N__36876\,
            in2 => \N__37024\,
            in3 => \N__37259\,
            lcout => \POWERLED.un1_dutycycle_53_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__36691\,
            in1 => \N__37007\,
            in2 => \N__37282\,
            in3 => \N__36522\,
            lcout => \POWERLED.un1_dutycycle_53_31_a1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_7_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100110011"
        )
    port map (
            in0 => \N__36693\,
            in1 => \N__37514\,
            in2 => \N__37283\,
            in3 => \N__37413\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_9_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011111011"
        )
    port map (
            in0 => \N__37414\,
            in1 => \N__36875\,
            in2 => \N__36910\,
            in3 => \N__36523\,
            lcout => \POWERLED.un1_dutycycle_53_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_8_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__36558\,
            in1 => \_gnd_net_\,
            in2 => \N__37416\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_31_a7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_7_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__36873\,
            in1 => \N__37513\,
            in2 => \N__36901\,
            in3 => \N__36894\,
            lcout => \POWERLED.un1_dutycycle_53_34_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__36478\,
            in1 => \N__36874\,
            in2 => \N__36898\,
            in3 => \N__37423\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__36872\,
            in1 => \N__36697\,
            in2 => \N__37293\,
            in3 => \N__36557\,
            lcout => \POWERLED.un1_dutycycle_53_39_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_10_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__36470\,
            in1 => \N__37290\,
            in2 => \N__36361\,
            in3 => \N__36351\,
            lcout => \POWERLED.un1_dutycycle_53_49_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37512\,
            in2 => \N__37294\,
            in3 => \N__37405\,
            lcout => \POWERLED.un1_dutycycle_53_39_c_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_8_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37417\,
            in3 => \N__37291\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_36_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_12_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \N__37149\,
            in1 => \N__37054\,
            in2 => \N__37048\,
            in3 => \N__37045\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
