-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 7 2022 10:06:35

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : out std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_1_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_0\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_16\ : std_logic;
signal \HDA_STRAP.curr_state_RNIH91AZ0Z_1\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \POWERLED.count_0_4\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \POWERLED.count_0_5\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.count_1_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_0_1\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.count_0_12\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.curr_state_3_0_cascade_\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \POWERLED.count_1_0_cascade_\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal \POWERLED.g0_i_o3_0\ : std_logic;
signal \POWERLED.un79_clk_100khzlt6_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_3\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \POWERLED.N_8\ : std_logic;
signal \POWERLED.un1_count_cry_0_i\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \POWERLED.N_5110_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.N_5111_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.N_5112_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.N_5113_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.N_5114_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.N_5115_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.N_5116_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.N_5117_i\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \POWERLED.N_5118_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.N_5119_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.N_5120_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.N_5121_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.N_5122_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.N_5123_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.N_5124_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_9\ : std_logic;
signal \POWERLED.un85_clk_100khz_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_10\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_3\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_0\ : std_logic;
signal \HDA_STRAP.un4_count_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_5\ : std_logic;
signal \HDA_STRAP.un4_count_10\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_17\ : std_logic;
signal \HDA_STRAP.countZ0Z_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \HDA_STRAP.un4_count_9_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_13\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_16\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.countZ0Z_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un4_count_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.un4_count_12\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_6\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_8\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.N_14_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal hda_sdo_atp : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \HDA_STRAP.curr_state_RNO_0Z0Z_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.N_5_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_14\ : std_logic;
signal \DSW_PWRGD.countZ0Z_13\ : std_logic;
signal \DSW_PWRGD.countZ0Z_15\ : std_logic;
signal \DSW_PWRGD.countZ0Z_12\ : std_logic;
signal \DSW_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_2\ : std_logic;
signal \DSW_PWRGD.countZ0Z_5\ : std_logic;
signal \DSW_PWRGD.countZ0Z_7\ : std_logic;
signal \DSW_PWRGD.countZ0Z_3\ : std_logic;
signal \DSW_PWRGD.un4_count_10\ : std_logic;
signal \DSW_PWRGD.countZ0Z_11\ : std_logic;
signal \DSW_PWRGD.countZ0Z_10\ : std_logic;
signal \DSW_PWRGD.countZ0Z_8\ : std_logic;
signal \DSW_PWRGD.countZ0Z_0\ : std_logic;
signal \DSW_PWRGD.un4_count_11\ : std_logic;
signal \DSW_PWRGD.un1_curr_state10_0\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal v33dsw_ok : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \DSW_PWRGD.N_1_i\ : std_logic;
signal \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal \G_27\ : std_logic;
signal \G_27_cascade_\ : std_logic;
signal \DSW_PWRGD.N_29_1\ : std_logic;
signal \POWERLED.d_i1_mux_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_16Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.d_i3_mux_cascade_\ : std_logic;
signal \POWERLED.un1_i3_mux\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal \POWERLED.count_0_2\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.count_1_2\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.count_1_3\ : std_logic;
signal \POWERLED.un1_count_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.count_1_4\ : std_logic;
signal \POWERLED.un1_count_cry_3\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.count_1_5\ : std_logic;
signal \POWERLED.un1_count_cry_4\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.count_1_10\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.count_1_11\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.count_1_12\ : std_logic;
signal \POWERLED.un1_count_cry_11_cZ0\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.count_1_13\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\ : std_logic;
signal \POWERLED.un1_count_cry_13_cZ0\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.count_1_9\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.count_1_6\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.count_1_7\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.count_1_8\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un85_clk_100khz_7\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2_c\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_c\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_c\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_c\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_c\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \POWERLED.count_offZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.count_off_0_3\ : std_logic;
signal \POWERLED.count_off_0_7\ : std_logic;
signal \DSW_PWRGD.countZ0Z_1\ : std_logic;
signal \DSW_PWRGD.countZ0Z_6\ : std_logic;
signal \DSW_PWRGD.countZ0Z_9\ : std_logic;
signal \DSW_PWRGD.countZ0Z_4\ : std_logic;
signal \DSW_PWRGD.un4_count_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_20_0_0\ : std_logic;
signal \POWERLED.o2_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_7_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_4_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_2_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_2_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_12_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_56_a0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_56_a1_1\ : std_logic;
signal \POWERLED.un1_clk_100khz_45_and_i_i_a3_0_0_cascade_\ : std_logic;
signal \POWERLED.N_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_3_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_3\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \POWERLED.dutycycle_eena_3_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_3_1\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_1_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_5_cascade_\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal v5s_enn : std_logic;
signal \POWERLED.mult1_un47_sum_i\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal v33a_enn : std_logic;
signal \POWERLED.un85_clk_100khz_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \POWERLED.mult1_un75_sum_i_8\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \bfn_5_1_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \POWERLED.count_off_0_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_off_0_11\ : std_logic;
signal \POWERLED.dutycycle_eena_8_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_8\ : std_logic;
signal \POWERLED.dutycycleZ1Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_4_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_4\ : std_logic;
signal \POWERLED.dutycycle_eena_4_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \POWERLED.dutycycle_eena_5_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_5_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_6_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_6\ : std_logic;
signal \POWERLED.dutycycle_eena_6_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \POWERLED.dutycycle_eena_5\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.N_4_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_12_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_48_and_i_i_a3_0_0\ : std_logic;
signal \POWERLED.dutycycle_en_12\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_12_cascade_\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_3\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.curr_state_1_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_9Z0Z_9\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_5\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_4_sf\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un85_clk_100khz_4\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal pch_pwrok : std_logic;
signal vccst_pwrgd : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.count_off_1_8\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_off_1_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_off_1_12\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \POWERLED.dutycycleZ1Z_14\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_13Z0Z_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_11_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_4\ : std_logic;
signal \POWERLED.dutycycle_en_7_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_39_and_i_0_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_30_and_i_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI4J2O7Z0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI4J2O7Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_11\ : std_logic;
signal \POWERLED.dutycycle_en_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_20_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_3_2_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_3_2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_10\ : std_logic;
signal \POWERLED.dutycycleZ1Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_50_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_12Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_15Z0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI_11Z0Z_9\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_2\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_3\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_4\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_9\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_11\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_12\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.mult1_un47_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.g2_1\ : std_logic;
signal \POWERLED.g2_5\ : std_logic;
signal \POWERLED.g0_4_4\ : std_logic;
signal \POWERLED.g0_4_5_cascade_\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.g3_1_0\ : std_logic;
signal \POWERLED.g3_1_4_cascade_\ : std_logic;
signal \POWERLED.g3_1_6_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un85_clk_100khz_2\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un145_sum\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_4_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \PCH_PWRGD_delayed_vccin_ok\ : std_logic;
signal \PCH_PWRGD.N_250_0\ : std_logic;
signal \PCH_PWRGD.N_250_0_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.dutycycle_eena_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_1\ : std_logic;
signal \POWERLED.dutycycle_eena_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_0\ : std_logic;
signal \POWERLED.func_state_RNISKPU6Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_1_13\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_off_1_14\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_96_0_a3_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_0\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_cascade_\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI765BZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI886BZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4AZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNICGABZ0Z1\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCBZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \POWERLED.N_115_f0_1\ : std_logic;
signal \POWERLED.N_366_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI2O4A1Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI2O4A1_2Z0Z_2\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_5\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI68EU3Z0Z_1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_0_1_5_cascade_\ : std_logic;
signal \SUSWARN_N_fast\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.m18_e_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_c_RNI919HZ0Z1\ : std_logic;
signal \POWERLED.dutycycle_1_0_5_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIT69J5Z0Z_1\ : std_logic;
signal \G_155_cascade_\ : std_logic;
signal \POWERLED.N_73\ : std_logic;
signal \POWERLED.dutycycle_eena_1\ : std_logic;
signal \POWERLED.N_73_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \POWERLED.N_277\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_2\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7_cascade_\ : std_logic;
signal \POWERLED.un85_clk_100khz_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2078\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_0\ : std_logic;
signal \G_9\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_13\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \POWERLED.count_off_RNIBQDB2Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.count_offZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_10\ : std_logic;
signal \POWERLED.un34_clk_100khz_8\ : std_logic;
signal \POWERLED.un34_clk_100khz_9_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\ : std_logic;
signal \POWERLED.N_220_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823\ : std_logic;
signal \POWERLED.N_304_cascade_\ : std_logic;
signal \POWERLED.N_2216_i_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_1_cascade_\ : std_logic;
signal \POWERLED.N_160\ : std_logic;
signal \POWERLED.N_3_0\ : std_logic;
signal \slp_s3n_signal_cascade_\ : std_logic;
signal \POWERLED.N_183\ : std_logic;
signal \POWERLED.func_state_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_162_i\ : std_logic;
signal \POWERLED.N_335\ : std_logic;
signal \POWERLED.func_state_RNI2O4A1Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.dutycycle_en_9\ : std_logic;
signal \POWERLED.func_state_RNI2O4A1_1Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_42_and_i_0_0\ : std_logic;
signal \POWERLED.func_state_RNI2O4A1Z0Z_1\ : std_logic;
signal \POWERLED.un1_clk_100khz_47_and_i_0_0_cascade_\ : std_logic;
signal \POWERLED.N_399_N\ : std_logic;
signal \POWERLED.dutycycle_en_11\ : std_logic;
signal \POWERLED.m18_e_5\ : std_logic;
signal \POWERLED.m18_e_6\ : std_logic;
signal \POWERLED.func_m2_0_a2Z0Z_0\ : std_logic;
signal \POWERLED.func_m2_0_a2Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNI2O4A1_0Z0Z_10\ : std_logic;
signal \POWERLED.func_state_RNI91IA4_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_0\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \POWERLED.func_state_1_m2_0_cascade_\ : std_logic;
signal \POWERLED.g0_9_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_fb_15_4_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_fb_15_0\ : std_logic;
signal \POWERLED.dutycycle_en_14_cascade_\ : std_logic;
signal \POWERLED.func_m2_0_a2_isoZ0\ : std_logic;
signal \POWERLED.dutycycle_eena_14_0Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_fb_15_1\ : std_logic;
signal \POWERLED.g1_0\ : std_logic;
signal \POWERLED.g1\ : std_logic;
signal \POWERLED.dutycycle_fb_15_2_0\ : std_logic;
signal \SUSWARN_N_rep1\ : std_logic;
signal \POWERLED.N_340_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIRAVV2Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_5\ : std_logic;
signal \POWERLED.dutycycle_fb_15_1_1\ : std_logic;
signal \POWERLED.g2_0\ : std_logic;
signal \POWERLED.N_398_0\ : std_logic;
signal \POWERLED.g0_1_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_10\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_a3_0\ : std_logic;
signal \POWERLED.dutycycle_0_5\ : std_logic;
signal \POWERLED.dutycycle_fb_14_a4_1\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.count_off_1_sqmuxa\ : std_logic;
signal \POWERLED.count_off_1_sqmuxa_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_6\ : std_logic;
signal \POWERLED.N_325\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNINH5P1Z0Z_2\ : std_logic;
signal \POWERLED.dutycycle_RNI4G9K2Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNO_2Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.N_240\ : std_logic;
signal \POWERLED.dutycycle_eena_13\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0\ : std_logic;
signal \POWERLED.g3\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m3_1_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNO_3Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_6\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m3s4_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_6\ : std_logic;
signal \POWERLED.N_239\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.N_271\ : std_logic;
signal \POWERLED.N_366\ : std_logic;
signal \POWERLED.N_331\ : std_logic;
signal \POWERLED.N_272\ : std_logic;
signal \POWERLED.dutycycle_N_3_mux_0_0\ : std_logic;
signal \PCH_PWRGD.count_rst_10\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \PCH_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_1_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_0_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_2_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_11_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \N_253_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.count_RNIM6A821Z0Z_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2173_i\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_11_0\ : std_logic;
signal \PCH_PWRGD.N_2173_i_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.m4_0_a2_11_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.m4_0_a2_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.m4_0_a2_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.m4_0_a2_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.m4_0_a2_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_10_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0\ : std_logic;
signal \PCH_PWRGD.curr_state_0_0\ : std_logic;
signal \PCH_PWRGD.m4_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_8_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2_1_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_10\ : std_logic;
signal v33a_ok : std_logic;
signal v5a_ok : std_logic;
signal slp_susn : std_logic;
signal v1p8a_ok : std_logic;
signal \rsmrst_pwrgd_signal_cascade_\ : std_logic;
signal \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\ : std_logic;
signal \N_382\ : std_logic;
signal \RSMRST_PWRGD.N_254_i\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD_curr_state_0\ : std_logic;
signal \POWERLED.N_301\ : std_logic;
signal \G_11\ : std_logic;
signal \RSMRST_PWRGD.N_29_2\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_N_3_mux_0\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_1_5\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_off_0_6\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.count_off_0_2\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.func_state_RNISKPU6Z0Z_0\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_15\ : std_logic;
signal \RSMRSTn_rep1\ : std_logic;
signal \POWERLED.N_4_0_3\ : std_logic;
signal \POWERLED.func_state_RNIOGRSZ0Z_0\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o2_1\ : std_logic;
signal \POWERLED.N_76\ : std_logic;
signal \POWERLED.func_state_RNI91IA4Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_1\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.func_state_1_m2_1_cascade_\ : std_logic;
signal \POWERLED.func_state_enZ0\ : std_logic;
signal \POWERLED.un1_N_3_mux_0\ : std_logic;
signal \N_4_1_cascade_\ : std_logic;
signal \G_34_0_a4_0_2_cascade_\ : std_logic;
signal \POWERLED_un1_dutycycle_172_m3_0_0\ : std_logic;
signal \POWERLED.N_8_0\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1_ns_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_10Z0Z_3\ : std_logic;
signal \N_11\ : std_logic;
signal \POWERLED.N_319_0\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.N_297\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_a2_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_296_N_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_1_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_2\ : std_logic;
signal \POWERLED.N_340\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_\ : std_logic;
signal \POWERLED.N_284\ : std_logic;
signal \POWERLED.func_state_RNIBQDB2Z0Z_0\ : std_logic;
signal \POWERLED.N_340_N\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_0\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_294_N\ : std_logic;
signal \POWERLED.func_state_1_m2_am_1_1\ : std_logic;
signal \POWERLED.func_N_5_mux_0\ : std_logic;
signal \POWERLED.func_state_RNIBL3Q3Z0Z_1\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_a2_0_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \func_state_RNI_7_1\ : std_logic;
signal \N_7\ : std_logic;
signal rsmrstn : std_logic;
signal \POWERLED.func_state_RNIZ0Z_1\ : std_logic;
signal slp_s3n : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_a2_6_0_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_a2_6_sx_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIPUGO_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_309_N\ : std_logic;
signal \POWERLED.count_clk_RNI2O4A1Z0Z_10\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_o2_4_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.N_145_N\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_a2_5_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_a2_5_0_cascade_\ : std_logic;
signal \RSMRSTn_fast\ : std_logic;
signal \POWERLED.func_state_RNIPUGOZ0Z_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \PCH_PWRGD.count_rst_13_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_6_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_3_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_12_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_5\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_4_0\ : std_logic;
signal \PCH_PWRGD.count_rst_7\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_5_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_7\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\ : std_logic;
signal \PCH_PWRGD.N_364\ : std_logic;
signal \G_1939_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \N_218\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \G_1939\ : std_logic;
signal \N_218_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2190_i\ : std_logic;
signal \PCH_PWRGD.N_2171_i\ : std_logic;
signal \PCH_PWRGD.N_2190_i_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.N_53_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_1\ : std_logic;
signal \VPP_VDDQ.N_55_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_2\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_1_7_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_7_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_14_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.count_clk_0_14\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_1\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_1\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_a2_0_0_cascade_\ : std_logic;
signal \POWERLED.N_285\ : std_logic;
signal \POWERLED.N_177\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_1_cascade_\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal slp_s4n : std_logic;
signal \POWERLED.un1_func_state25_4_i_a2_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIBVNSZ0Z_0\ : std_logic;
signal \POWERLED.N_291\ : std_logic;
signal \POWERLED.count_clk_en_0_cascade_\ : std_logic;
signal \POWERLED.N_396\ : std_logic;
signal \POWERLED.func_state_RNI2O4A1_1Z0Z_1\ : std_logic;
signal \POWERLED.count_clk_en_2_cascade_\ : std_logic;
signal \G_155\ : std_logic;
signal \POWERLED.func_state_RNI_2Z0Z_1\ : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.N_176\ : std_logic;
signal \POWERLED.N_176_cascade_\ : std_logic;
signal \POWERLED.N_2218_i\ : std_logic;
signal \POWERLED.N_2216_i\ : std_logic;
signal \POWERLED.N_27\ : std_logic;
signal \POWERLED.func_state\ : std_logic;
signal \POWERLED.N_219\ : std_logic;
signal vpp_en : std_logic;
signal \VPP_VDDQ.N_64_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ.curr_state_7_0\ : std_logic;
signal \VPP_VDDQ.curr_state_7_0_cascade_\ : std_logic;
signal \N_246\ : std_logic;
signal \N_246_cascade_\ : std_logic;
signal \N_381\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal vccst_en : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_0\ : std_logic;
signal \VPP_VDDQ.un6_count_10_cascade_\ : std_logic;
signal \VPP_VDDQ_un6_count\ : std_logic;
signal \VPP_VDDQ.un6_count_8\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal suswarn_n : std_logic;
signal \VPP_VDDQ.N_361_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_62_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en_cascade_\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_ok\ : std_logic;
signal vddq_ok : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ.N_361_0\ : std_logic;
signal \N_570_g\ : std_logic;
signal \VPP_VDDQ.N_2192_i\ : std_logic;
signal \VPP_VDDQ.N_62\ : std_logic;
signal \VPP_VDDQ.N_62_i\ : std_logic;
signal \VPP_VDDQ.count_2_1_14_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_4_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_0_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_0_5\ : std_logic;
signal \VPP_VDDQ.count_2_1_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_174\ : std_logic;
signal dsw_pwrok : std_logic;
signal vccst_cpu_ok : std_logic;
signal v5s_ok : std_logic;
signal v33s_ok : std_logic;
signal slp_s3n_signal : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\ : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal vccin_en : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_9\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_0_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\ : std_logic;
signal \VPP_VDDQ.N_1_i_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.count_2_1_11_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.count_clkZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.count_clk_0_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.count_clkZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_cascade_\ : std_logic;
signal \POWERLED.N_352\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.un2_count_clk_15_0_9_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_15_0_8\ : std_logic;
signal \POWERLED.un2_count_clk_15_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.un2_count_clk_15_0_10\ : std_logic;
signal \POWERLED.count_clk_0_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_12_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_12_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_15_0_7\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_15\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1\ : std_logic;
signal \POWERLED.func_state_RNIH9594_0_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.count_clk_en\ : std_logic;
signal \VPP_VDDQ.N_66_i\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \N_29_g\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal fpga_osc : std_logic;
signal \VPP_VDDQ.N_29_0\ : std_logic;
signal \G_43\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    SLP_S0n <= \SLP_S0n_wire\;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35432\,
            DIN => \N__35431\,
            DOUT => \N__35430\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35432\,
            PADOUT => \N__35431\,
            PADIN => \N__35430\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35423\,
            DIN => \N__35422\,
            DOUT => \N__35421\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35423\,
            PADOUT => \N__35422\,
            PADIN => \N__35421\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16753\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35414\,
            DIN => \N__35413\,
            DOUT => \N__35412\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35414\,
            PADOUT => \N__35413\,
            PADIN => \N__35412\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24942\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35405\,
            DIN => \N__35404\,
            DOUT => \N__35403\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35405\,
            PADOUT => \N__35404\,
            PADIN => \N__35403\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17059\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35396\,
            DIN => \N__35395\,
            DOUT => \N__35394\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35396\,
            PADOUT => \N__35395\,
            PADIN => \N__35394\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35387\,
            DIN => \N__35386\,
            DOUT => \N__35385\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35387\,
            PADOUT => \N__35386\,
            PADIN => \N__35385\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35378\,
            DIN => \N__35377\,
            DOUT => \N__35376\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35378\,
            PADOUT => \N__35377\,
            PADIN => \N__35376\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35369\,
            DIN => \N__35368\,
            DOUT => \N__35367\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35369\,
            PADOUT => \N__35368\,
            PADIN => \N__35367\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35360\,
            DIN => \N__35359\,
            DOUT => \N__35358\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35360\,
            PADOUT => \N__35359\,
            PADIN => \N__35358\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16791\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35351\,
            DIN => \N__35350\,
            DOUT => \N__35349\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35351\,
            PADOUT => \N__35350\,
            PADIN => \N__35349\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35342\,
            DIN => \N__35341\,
            DOUT => \N__35340\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35342\,
            PADOUT => \N__35341\,
            PADIN => \N__35340\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35333\,
            DIN => \N__35332\,
            DOUT => \N__35331\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35333\,
            PADOUT => \N__35332\,
            PADIN => \N__35331\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14140\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35324\,
            DIN => \N__35323\,
            DOUT => \N__35322\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35324\,
            PADOUT => \N__35323\,
            PADIN => \N__35322\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35315\,
            DIN => \N__35314\,
            DOUT => \N__35313\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35315\,
            PADOUT => \N__35314\,
            PADIN => \N__35313\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35306\,
            DIN => \N__35305\,
            DOUT => \N__35304\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35306\,
            PADOUT => \N__35305\,
            PADIN => \N__35304\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35297\,
            DIN => \N__35296\,
            DOUT => \N__35295\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35297\,
            PADOUT => \N__35296\,
            PADIN => \N__35295\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35288\,
            DIN => \N__35287\,
            DOUT => \N__35286\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35288\,
            PADOUT => \N__35287\,
            PADIN => \N__35286\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30212\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35279\,
            DIN => \N__35278\,
            DOUT => \N__35277\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35279\,
            PADOUT => \N__35278\,
            PADIN => \N__35277\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35270\,
            DIN => \N__35269\,
            DOUT => \N__35268\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35270\,
            PADOUT => \N__35269\,
            PADIN => \N__35268\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35261\,
            DIN => \N__35260\,
            DOUT => \N__35259\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35261\,
            PADOUT => \N__35260\,
            PADIN => \N__35259\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30637\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35252\,
            DIN => \N__35251\,
            DOUT => \N__35250\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35252\,
            PADOUT => \N__35251\,
            PADIN => \N__35250\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35243\,
            DIN => \N__35242\,
            DOUT => \N__35241\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35243\,
            PADOUT => \N__35242\,
            PADIN => \N__35241\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35234\,
            DIN => \N__35233\,
            DOUT => \N__35232\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35234\,
            PADOUT => \N__35233\,
            PADIN => \N__35232\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35225\,
            DIN => \N__35224\,
            DOUT => \N__35223\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35225\,
            PADOUT => \N__35224\,
            PADIN => \N__35223\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35216\,
            DIN => \N__35215\,
            DOUT => \N__35214\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35216\,
            PADOUT => \N__35215\,
            PADIN => \N__35214\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26413\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35207\,
            DIN => \N__35206\,
            DOUT => \N__35205\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35207\,
            PADOUT => \N__35206\,
            PADIN => \N__35205\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35198\,
            DIN => \N__35197\,
            DOUT => \N__35196\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35198\,
            PADOUT => \N__35197\,
            PADIN => \N__35196\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18721\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35189\,
            DIN => \N__35188\,
            DOUT => \N__35187\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35189\,
            PADOUT => \N__35188\,
            PADIN => \N__35187\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18781\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35180\,
            DIN => \N__35179\,
            DOUT => \N__35178\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35180\,
            PADOUT => \N__35179\,
            PADIN => \N__35178\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35171\,
            DIN => \N__35170\,
            DOUT => \N__35169\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35171\,
            PADOUT => \N__35170\,
            PADIN => \N__35169\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35162\,
            DIN => \N__35161\,
            DOUT => \N__35160\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35162\,
            PADOUT => \N__35161\,
            PADIN => \N__35160\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35153\,
            DIN => \N__35152\,
            DOUT => \N__35151\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35153\,
            PADOUT => \N__35152\,
            PADIN => \N__35151\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35144\,
            DIN => \N__35143\,
            DOUT => \N__35142\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35144\,
            PADOUT => \N__35143\,
            PADIN => \N__35142\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34566\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35135\,
            DIN => \N__35134\,
            DOUT => \N__35133\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35135\,
            PADOUT => \N__35134\,
            PADIN => \N__35133\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14665\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35126\,
            DIN => \N__35125\,
            DOUT => \N__35124\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35126\,
            PADOUT => \N__35125\,
            PADIN => \N__35124\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35117\,
            DIN => \N__35116\,
            DOUT => \N__35115\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35117\,
            PADOUT => \N__35116\,
            PADIN => \N__35115\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29143\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35108\,
            DIN => \N__35107\,
            DOUT => \N__35106\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35108\,
            PADOUT => \N__35107\,
            PADIN => \N__35106\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35099\,
            DIN => \N__35098\,
            DOUT => \N__35097\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35099\,
            PADOUT => \N__35098\,
            PADIN => \N__35097\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35090\,
            DIN => \N__35089\,
            DOUT => \N__35088\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35090\,
            PADOUT => \N__35089\,
            PADIN => \N__35088\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35081\,
            DIN => \N__35080\,
            DOUT => \N__35079\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35081\,
            PADOUT => \N__35080\,
            PADIN => \N__35079\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35072\,
            DIN => \N__35071\,
            DOUT => \N__35070\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35072\,
            PADOUT => \N__35071\,
            PADIN => \N__35070\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24859\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35063\,
            DIN => \N__35062\,
            DOUT => \N__35061\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35063\,
            PADOUT => \N__35062\,
            PADIN => \N__35061\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35054\,
            DIN => \N__35053\,
            DOUT => \N__35052\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35054\,
            PADOUT => \N__35053\,
            PADIN => \N__35052\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16795\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35045\,
            DIN => \N__35044\,
            DOUT => \N__35043\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35045\,
            PADOUT => \N__35044\,
            PADIN => \N__35043\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35036\,
            DIN => \N__35035\,
            DOUT => \N__35034\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35036\,
            PADOUT => \N__35035\,
            PADIN => \N__35034\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31237\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35027\,
            DIN => \N__35026\,
            DOUT => \N__35025\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35027\,
            PADOUT => \N__35026\,
            PADIN => \N__35025\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24949\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35018\,
            DIN => \N__35017\,
            DOUT => \N__35016\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35018\,
            PADOUT => \N__35017\,
            PADIN => \N__35016\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35009\,
            DIN => \N__35008\,
            DOUT => \N__35007\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35009\,
            PADOUT => \N__35008\,
            PADIN => \N__35007\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35000\,
            DIN => \N__34999\,
            DOUT => \N__34998\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35000\,
            PADOUT => \N__34999\,
            PADIN => \N__34998\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34991\,
            DIN => \N__34990\,
            DOUT => \N__34989\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34991\,
            PADOUT => \N__34990\,
            PADIN => \N__34989\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34982\,
            DIN => \N__34981\,
            DOUT => \N__34980\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34982\,
            PADOUT => \N__34981\,
            PADIN => \N__34980\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30916\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34973\,
            DIN => \N__34972\,
            DOUT => \N__34971\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34973\,
            PADOUT => \N__34972\,
            PADIN => \N__34971\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34964\,
            DIN => \N__34963\,
            DOUT => \N__34962\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34964\,
            PADOUT => \N__34963\,
            PADIN => \N__34962\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34955\,
            DIN => \N__34954\,
            DOUT => \N__34953\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34955\,
            PADOUT => \N__34954\,
            PADIN => \N__34953\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34946\,
            DIN => \N__34945\,
            DOUT => \N__34944\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34946\,
            PADOUT => \N__34945\,
            PADIN => \N__34944\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34937\,
            DIN => \N__34936\,
            DOUT => \N__34935\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34937\,
            PADOUT => \N__34936\,
            PADIN => \N__34935\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34928\,
            DIN => \N__34927\,
            DOUT => \N__34926\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34928\,
            PADOUT => \N__34927\,
            PADIN => \N__34926\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34919\,
            DIN => \N__34918\,
            DOUT => \N__34917\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34919\,
            PADOUT => \N__34918\,
            PADIN => \N__34917\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18771\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34910\,
            DIN => \N__34909\,
            DOUT => \N__34908\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34910\,
            PADOUT => \N__34909\,
            PADIN => \N__34908\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__8159\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34830\
        );

    \I__8158\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34830\
        );

    \I__8157\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34830\
        );

    \I__8156\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34830\
        );

    \I__8155\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34821\
        );

    \I__8154\ : InMux
    port map (
            O => \N__34886\,
            I => \N__34821\
        );

    \I__8153\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34821\
        );

    \I__8152\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34821\
        );

    \I__8151\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34812\
        );

    \I__8150\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34812\
        );

    \I__8149\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34812\
        );

    \I__8148\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34812\
        );

    \I__8147\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34805\
        );

    \I__8146\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34805\
        );

    \I__8145\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34805\
        );

    \I__8144\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34798\
        );

    \I__8143\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34798\
        );

    \I__8142\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34798\
        );

    \I__8141\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34789\
        );

    \I__8140\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34789\
        );

    \I__8139\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34789\
        );

    \I__8138\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34789\
        );

    \I__8137\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34780\
        );

    \I__8136\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34780\
        );

    \I__8135\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34780\
        );

    \I__8134\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34780\
        );

    \I__8133\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34771\
        );

    \I__8132\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34771\
        );

    \I__8131\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34771\
        );

    \I__8130\ : InMux
    port map (
            O => \N__34862\,
            I => \N__34771\
        );

    \I__8129\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34762\
        );

    \I__8128\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34762\
        );

    \I__8127\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34762\
        );

    \I__8126\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34762\
        );

    \I__8125\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34759\
        );

    \I__8124\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34754\
        );

    \I__8123\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34754\
        );

    \I__8122\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34745\
        );

    \I__8121\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34745\
        );

    \I__8120\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34745\
        );

    \I__8119\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34745\
        );

    \I__8118\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34736\
        );

    \I__8117\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34736\
        );

    \I__8116\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34736\
        );

    \I__8115\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34736\
        );

    \I__8114\ : InMux
    port map (
            O => \N__34846\,
            I => \N__34729\
        );

    \I__8113\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34729\
        );

    \I__8112\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34729\
        );

    \I__8111\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34726\
        );

    \I__8110\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34721\
        );

    \I__8109\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34721\
        );

    \I__8108\ : InMux
    port map (
            O => \N__34840\,
            I => \N__34718\
        );

    \I__8107\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34715\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__34830\,
            I => \N__34707\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__34821\,
            I => \N__34703\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__34812\,
            I => \N__34700\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__34805\,
            I => \N__34697\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__34798\,
            I => \N__34693\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__34789\,
            I => \N__34690\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__34780\,
            I => \N__34684\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34681\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34678\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__34759\,
            I => \N__34675\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34672\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__34745\,
            I => \N__34669\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34666\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__34729\,
            I => \N__34663\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__34726\,
            I => \N__34660\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34657\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__34718\,
            I => \N__34654\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__34715\,
            I => \N__34651\
        );

    \I__8088\ : CEMux
    port map (
            O => \N__34714\,
            I => \N__34594\
        );

    \I__8087\ : CEMux
    port map (
            O => \N__34713\,
            I => \N__34594\
        );

    \I__8086\ : CEMux
    port map (
            O => \N__34712\,
            I => \N__34594\
        );

    \I__8085\ : CEMux
    port map (
            O => \N__34711\,
            I => \N__34594\
        );

    \I__8084\ : CEMux
    port map (
            O => \N__34710\,
            I => \N__34594\
        );

    \I__8083\ : Glb2LocalMux
    port map (
            O => \N__34707\,
            I => \N__34594\
        );

    \I__8082\ : CEMux
    port map (
            O => \N__34706\,
            I => \N__34594\
        );

    \I__8081\ : Glb2LocalMux
    port map (
            O => \N__34703\,
            I => \N__34594\
        );

    \I__8080\ : Glb2LocalMux
    port map (
            O => \N__34700\,
            I => \N__34594\
        );

    \I__8079\ : Glb2LocalMux
    port map (
            O => \N__34697\,
            I => \N__34594\
        );

    \I__8078\ : CEMux
    port map (
            O => \N__34696\,
            I => \N__34594\
        );

    \I__8077\ : Glb2LocalMux
    port map (
            O => \N__34693\,
            I => \N__34594\
        );

    \I__8076\ : Glb2LocalMux
    port map (
            O => \N__34690\,
            I => \N__34594\
        );

    \I__8075\ : CEMux
    port map (
            O => \N__34689\,
            I => \N__34594\
        );

    \I__8074\ : CEMux
    port map (
            O => \N__34688\,
            I => \N__34594\
        );

    \I__8073\ : CEMux
    port map (
            O => \N__34687\,
            I => \N__34594\
        );

    \I__8072\ : Glb2LocalMux
    port map (
            O => \N__34684\,
            I => \N__34594\
        );

    \I__8071\ : Glb2LocalMux
    port map (
            O => \N__34681\,
            I => \N__34594\
        );

    \I__8070\ : Glb2LocalMux
    port map (
            O => \N__34678\,
            I => \N__34594\
        );

    \I__8069\ : Glb2LocalMux
    port map (
            O => \N__34675\,
            I => \N__34594\
        );

    \I__8068\ : Glb2LocalMux
    port map (
            O => \N__34672\,
            I => \N__34594\
        );

    \I__8067\ : Glb2LocalMux
    port map (
            O => \N__34669\,
            I => \N__34594\
        );

    \I__8066\ : Glb2LocalMux
    port map (
            O => \N__34666\,
            I => \N__34594\
        );

    \I__8065\ : Glb2LocalMux
    port map (
            O => \N__34663\,
            I => \N__34594\
        );

    \I__8064\ : Glb2LocalMux
    port map (
            O => \N__34660\,
            I => \N__34594\
        );

    \I__8063\ : Glb2LocalMux
    port map (
            O => \N__34657\,
            I => \N__34594\
        );

    \I__8062\ : Glb2LocalMux
    port map (
            O => \N__34654\,
            I => \N__34594\
        );

    \I__8061\ : Glb2LocalMux
    port map (
            O => \N__34651\,
            I => \N__34594\
        );

    \I__8060\ : GlobalMux
    port map (
            O => \N__34594\,
            I => \N__34591\
        );

    \I__8059\ : gio2CtrlBuf
    port map (
            O => \N__34591\,
            I => \N_29_g\
        );

    \I__8058\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34584\
        );

    \I__8057\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34581\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__34584\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__34581\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__8054\ : InMux
    port map (
            O => \N__34576\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__8053\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__8051\ : Span4Mux_s3_v
    port map (
            O => \N__34567\,
            I => \N__34562\
        );

    \I__8050\ : IoInMux
    port map (
            O => \N__34566\,
            I => \N__34558\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34553\
        );

    \I__8048\ : Span4Mux_h
    port map (
            O => \N__34562\,
            I => \N__34550\
        );

    \I__8047\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34547\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34544\
        );

    \I__8045\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34541\
        );

    \I__8044\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34538\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__34553\,
            I => \N__34534\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__34550\,
            I => \N__34529\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34529\
        );

    \I__8040\ : Span4Mux_s3_h
    port map (
            O => \N__34544\,
            I => \N__34526\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34523\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34520\
        );

    \I__8037\ : InMux
    port map (
            O => \N__34537\,
            I => \N__34517\
        );

    \I__8036\ : Span4Mux_v
    port map (
            O => \N__34534\,
            I => \N__34514\
        );

    \I__8035\ : Span4Mux_v
    port map (
            O => \N__34529\,
            I => \N__34511\
        );

    \I__8034\ : Span4Mux_v
    port map (
            O => \N__34526\,
            I => \N__34506\
        );

    \I__8033\ : Span4Mux_v
    port map (
            O => \N__34523\,
            I => \N__34506\
        );

    \I__8032\ : Span4Mux_v
    port map (
            O => \N__34520\,
            I => \N__34501\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__34517\,
            I => \N__34501\
        );

    \I__8030\ : Span4Mux_h
    port map (
            O => \N__34514\,
            I => \N__34497\
        );

    \I__8029\ : Span4Mux_v
    port map (
            O => \N__34511\,
            I => \N__34494\
        );

    \I__8028\ : Span4Mux_h
    port map (
            O => \N__34506\,
            I => \N__34489\
        );

    \I__8027\ : Span4Mux_v
    port map (
            O => \N__34501\,
            I => \N__34489\
        );

    \I__8026\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34486\
        );

    \I__8025\ : Odrv4
    port map (
            O => \N__34497\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__34494\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__34489\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__34486\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8021\ : InMux
    port map (
            O => \N__34477\,
            I => \bfn_12_16_0_\
        );

    \I__8020\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34470\
        );

    \I__8019\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34467\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__34470\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__34467\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__8016\ : ClkMux
    port map (
            O => \N__34462\,
            I => \N__34455\
        );

    \I__8015\ : ClkMux
    port map (
            O => \N__34461\,
            I => \N__34452\
        );

    \I__8014\ : ClkMux
    port map (
            O => \N__34460\,
            I => \N__34446\
        );

    \I__8013\ : ClkMux
    port map (
            O => \N__34459\,
            I => \N__34441\
        );

    \I__8012\ : ClkMux
    port map (
            O => \N__34458\,
            I => \N__34435\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__34455\,
            I => \N__34426\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__34452\,
            I => \N__34422\
        );

    \I__8009\ : ClkMux
    port map (
            O => \N__34451\,
            I => \N__34418\
        );

    \I__8008\ : ClkMux
    port map (
            O => \N__34450\,
            I => \N__34413\
        );

    \I__8007\ : ClkMux
    port map (
            O => \N__34449\,
            I => \N__34409\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__34446\,
            I => \N__34406\
        );

    \I__8005\ : ClkMux
    port map (
            O => \N__34445\,
            I => \N__34403\
        );

    \I__8004\ : ClkMux
    port map (
            O => \N__34444\,
            I => \N__34400\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34397\
        );

    \I__8002\ : ClkMux
    port map (
            O => \N__34440\,
            I => \N__34394\
        );

    \I__8001\ : ClkMux
    port map (
            O => \N__34439\,
            I => \N__34391\
        );

    \I__8000\ : ClkMux
    port map (
            O => \N__34438\,
            I => \N__34385\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__34435\,
            I => \N__34382\
        );

    \I__7998\ : ClkMux
    port map (
            O => \N__34434\,
            I => \N__34379\
        );

    \I__7997\ : ClkMux
    port map (
            O => \N__34433\,
            I => \N__34375\
        );

    \I__7996\ : ClkMux
    port map (
            O => \N__34432\,
            I => \N__34369\
        );

    \I__7995\ : ClkMux
    port map (
            O => \N__34431\,
            I => \N__34365\
        );

    \I__7994\ : ClkMux
    port map (
            O => \N__34430\,
            I => \N__34362\
        );

    \I__7993\ : ClkMux
    port map (
            O => \N__34429\,
            I => \N__34358\
        );

    \I__7992\ : Span4Mux_s1_h
    port map (
            O => \N__34426\,
            I => \N__34354\
        );

    \I__7991\ : ClkMux
    port map (
            O => \N__34425\,
            I => \N__34351\
        );

    \I__7990\ : Span4Mux_s1_h
    port map (
            O => \N__34422\,
            I => \N__34345\
        );

    \I__7989\ : ClkMux
    port map (
            O => \N__34421\,
            I => \N__34342\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__34418\,
            I => \N__34339\
        );

    \I__7987\ : ClkMux
    port map (
            O => \N__34417\,
            I => \N__34336\
        );

    \I__7986\ : ClkMux
    port map (
            O => \N__34416\,
            I => \N__34333\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__34413\,
            I => \N__34329\
        );

    \I__7984\ : ClkMux
    port map (
            O => \N__34412\,
            I => \N__34325\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34318\
        );

    \I__7982\ : Span4Mux_v
    port map (
            O => \N__34406\,
            I => \N__34311\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34311\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__34400\,
            I => \N__34311\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__34397\,
            I => \N__34304\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__34394\,
            I => \N__34304\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34304\
        );

    \I__7976\ : ClkMux
    port map (
            O => \N__34390\,
            I => \N__34301\
        );

    \I__7975\ : ClkMux
    port map (
            O => \N__34389\,
            I => \N__34298\
        );

    \I__7974\ : ClkMux
    port map (
            O => \N__34388\,
            I => \N__34295\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__34385\,
            I => \N__34285\
        );

    \I__7972\ : Span4Mux_h
    port map (
            O => \N__34382\,
            I => \N__34285\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__34379\,
            I => \N__34285\
        );

    \I__7970\ : ClkMux
    port map (
            O => \N__34378\,
            I => \N__34282\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__34375\,
            I => \N__34279\
        );

    \I__7968\ : ClkMux
    port map (
            O => \N__34374\,
            I => \N__34276\
        );

    \I__7967\ : ClkMux
    port map (
            O => \N__34373\,
            I => \N__34272\
        );

    \I__7966\ : ClkMux
    port map (
            O => \N__34372\,
            I => \N__34268\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__34369\,
            I => \N__34264\
        );

    \I__7964\ : ClkMux
    port map (
            O => \N__34368\,
            I => \N__34261\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__34365\,
            I => \N__34258\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__34362\,
            I => \N__34255\
        );

    \I__7961\ : ClkMux
    port map (
            O => \N__34361\,
            I => \N__34252\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__34358\,
            I => \N__34249\
        );

    \I__7959\ : ClkMux
    port map (
            O => \N__34357\,
            I => \N__34246\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__34354\,
            I => \N__34241\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__34351\,
            I => \N__34241\
        );

    \I__7956\ : ClkMux
    port map (
            O => \N__34350\,
            I => \N__34237\
        );

    \I__7955\ : ClkMux
    port map (
            O => \N__34349\,
            I => \N__34234\
        );

    \I__7954\ : ClkMux
    port map (
            O => \N__34348\,
            I => \N__34230\
        );

    \I__7953\ : Span4Mux_v
    port map (
            O => \N__34345\,
            I => \N__34225\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34225\
        );

    \I__7951\ : Span4Mux_s2_h
    port map (
            O => \N__34339\,
            I => \N__34217\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__34336\,
            I => \N__34217\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__34333\,
            I => \N__34214\
        );

    \I__7948\ : ClkMux
    port map (
            O => \N__34332\,
            I => \N__34211\
        );

    \I__7947\ : Span4Mux_s2_h
    port map (
            O => \N__34329\,
            I => \N__34207\
        );

    \I__7946\ : ClkMux
    port map (
            O => \N__34328\,
            I => \N__34204\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__34325\,
            I => \N__34201\
        );

    \I__7944\ : ClkMux
    port map (
            O => \N__34324\,
            I => \N__34198\
        );

    \I__7943\ : ClkMux
    port map (
            O => \N__34323\,
            I => \N__34192\
        );

    \I__7942\ : ClkMux
    port map (
            O => \N__34322\,
            I => \N__34189\
        );

    \I__7941\ : ClkMux
    port map (
            O => \N__34321\,
            I => \N__34186\
        );

    \I__7940\ : Span4Mux_h
    port map (
            O => \N__34318\,
            I => \N__34182\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__34311\,
            I => \N__34171\
        );

    \I__7938\ : Span4Mux_v
    port map (
            O => \N__34304\,
            I => \N__34171\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__34301\,
            I => \N__34171\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__34298\,
            I => \N__34171\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__34295\,
            I => \N__34171\
        );

    \I__7934\ : ClkMux
    port map (
            O => \N__34294\,
            I => \N__34167\
        );

    \I__7933\ : ClkMux
    port map (
            O => \N__34293\,
            I => \N__34164\
        );

    \I__7932\ : ClkMux
    port map (
            O => \N__34292\,
            I => \N__34158\
        );

    \I__7931\ : Span4Mux_v
    port map (
            O => \N__34285\,
            I => \N__34153\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__34282\,
            I => \N__34153\
        );

    \I__7929\ : Span4Mux_s1_h
    port map (
            O => \N__34279\,
            I => \N__34148\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34148\
        );

    \I__7927\ : ClkMux
    port map (
            O => \N__34275\,
            I => \N__34145\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__34272\,
            I => \N__34140\
        );

    \I__7925\ : ClkMux
    port map (
            O => \N__34271\,
            I => \N__34137\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__34268\,
            I => \N__34134\
        );

    \I__7923\ : ClkMux
    port map (
            O => \N__34267\,
            I => \N__34131\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__34264\,
            I => \N__34126\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34126\
        );

    \I__7920\ : Span4Mux_v
    port map (
            O => \N__34258\,
            I => \N__34119\
        );

    \I__7919\ : Span4Mux_s1_h
    port map (
            O => \N__34255\,
            I => \N__34119\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__34252\,
            I => \N__34119\
        );

    \I__7917\ : Span4Mux_s2_h
    port map (
            O => \N__34249\,
            I => \N__34114\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34114\
        );

    \I__7915\ : Span4Mux_h
    port map (
            O => \N__34241\,
            I => \N__34111\
        );

    \I__7914\ : ClkMux
    port map (
            O => \N__34240\,
            I => \N__34108\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__34237\,
            I => \N__34105\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__34234\,
            I => \N__34102\
        );

    \I__7911\ : ClkMux
    port map (
            O => \N__34233\,
            I => \N__34099\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34096\
        );

    \I__7909\ : Span4Mux_s1_h
    port map (
            O => \N__34225\,
            I => \N__34093\
        );

    \I__7908\ : ClkMux
    port map (
            O => \N__34224\,
            I => \N__34090\
        );

    \I__7907\ : ClkMux
    port map (
            O => \N__34223\,
            I => \N__34087\
        );

    \I__7906\ : ClkMux
    port map (
            O => \N__34222\,
            I => \N__34081\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__34217\,
            I => \N__34073\
        );

    \I__7904\ : Span4Mux_s2_h
    port map (
            O => \N__34214\,
            I => \N__34073\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__34211\,
            I => \N__34073\
        );

    \I__7902\ : ClkMux
    port map (
            O => \N__34210\,
            I => \N__34070\
        );

    \I__7901\ : Span4Mux_v
    port map (
            O => \N__34207\,
            I => \N__34064\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__34204\,
            I => \N__34064\
        );

    \I__7899\ : Span4Mux_s2_h
    port map (
            O => \N__34201\,
            I => \N__34059\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34059\
        );

    \I__7897\ : ClkMux
    port map (
            O => \N__34197\,
            I => \N__34056\
        );

    \I__7896\ : ClkMux
    port map (
            O => \N__34196\,
            I => \N__34052\
        );

    \I__7895\ : ClkMux
    port map (
            O => \N__34195\,
            I => \N__34049\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__34192\,
            I => \N__34046\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34041\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__34186\,
            I => \N__34041\
        );

    \I__7891\ : ClkMux
    port map (
            O => \N__34185\,
            I => \N__34038\
        );

    \I__7890\ : Span4Mux_v
    port map (
            O => \N__34182\,
            I => \N__34035\
        );

    \I__7889\ : Span4Mux_v
    port map (
            O => \N__34171\,
            I => \N__34032\
        );

    \I__7888\ : ClkMux
    port map (
            O => \N__34170\,
            I => \N__34029\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34024\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__34164\,
            I => \N__34024\
        );

    \I__7885\ : ClkMux
    port map (
            O => \N__34163\,
            I => \N__34021\
        );

    \I__7884\ : ClkMux
    port map (
            O => \N__34162\,
            I => \N__34017\
        );

    \I__7883\ : ClkMux
    port map (
            O => \N__34161\,
            I => \N__34014\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__34158\,
            I => \N__34010\
        );

    \I__7881\ : Span4Mux_v
    port map (
            O => \N__34153\,
            I => \N__34003\
        );

    \I__7880\ : Span4Mux_v
    port map (
            O => \N__34148\,
            I => \N__34003\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__34145\,
            I => \N__34003\
        );

    \I__7878\ : ClkMux
    port map (
            O => \N__34144\,
            I => \N__34000\
        );

    \I__7877\ : ClkMux
    port map (
            O => \N__34143\,
            I => \N__33993\
        );

    \I__7876\ : Span4Mux_s3_h
    port map (
            O => \N__34140\,
            I => \N__33984\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__33984\
        );

    \I__7874\ : Span4Mux_s3_h
    port map (
            O => \N__34134\,
            I => \N__33984\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__34131\,
            I => \N__33984\
        );

    \I__7872\ : Span4Mux_v
    port map (
            O => \N__34126\,
            I => \N__33980\
        );

    \I__7871\ : Span4Mux_h
    port map (
            O => \N__34119\,
            I => \N__33975\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__34114\,
            I => \N__33975\
        );

    \I__7869\ : Span4Mux_h
    port map (
            O => \N__34111\,
            I => \N__33970\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__34108\,
            I => \N__33970\
        );

    \I__7867\ : Span4Mux_s1_h
    port map (
            O => \N__34105\,
            I => \N__33963\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__34102\,
            I => \N__33963\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__33963\
        );

    \I__7864\ : Span4Mux_s1_h
    port map (
            O => \N__34096\,
            I => \N__33960\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__34093\,
            I => \N__33955\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__34090\,
            I => \N__33955\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__34087\,
            I => \N__33952\
        );

    \I__7860\ : ClkMux
    port map (
            O => \N__34086\,
            I => \N__33949\
        );

    \I__7859\ : ClkMux
    port map (
            O => \N__34085\,
            I => \N__33946\
        );

    \I__7858\ : ClkMux
    port map (
            O => \N__34084\,
            I => \N__33943\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__34081\,
            I => \N__33940\
        );

    \I__7856\ : ClkMux
    port map (
            O => \N__34080\,
            I => \N__33937\
        );

    \I__7855\ : Span4Mux_v
    port map (
            O => \N__34073\,
            I => \N__33932\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__34070\,
            I => \N__33932\
        );

    \I__7853\ : ClkMux
    port map (
            O => \N__34069\,
            I => \N__33929\
        );

    \I__7852\ : Span4Mux_v
    port map (
            O => \N__34064\,
            I => \N__33922\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__34059\,
            I => \N__33922\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__34056\,
            I => \N__33922\
        );

    \I__7849\ : ClkMux
    port map (
            O => \N__34055\,
            I => \N__33919\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__34052\,
            I => \N__33916\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__34049\,
            I => \N__33913\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__34046\,
            I => \N__33906\
        );

    \I__7845\ : Span4Mux_h
    port map (
            O => \N__34041\,
            I => \N__33906\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__33906\
        );

    \I__7843\ : Span4Mux_h
    port map (
            O => \N__34035\,
            I => \N__33895\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__34032\,
            I => \N__33895\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__33895\
        );

    \I__7840\ : Span4Mux_h
    port map (
            O => \N__34024\,
            I => \N__33895\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__34021\,
            I => \N__33895\
        );

    \I__7838\ : ClkMux
    port map (
            O => \N__34020\,
            I => \N__33892\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__34017\,
            I => \N__33889\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__34014\,
            I => \N__33886\
        );

    \I__7835\ : ClkMux
    port map (
            O => \N__34013\,
            I => \N__33883\
        );

    \I__7834\ : Span4Mux_s1_h
    port map (
            O => \N__34010\,
            I => \N__33876\
        );

    \I__7833\ : Span4Mux_s2_v
    port map (
            O => \N__34003\,
            I => \N__33876\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34000\,
            I => \N__33876\
        );

    \I__7831\ : ClkMux
    port map (
            O => \N__33999\,
            I => \N__33872\
        );

    \I__7830\ : ClkMux
    port map (
            O => \N__33998\,
            I => \N__33869\
        );

    \I__7829\ : ClkMux
    port map (
            O => \N__33997\,
            I => \N__33866\
        );

    \I__7828\ : ClkMux
    port map (
            O => \N__33996\,
            I => \N__33863\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33860\
        );

    \I__7826\ : Span4Mux_v
    port map (
            O => \N__33984\,
            I => \N__33857\
        );

    \I__7825\ : ClkMux
    port map (
            O => \N__33983\,
            I => \N__33854\
        );

    \I__7824\ : Span4Mux_v
    port map (
            O => \N__33980\,
            I => \N__33850\
        );

    \I__7823\ : Span4Mux_v
    port map (
            O => \N__33975\,
            I => \N__33843\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__33970\,
            I => \N__33843\
        );

    \I__7821\ : Span4Mux_h
    port map (
            O => \N__33963\,
            I => \N__33843\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__33960\,
            I => \N__33830\
        );

    \I__7819\ : Span4Mux_v
    port map (
            O => \N__33955\,
            I => \N__33830\
        );

    \I__7818\ : Span4Mux_h
    port map (
            O => \N__33952\,
            I => \N__33830\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__33949\,
            I => \N__33830\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33830\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__33943\,
            I => \N__33830\
        );

    \I__7814\ : Span4Mux_s1_h
    port map (
            O => \N__33940\,
            I => \N__33825\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__33937\,
            I => \N__33825\
        );

    \I__7812\ : Span4Mux_v
    port map (
            O => \N__33932\,
            I => \N__33820\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__33929\,
            I => \N__33820\
        );

    \I__7810\ : Span4Mux_v
    port map (
            O => \N__33922\,
            I => \N__33815\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__33919\,
            I => \N__33815\
        );

    \I__7808\ : Span4Mux_v
    port map (
            O => \N__33916\,
            I => \N__33804\
        );

    \I__7807\ : Span4Mux_h
    port map (
            O => \N__33913\,
            I => \N__33804\
        );

    \I__7806\ : IoSpan4Mux
    port map (
            O => \N__33906\,
            I => \N__33804\
        );

    \I__7805\ : Span4Mux_v
    port map (
            O => \N__33895\,
            I => \N__33804\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__33892\,
            I => \N__33804\
        );

    \I__7803\ : Span4Mux_v
    port map (
            O => \N__33889\,
            I => \N__33795\
        );

    \I__7802\ : Span4Mux_h
    port map (
            O => \N__33886\,
            I => \N__33795\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__33883\,
            I => \N__33795\
        );

    \I__7800\ : Span4Mux_h
    port map (
            O => \N__33876\,
            I => \N__33795\
        );

    \I__7799\ : ClkMux
    port map (
            O => \N__33875\,
            I => \N__33792\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__33872\,
            I => \N__33789\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__33869\,
            I => \N__33786\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__33866\,
            I => \N__33781\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__33863\,
            I => \N__33781\
        );

    \I__7794\ : Span12Mux_s5_h
    port map (
            O => \N__33860\,
            I => \N__33778\
        );

    \I__7793\ : Sp12to4
    port map (
            O => \N__33857\,
            I => \N__33775\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__33854\,
            I => \N__33772\
        );

    \I__7791\ : ClkMux
    port map (
            O => \N__33853\,
            I => \N__33769\
        );

    \I__7790\ : IoSpan4Mux
    port map (
            O => \N__33850\,
            I => \N__33766\
        );

    \I__7789\ : Span4Mux_v
    port map (
            O => \N__33843\,
            I => \N__33763\
        );

    \I__7788\ : Span4Mux_v
    port map (
            O => \N__33830\,
            I => \N__33758\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__33825\,
            I => \N__33758\
        );

    \I__7786\ : IoSpan4Mux
    port map (
            O => \N__33820\,
            I => \N__33751\
        );

    \I__7785\ : IoSpan4Mux
    port map (
            O => \N__33815\,
            I => \N__33751\
        );

    \I__7784\ : IoSpan4Mux
    port map (
            O => \N__33804\,
            I => \N__33751\
        );

    \I__7783\ : Span4Mux_v
    port map (
            O => \N__33795\,
            I => \N__33746\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__33792\,
            I => \N__33746\
        );

    \I__7781\ : Span12Mux_s5_h
    port map (
            O => \N__33789\,
            I => \N__33739\
        );

    \I__7780\ : Sp12to4
    port map (
            O => \N__33786\,
            I => \N__33739\
        );

    \I__7779\ : Sp12to4
    port map (
            O => \N__33781\,
            I => \N__33739\
        );

    \I__7778\ : Span12Mux_v
    port map (
            O => \N__33778\,
            I => \N__33730\
        );

    \I__7777\ : Span12Mux_s6_h
    port map (
            O => \N__33775\,
            I => \N__33730\
        );

    \I__7776\ : Span12Mux_s5_h
    port map (
            O => \N__33772\,
            I => \N__33730\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__33769\,
            I => \N__33730\
        );

    \I__7774\ : Odrv4
    port map (
            O => \N__33766\,
            I => fpga_osc
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__33763\,
            I => fpga_osc
        );

    \I__7772\ : Odrv4
    port map (
            O => \N__33758\,
            I => fpga_osc
        );

    \I__7771\ : Odrv4
    port map (
            O => \N__33751\,
            I => fpga_osc
        );

    \I__7770\ : Odrv4
    port map (
            O => \N__33746\,
            I => fpga_osc
        );

    \I__7769\ : Odrv12
    port map (
            O => \N__33739\,
            I => fpga_osc
        );

    \I__7768\ : Odrv12
    port map (
            O => \N__33730\,
            I => fpga_osc
        );

    \I__7767\ : CEMux
    port map (
            O => \N__33715\,
            I => \N__33712\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__33712\,
            I => \VPP_VDDQ.N_29_0\
        );

    \I__7765\ : SRMux
    port map (
            O => \N__33709\,
            I => \N__33706\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__33706\,
            I => \N__33700\
        );

    \I__7763\ : SRMux
    port map (
            O => \N__33705\,
            I => \N__33697\
        );

    \I__7762\ : SRMux
    port map (
            O => \N__33704\,
            I => \N__33694\
        );

    \I__7761\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33691\
        );

    \I__7760\ : Span4Mux_s1_h
    port map (
            O => \N__33700\,
            I => \N__33688\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__33697\,
            I => \N__33683\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33683\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__33691\,
            I => \N__33680\
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__33688\,
            I => \G_43\
        );

    \I__7755\ : Odrv4
    port map (
            O => \N__33683\,
            I => \G_43\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__33680\,
            I => \G_43\
        );

    \I__7753\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33669\
        );

    \I__7752\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33666\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__33669\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__33666\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__7749\ : InMux
    port map (
            O => \N__33661\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__7748\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33654\
        );

    \I__7747\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33651\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__33654\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__33651\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__7744\ : InMux
    port map (
            O => \N__33646\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__7743\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33639\
        );

    \I__7742\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33636\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__33639\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__33636\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__7739\ : InMux
    port map (
            O => \N__33631\,
            I => \bfn_12_15_0_\
        );

    \I__7738\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33624\
        );

    \I__7737\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33621\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__33624\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__33621\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__7734\ : InMux
    port map (
            O => \N__33616\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__7733\ : CascadeMux
    port map (
            O => \N__33613\,
            I => \N__33609\
        );

    \I__7732\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33606\
        );

    \I__7731\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33603\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__33606\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__33603\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__7728\ : InMux
    port map (
            O => \N__33598\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__7727\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33591\
        );

    \I__7726\ : InMux
    port map (
            O => \N__33594\,
            I => \N__33588\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__33591\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__33588\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__7723\ : InMux
    port map (
            O => \N__33583\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33580\,
            I => \N__33576\
        );

    \I__7721\ : InMux
    port map (
            O => \N__33579\,
            I => \N__33573\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__33576\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__33573\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33568\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__33565\,
            I => \N__33561\
        );

    \I__7716\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33558\
        );

    \I__7715\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33555\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__33558\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__33555\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33550\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__7711\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33544\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33540\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__33543\,
            I => \N__33536\
        );

    \I__7708\ : Span4Mux_s1_h
    port map (
            O => \N__33540\,
            I => \N__33533\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33539\,
            I => \N__33530\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33527\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__33533\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33530\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33527\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33517\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__33517\,
            I => \POWERLED.count_clk_RNIZ0Z_12\
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__33514\,
            I => \POWERLED.count_clkZ0Z_2_cascade_\
        );

    \I__7699\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__33508\,
            I => \N__33504\
        );

    \I__7697\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33501\
        );

    \I__7696\ : Odrv4
    port map (
            O => \N__33504\,
            I => \POWERLED.count_clk_RNIZ0Z_15\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__33501\,
            I => \POWERLED.count_clk_RNIZ0Z_15\
        );

    \I__7694\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__33493\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1\
        );

    \I__7692\ : CascadeMux
    port map (
            O => \N__33490\,
            I => \N__33480\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__33489\,
            I => \N__33477\
        );

    \I__7690\ : CascadeMux
    port map (
            O => \N__33488\,
            I => \N__33472\
        );

    \I__7689\ : InMux
    port map (
            O => \N__33487\,
            I => \N__33466\
        );

    \I__7688\ : InMux
    port map (
            O => \N__33486\,
            I => \N__33461\
        );

    \I__7687\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33461\
        );

    \I__7686\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33444\
        );

    \I__7685\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33444\
        );

    \I__7684\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33444\
        );

    \I__7683\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33444\
        );

    \I__7682\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33437\
        );

    \I__7681\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33437\
        );

    \I__7680\ : InMux
    port map (
            O => \N__33472\,
            I => \N__33437\
        );

    \I__7679\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33434\
        );

    \I__7678\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33429\
        );

    \I__7677\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33429\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33424\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__33461\,
            I => \N__33424\
        );

    \I__7674\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33419\
        );

    \I__7673\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33419\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__33458\,
            I => \N__33413\
        );

    \I__7671\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33408\
        );

    \I__7670\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33403\
        );

    \I__7669\ : InMux
    port map (
            O => \N__33455\,
            I => \N__33403\
        );

    \I__7668\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33400\
        );

    \I__7667\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33397\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__33444\,
            I => \N__33392\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__33437\,
            I => \N__33392\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__33434\,
            I => \N__33383\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33383\
        );

    \I__7662\ : Span4Mux_v
    port map (
            O => \N__33424\,
            I => \N__33383\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33419\,
            I => \N__33383\
        );

    \I__7660\ : InMux
    port map (
            O => \N__33418\,
            I => \N__33370\
        );

    \I__7659\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33370\
        );

    \I__7658\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33370\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33370\
        );

    \I__7656\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33370\
        );

    \I__7655\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33370\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__33408\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__33403\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__33400\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__33397\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7650\ : Odrv12
    port map (
            O => \N__33392\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7649\ : Odrv4
    port map (
            O => \N__33383\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__33370\,
            I => \POWERLED.func_state_RNIH9594_0_1\
        );

    \I__7647\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33349\
        );

    \I__7646\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33349\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__33349\,
            I => \N__33346\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__33346\,
            I => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\
        );

    \I__7643\ : CascadeMux
    port map (
            O => \N__33343\,
            I => \N__33340\
        );

    \I__7642\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33337\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__33337\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__7640\ : CEMux
    port map (
            O => \N__33334\,
            I => \N__33328\
        );

    \I__7639\ : CEMux
    port map (
            O => \N__33333\,
            I => \N__33325\
        );

    \I__7638\ : CEMux
    port map (
            O => \N__33332\,
            I => \N__33321\
        );

    \I__7637\ : CEMux
    port map (
            O => \N__33331\,
            I => \N__33313\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__33328\,
            I => \N__33310\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__33325\,
            I => \N__33307\
        );

    \I__7634\ : CEMux
    port map (
            O => \N__33324\,
            I => \N__33304\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33321\,
            I => \N__33301\
        );

    \I__7632\ : CascadeMux
    port map (
            O => \N__33320\,
            I => \N__33298\
        );

    \I__7631\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33293\
        );

    \I__7630\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33293\
        );

    \I__7629\ : CEMux
    port map (
            O => \N__33317\,
            I => \N__33282\
        );

    \I__7628\ : CEMux
    port map (
            O => \N__33316\,
            I => \N__33279\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33276\
        );

    \I__7626\ : Span4Mux_v
    port map (
            O => \N__33310\,
            I => \N__33271\
        );

    \I__7625\ : Span4Mux_s0_h
    port map (
            O => \N__33307\,
            I => \N__33271\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__33304\,
            I => \N__33268\
        );

    \I__7623\ : Span4Mux_v
    port map (
            O => \N__33301\,
            I => \N__33264\
        );

    \I__7622\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33261\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__33293\,
            I => \N__33258\
        );

    \I__7620\ : CascadeMux
    port map (
            O => \N__33292\,
            I => \N__33254\
        );

    \I__7619\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33247\
        );

    \I__7618\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33247\
        );

    \I__7617\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33247\
        );

    \I__7616\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33238\
        );

    \I__7615\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33238\
        );

    \I__7614\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33238\
        );

    \I__7613\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33238\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33232\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__33279\,
            I => \N__33229\
        );

    \I__7610\ : Span4Mux_v
    port map (
            O => \N__33276\,
            I => \N__33224\
        );

    \I__7609\ : Span4Mux_h
    port map (
            O => \N__33271\,
            I => \N__33224\
        );

    \I__7608\ : Sp12to4
    port map (
            O => \N__33268\,
            I => \N__33221\
        );

    \I__7607\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33218\
        );

    \I__7606\ : Span4Mux_h
    port map (
            O => \N__33264\,
            I => \N__33211\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__33261\,
            I => \N__33211\
        );

    \I__7604\ : Span4Mux_v
    port map (
            O => \N__33258\,
            I => \N__33211\
        );

    \I__7603\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33206\
        );

    \I__7602\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33206\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__33247\,
            I => \N__33201\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33201\
        );

    \I__7599\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33194\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33194\
        );

    \I__7597\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33194\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__33232\,
            I => \POWERLED.count_clk_en\
        );

    \I__7595\ : Odrv12
    port map (
            O => \N__33229\,
            I => \POWERLED.count_clk_en\
        );

    \I__7594\ : Odrv4
    port map (
            O => \N__33224\,
            I => \POWERLED.count_clk_en\
        );

    \I__7593\ : Odrv12
    port map (
            O => \N__33221\,
            I => \POWERLED.count_clk_en\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__33218\,
            I => \POWERLED.count_clk_en\
        );

    \I__7591\ : Odrv4
    port map (
            O => \N__33211\,
            I => \POWERLED.count_clk_en\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__33206\,
            I => \POWERLED.count_clk_en\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__33201\,
            I => \POWERLED.count_clk_en\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__33194\,
            I => \POWERLED.count_clk_en\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__33175\,
            I => \N__33171\
        );

    \I__7586\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33168\
        );

    \I__7585\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33165\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__33168\,
            I => \VPP_VDDQ.N_66_i\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__33165\,
            I => \VPP_VDDQ.N_66_i\
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__33160\,
            I => \N__33156\
        );

    \I__7581\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33153\
        );

    \I__7580\ : InMux
    port map (
            O => \N__33156\,
            I => \N__33150\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__33153\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__33150\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__7577\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33141\
        );

    \I__7576\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33138\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__33141\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__33138\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__7573\ : InMux
    port map (
            O => \N__33133\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__7572\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33126\
        );

    \I__7571\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33123\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__33126\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__33123\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__7568\ : InMux
    port map (
            O => \N__33118\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__33115\,
            I => \N__33111\
        );

    \I__7566\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33108\
        );

    \I__7565\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33105\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__33108\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__33105\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__7562\ : InMux
    port map (
            O => \N__33100\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__7561\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33093\
        );

    \I__7560\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33090\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__33093\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__33090\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__7557\ : InMux
    port map (
            O => \N__33085\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__7556\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33078\
        );

    \I__7555\ : InMux
    port map (
            O => \N__33081\,
            I => \N__33075\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__33078\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__33075\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__7552\ : InMux
    port map (
            O => \N__33070\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__7551\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33061\
        );

    \I__7550\ : InMux
    port map (
            O => \N__33066\,
            I => \N__33061\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__33061\,
            I => \N__33057\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__33060\,
            I => \N__33054\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__33057\,
            I => \N__33051\
        );

    \I__7546\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33048\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__33051\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__33048\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__7543\ : CascadeMux
    port map (
            O => \N__33043\,
            I => \N__33040\
        );

    \I__7542\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33036\
        );

    \I__7541\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33033\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__33036\,
            I => \N__33030\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__33033\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__7538\ : Odrv4
    port map (
            O => \N__33030\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__7537\ : CascadeMux
    port map (
            O => \N__33025\,
            I => \N__33021\
        );

    \I__7536\ : CascadeMux
    port map (
            O => \N__33024\,
            I => \N__33015\
        );

    \I__7535\ : InMux
    port map (
            O => \N__33021\,
            I => \N__33011\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__33020\,
            I => \N__33008\
        );

    \I__7533\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33005\
        );

    \I__7532\ : InMux
    port map (
            O => \N__33018\,
            I => \N__33002\
        );

    \I__7531\ : InMux
    port map (
            O => \N__33015\,
            I => \N__32997\
        );

    \I__7530\ : InMux
    port map (
            O => \N__33014\,
            I => \N__32997\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__33011\,
            I => \N__32994\
        );

    \I__7528\ : InMux
    port map (
            O => \N__33008\,
            I => \N__32991\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__33005\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__33002\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__32997\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__7524\ : Odrv4
    port map (
            O => \N__32994\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__32991\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__32980\,
            I => \POWERLED.un2_count_clk_15_0_9_cascade_\
        );

    \I__7521\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__32974\,
            I => \POWERLED.un2_count_clk_15_0_8\
        );

    \I__7519\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32960\
        );

    \I__7518\ : CascadeMux
    port map (
            O => \N__32970\,
            I => \N__32957\
        );

    \I__7517\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32953\
        );

    \I__7516\ : InMux
    port map (
            O => \N__32968\,
            I => \N__32948\
        );

    \I__7515\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \N__32945\
        );

    \I__7514\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32939\
        );

    \I__7513\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32939\
        );

    \I__7512\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32934\
        );

    \I__7511\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32934\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32931\
        );

    \I__7509\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32928\
        );

    \I__7508\ : InMux
    port map (
            O => \N__32956\,
            I => \N__32925\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__32953\,
            I => \N__32922\
        );

    \I__7506\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32919\
        );

    \I__7505\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32916\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__32948\,
            I => \N__32912\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32909\
        );

    \I__7502\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32906\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__32939\,
            I => \N__32901\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__32934\,
            I => \N__32901\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__32931\,
            I => \N__32898\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__32928\,
            I => \N__32893\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32893\
        );

    \I__7496\ : Span4Mux_v
    port map (
            O => \N__32922\,
            I => \N__32886\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32886\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__32916\,
            I => \N__32886\
        );

    \I__7493\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32883\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__32912\,
            I => \N__32877\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32877\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32874\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__32901\,
            I => \N__32867\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__32898\,
            I => \N__32867\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__32893\,
            I => \N__32867\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__32886\,
            I => \N__32862\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32862\
        );

    \I__7484\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32859\
        );

    \I__7483\ : Span4Mux_h
    port map (
            O => \N__32877\,
            I => \N__32854\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__32874\,
            I => \N__32854\
        );

    \I__7481\ : Span4Mux_h
    port map (
            O => \N__32867\,
            I => \N__32849\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__32862\,
            I => \N__32849\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__32859\,
            I => \POWERLED.un2_count_clk_15_1\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__32854\,
            I => \POWERLED.un2_count_clk_15_1\
        );

    \I__7477\ : Odrv4
    port map (
            O => \N__32849\,
            I => \POWERLED.un2_count_clk_15_1\
        );

    \I__7476\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32837\
        );

    \I__7475\ : InMux
    port map (
            O => \N__32841\,
            I => \N__32832\
        );

    \I__7474\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32832\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32829\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__32832\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__7471\ : Odrv4
    port map (
            O => \N__32829\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__7470\ : CascadeMux
    port map (
            O => \N__32824\,
            I => \N__32818\
        );

    \I__7469\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32813\
        );

    \I__7468\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32813\
        );

    \I__7467\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32810\
        );

    \I__7466\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32807\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__32813\,
            I => \N__32804\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__32810\,
            I => \N__32801\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32798\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__32804\,
            I => \N__32795\
        );

    \I__7461\ : Span4Mux_s2_h
    port map (
            O => \N__32801\,
            I => \N__32792\
        );

    \I__7460\ : Span4Mux_s2_h
    port map (
            O => \N__32798\,
            I => \N__32789\
        );

    \I__7459\ : Odrv4
    port map (
            O => \N__32795\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__32792\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__32789\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__7456\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32779\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__32779\,
            I => \POWERLED.un2_count_clk_15_0_10\
        );

    \I__7454\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32773\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__32773\,
            I => \N__32770\
        );

    \I__7452\ : Odrv12
    port map (
            O => \N__32770\,
            I => \POWERLED.count_clk_0_12\
        );

    \I__7451\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32763\
        );

    \I__7450\ : InMux
    port map (
            O => \N__32766\,
            I => \N__32760\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__32763\,
            I => \N__32757\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__32760\,
            I => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__32757\,
            I => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__32752\,
            I => \N__32749\
        );

    \I__7445\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32746\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__32746\,
            I => \N__32743\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__32743\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__32740\,
            I => \POWERLED.count_clkZ0Z_12_cascade_\
        );

    \I__7441\ : CascadeMux
    port map (
            O => \N__32737\,
            I => \N__32732\
        );

    \I__7440\ : InMux
    port map (
            O => \N__32736\,
            I => \N__32729\
        );

    \I__7439\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32723\
        );

    \I__7438\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32723\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32720\
        );

    \I__7436\ : CascadeMux
    port map (
            O => \N__32728\,
            I => \N__32717\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__32723\,
            I => \N__32714\
        );

    \I__7434\ : Span4Mux_s3_h
    port map (
            O => \N__32720\,
            I => \N__32711\
        );

    \I__7433\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32708\
        );

    \I__7432\ : Span4Mux_s2_h
    port map (
            O => \N__32714\,
            I => \N__32705\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__32711\,
            I => \N__32700\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32700\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__32705\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__32700\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__7427\ : CascadeMux
    port map (
            O => \N__32695\,
            I => \POWERLED.count_clk_RNIZ0Z_12_cascade_\
        );

    \I__7426\ : CascadeMux
    port map (
            O => \N__32692\,
            I => \N__32689\
        );

    \I__7425\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32686\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__32686\,
            I => \POWERLED.un2_count_clk_15_0_7\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__32683\,
            I => \N__32680\
        );

    \I__7422\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32675\
        );

    \I__7421\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32672\
        );

    \I__7420\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32669\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__32675\,
            I => \N__32666\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__32672\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__32669\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__7416\ : Odrv4
    port map (
            O => \N__32666\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__7415\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32653\
        );

    \I__7414\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32653\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32650\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__32650\,
            I => \N__32647\
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__32647\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__7410\ : CascadeMux
    port map (
            O => \N__32644\,
            I => \N__32641\
        );

    \I__7409\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32638\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__32638\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__7407\ : CascadeMux
    port map (
            O => \N__32635\,
            I => \N__32632\
        );

    \I__7406\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32628\
        );

    \I__7405\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32625\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__32628\,
            I => \N__32622\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__32625\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__7402\ : Odrv12
    port map (
            O => \N__32622\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__32617\,
            I => \POWERLED.count_clkZ0Z_15_cascade_\
        );

    \I__7400\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32607\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32602\
        );

    \I__7398\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32602\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32599\
        );

    \I__7396\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32596\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32607\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__32602\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__32599\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__32596\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__7391\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32584\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__32584\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__7389\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32575\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32575\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__32575\,
            I => \N__32572\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__32572\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__7385\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32566\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__32566\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__7383\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32560\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__32560\,
            I => \POWERLED.count_clk_0_10\
        );

    \I__7381\ : InMux
    port map (
            O => \N__32557\,
            I => \N__32551\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32556\,
            I => \N__32551\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__32551\,
            I => \N__32548\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__32548\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__7377\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32541\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__32544\,
            I => \N__32537\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__32541\,
            I => \N__32534\
        );

    \I__7374\ : InMux
    port map (
            O => \N__32540\,
            I => \N__32531\
        );

    \I__7373\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32528\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__32534\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__32531\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32528\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__32521\,
            I => \POWERLED.count_clkZ0Z_10_cascade_\
        );

    \I__7368\ : InMux
    port map (
            O => \N__32518\,
            I => \N__32515\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32511\
        );

    \I__7366\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32508\
        );

    \I__7365\ : Span4Mux_s1_h
    port map (
            O => \N__32511\,
            I => \N__32503\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__32508\,
            I => \N__32503\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__32503\,
            I => \POWERLED.count_clk_RNIZ0Z_13\
        );

    \I__7362\ : CascadeMux
    port map (
            O => \N__32500\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_cascade_\
        );

    \I__7361\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32485\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32485\
        );

    \I__7359\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32485\
        );

    \I__7358\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32485\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__32485\,
            I => \N__32481\
        );

    \I__7356\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32478\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__32481\,
            I => \POWERLED.N_352\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__32478\,
            I => \POWERLED.N_352\
        );

    \I__7353\ : InMux
    port map (
            O => \N__32473\,
            I => \POWERLED.un1_count_clk_2_cry_11\
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__32470\,
            I => \N__32466\
        );

    \I__7351\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32463\
        );

    \I__7350\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32460\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__32463\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__32460\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__7347\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32449\
        );

    \I__7346\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32449\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__32449\,
            I => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\
        );

    \I__7344\ : InMux
    port map (
            O => \N__32446\,
            I => \POWERLED.un1_count_clk_2_cry_12\
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__32443\,
            I => \N__32440\
        );

    \I__7342\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32437\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32437\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__7340\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32428\
        );

    \I__7339\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32428\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__32428\,
            I => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\
        );

    \I__7337\ : InMux
    port map (
            O => \N__32425\,
            I => \POWERLED.un1_count_clk_2_cry_13\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32422\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__32419\,
            I => \N__32415\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__32418\,
            I => \N__32410\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32407\
        );

    \I__7332\ : InMux
    port map (
            O => \N__32414\,
            I => \N__32402\
        );

    \I__7331\ : InMux
    port map (
            O => \N__32413\,
            I => \N__32402\
        );

    \I__7330\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32399\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32396\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__32402\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__32399\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__32396\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__7325\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32383\
        );

    \I__7324\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32383\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__32383\,
            I => \N__32380\
        );

    \I__7322\ : Odrv4
    port map (
            O => \N__32380\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__7321\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32374\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__32374\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__7319\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32368\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__32368\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__7317\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32359\
        );

    \I__7316\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32359\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__32359\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__7314\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32353\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__32353\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__7312\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32346\
        );

    \I__7311\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32343\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__32346\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__32343\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__7308\ : InMux
    port map (
            O => \N__32338\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__7307\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32331\
        );

    \I__7306\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32328\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__32331\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__32328\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__7303\ : InMux
    port map (
            O => \N__32323\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__7302\ : InMux
    port map (
            O => \N__32320\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__7301\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32311\
        );

    \I__7300\ : InMux
    port map (
            O => \N__32316\,
            I => \N__32311\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__32311\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32308\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__7297\ : CascadeMux
    port map (
            O => \N__32305\,
            I => \N__32301\
        );

    \I__7296\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32296\
        );

    \I__7295\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32296\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32293\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__32293\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__7292\ : InMux
    port map (
            O => \N__32290\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__7291\ : InMux
    port map (
            O => \N__32287\,
            I => \POWERLED.un1_count_clk_2_cry_7\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__32284\,
            I => \N__32280\
        );

    \I__7289\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32275\
        );

    \I__7288\ : InMux
    port map (
            O => \N__32280\,
            I => \N__32275\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__32275\,
            I => \N__32272\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__32272\,
            I => \N__32269\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__32269\,
            I => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\
        );

    \I__7284\ : InMux
    port map (
            O => \N__32266\,
            I => \bfn_12_10_0_\
        );

    \I__7283\ : InMux
    port map (
            O => \N__32263\,
            I => \POWERLED.un1_count_clk_2_cry_9\
        );

    \I__7282\ : InMux
    port map (
            O => \N__32260\,
            I => \POWERLED.un1_count_clk_2_cry_10\
        );

    \I__7281\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32251\
        );

    \I__7280\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32251\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__32251\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__7278\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32245\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__32245\,
            I => \N__32242\
        );

    \I__7276\ : Odrv4
    port map (
            O => \N__32242\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__7275\ : CascadeMux
    port map (
            O => \N__32239\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1_cascade_\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__32236\,
            I => \N__32232\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__32235\,
            I => \N__32229\
        );

    \I__7272\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32224\
        );

    \I__7271\ : InMux
    port map (
            O => \N__32229\,
            I => \N__32221\
        );

    \I__7270\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32216\
        );

    \I__7269\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32216\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32213\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__32221\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__32216\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7265\ : Odrv12
    port map (
            O => \N__32213\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__32206\,
            I => \N__32203\
        );

    \I__7263\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32200\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__32200\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__32197\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__32194\,
            I => \N__32191\
        );

    \I__7259\ : InMux
    port map (
            O => \N__32191\,
            I => \N__32185\
        );

    \I__7258\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32185\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__32185\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__32182\,
            I => \N__32178\
        );

    \I__7255\ : CascadeMux
    port map (
            O => \N__32181\,
            I => \N__32174\
        );

    \I__7254\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32155\
        );

    \I__7253\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32155\
        );

    \I__7252\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32155\
        );

    \I__7251\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32155\
        );

    \I__7250\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32143\
        );

    \I__7249\ : InMux
    port map (
            O => \N__32171\,
            I => \N__32130\
        );

    \I__7248\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32130\
        );

    \I__7247\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32130\
        );

    \I__7246\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32130\
        );

    \I__7245\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32130\
        );

    \I__7244\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32130\
        );

    \I__7243\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32127\
        );

    \I__7242\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32124\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__32155\,
            I => \N__32121\
        );

    \I__7240\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32112\
        );

    \I__7239\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32112\
        );

    \I__7238\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32112\
        );

    \I__7237\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32112\
        );

    \I__7236\ : CascadeMux
    port map (
            O => \N__32150\,
            I => \N__32108\
        );

    \I__7235\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32098\
        );

    \I__7234\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32098\
        );

    \I__7233\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32098\
        );

    \I__7232\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32098\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32095\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32092\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__32127\,
            I => \N__32074\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__32124\,
            I => \N__32074\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__32121\,
            I => \N__32074\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__32112\,
            I => \N__32074\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__32111\,
            I => \N__32070\
        );

    \I__7224\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32065\
        );

    \I__7223\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32062\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__32098\,
            I => \N__32059\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__32095\,
            I => \N__32056\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__32092\,
            I => \N__32053\
        );

    \I__7219\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32044\
        );

    \I__7218\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32044\
        );

    \I__7217\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32044\
        );

    \I__7216\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32044\
        );

    \I__7215\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32033\
        );

    \I__7214\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32033\
        );

    \I__7213\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32033\
        );

    \I__7212\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32033\
        );

    \I__7211\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32033\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__32074\,
            I => \N__32030\
        );

    \I__7209\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32021\
        );

    \I__7208\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32021\
        );

    \I__7207\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32021\
        );

    \I__7206\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32021\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__32065\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__32062\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__32059\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__32056\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7201\ : Odrv4
    port map (
            O => \N__32053\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__32044\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__32033\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7198\ : Odrv4
    port map (
            O => \N__32030\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__32021\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__32002\,
            I => \N__31998\
        );

    \I__7195\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31993\
        );

    \I__7194\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31993\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31993\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__7192\ : CascadeMux
    port map (
            O => \N__31990\,
            I => \N__31985\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__31989\,
            I => \N__31976\
        );

    \I__7190\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31968\
        );

    \I__7189\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31957\
        );

    \I__7188\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31957\
        );

    \I__7187\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31957\
        );

    \I__7186\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31957\
        );

    \I__7185\ : InMux
    port map (
            O => \N__31981\,
            I => \N__31957\
        );

    \I__7184\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31954\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__31979\,
            I => \N__31944\
        );

    \I__7182\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31936\
        );

    \I__7181\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31936\
        );

    \I__7180\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31931\
        );

    \I__7179\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31931\
        );

    \I__7178\ : CascadeMux
    port map (
            O => \N__31972\,
            I => \N__31928\
        );

    \I__7177\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31922\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__31968\,
            I => \N__31915\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31915\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31915\
        );

    \I__7173\ : CascadeMux
    port map (
            O => \N__31953\,
            I => \N__31903\
        );

    \I__7172\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31898\
        );

    \I__7171\ : InMux
    port map (
            O => \N__31951\,
            I => \N__31889\
        );

    \I__7170\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31889\
        );

    \I__7169\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31889\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31889\
        );

    \I__7167\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31884\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31884\
        );

    \I__7165\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31881\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31876\
        );

    \I__7163\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31876\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31871\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31871\
        );

    \I__7160\ : InMux
    port map (
            O => \N__31928\,
            I => \N__31866\
        );

    \I__7159\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31866\
        );

    \I__7158\ : InMux
    port map (
            O => \N__31926\,
            I => \N__31861\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31861\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__31922\,
            I => \N__31856\
        );

    \I__7155\ : Span4Mux_v
    port map (
            O => \N__31915\,
            I => \N__31856\
        );

    \I__7154\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31845\
        );

    \I__7153\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31845\
        );

    \I__7152\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31845\
        );

    \I__7151\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31845\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31845\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31836\
        );

    \I__7148\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31836\
        );

    \I__7147\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31836\
        );

    \I__7146\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31836\
        );

    \I__7145\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31829\
        );

    \I__7144\ : InMux
    port map (
            O => \N__31902\,
            I => \N__31829\
        );

    \I__7143\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31829\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31824\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__31889\,
            I => \N__31824\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__31884\,
            I => \N__31815\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__31881\,
            I => \N__31815\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__31876\,
            I => \N__31815\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__31871\,
            I => \N__31815\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__31866\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__31861\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__31856\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__31845\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__31836\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__31829\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7130\ : Odrv12
    port map (
            O => \N__31824\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__31815\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7128\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31787\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__31797\,
            I => \N__31771\
        );

    \I__7126\ : CascadeMux
    port map (
            O => \N__31796\,
            I => \N__31767\
        );

    \I__7125\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31749\
        );

    \I__7124\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31749\
        );

    \I__7123\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31749\
        );

    \I__7122\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31749\
        );

    \I__7121\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31749\
        );

    \I__7120\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31749\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__31787\,
            I => \N__31739\
        );

    \I__7118\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31730\
        );

    \I__7117\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31730\
        );

    \I__7116\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31730\
        );

    \I__7115\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31730\
        );

    \I__7114\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31721\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31721\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31721\
        );

    \I__7111\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31721\
        );

    \I__7110\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31710\
        );

    \I__7109\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31710\
        );

    \I__7108\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31710\
        );

    \I__7107\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31710\
        );

    \I__7106\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31710\
        );

    \I__7105\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31707\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31702\
        );

    \I__7103\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31702\
        );

    \I__7102\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31699\
        );

    \I__7101\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31690\
        );

    \I__7100\ : InMux
    port map (
            O => \N__31764\,
            I => \N__31690\
        );

    \I__7099\ : InMux
    port map (
            O => \N__31763\,
            I => \N__31690\
        );

    \I__7098\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31690\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__31749\,
            I => \N__31687\
        );

    \I__7096\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31680\
        );

    \I__7095\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31680\
        );

    \I__7094\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31680\
        );

    \I__7093\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31671\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31671\
        );

    \I__7091\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31671\
        );

    \I__7090\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31671\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__31739\,
            I => \N__31664\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__31730\,
            I => \N__31664\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__31721\,
            I => \N__31664\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__31710\,
            I => \N__31661\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31707\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__31702\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__31699\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__31690\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7081\ : Odrv4
    port map (
            O => \N__31687\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__31680\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__31671\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__31664\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__31661\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7076\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31639\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__31639\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__31636\,
            I => \VPP_VDDQ.count_2_1_11_cascade_\
        );

    \I__7073\ : CEMux
    port map (
            O => \N__31633\,
            I => \N__31628\
        );

    \I__7072\ : CEMux
    port map (
            O => \N__31632\,
            I => \N__31623\
        );

    \I__7071\ : CEMux
    port map (
            O => \N__31631\,
            I => \N__31615\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__31628\,
            I => \N__31612\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31607\
        );

    \I__7068\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31607\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__31623\,
            I => \N__31601\
        );

    \I__7066\ : CEMux
    port map (
            O => \N__31622\,
            I => \N__31598\
        );

    \I__7065\ : CEMux
    port map (
            O => \N__31621\,
            I => \N__31595\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31620\,
            I => \N__31591\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31584\
        );

    \I__7062\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31584\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31577\
        );

    \I__7060\ : Span4Mux_v
    port map (
            O => \N__31612\,
            I => \N__31577\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31577\
        );

    \I__7058\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31570\
        );

    \I__7057\ : InMux
    port map (
            O => \N__31605\,
            I => \N__31570\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31570\
        );

    \I__7055\ : Span4Mux_h
    port map (
            O => \N__31601\,
            I => \N__31559\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__31598\,
            I => \N__31559\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31559\
        );

    \I__7052\ : CEMux
    port map (
            O => \N__31594\,
            I => \N__31556\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__31591\,
            I => \N__31553\
        );

    \I__7050\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31542\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31542\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__31584\,
            I => \N__31535\
        );

    \I__7047\ : Span4Mux_h
    port map (
            O => \N__31577\,
            I => \N__31535\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__31570\,
            I => \N__31535\
        );

    \I__7045\ : CEMux
    port map (
            O => \N__31569\,
            I => \N__31526\
        );

    \I__7044\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31526\
        );

    \I__7043\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31526\
        );

    \I__7042\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31526\
        );

    \I__7041\ : Span4Mux_v
    port map (
            O => \N__31559\,
            I => \N__31523\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31520\
        );

    \I__7039\ : Span4Mux_v
    port map (
            O => \N__31553\,
            I => \N__31517\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31510\
        );

    \I__7037\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31510\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31510\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31507\
        );

    \I__7034\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31502\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31502\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31495\
        );

    \I__7031\ : Sp12to4
    port map (
            O => \N__31535\,
            I => \N__31495\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__31526\,
            I => \N__31495\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__31523\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__31520\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7027\ : Odrv4
    port map (
            O => \N__31517\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__31510\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__31507\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__31502\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7023\ : Odrv12
    port map (
            O => \N__31495\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7022\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31476\
        );

    \I__7021\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31473\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__31476\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__31473\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__7018\ : InMux
    port map (
            O => \N__31468\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__7017\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31462\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__31462\,
            I => \VPP_VDDQ.count_2_1_12\
        );

    \I__7015\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31456\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__31456\,
            I => \VPP_VDDQ.count_2_1_13\
        );

    \I__7013\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31450\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__31450\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__7011\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31443\
        );

    \I__7010\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31440\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__31443\,
            I => \N__31437\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__31440\,
            I => \N__31434\
        );

    \I__7007\ : Odrv4
    port map (
            O => \N__31437\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__31434\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__7005\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31425\
        );

    \I__7004\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__31425\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__31422\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \VPP_VDDQ.count_2Z0Z_13_cascade_\
        );

    \I__7000\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31411\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__31411\,
            I => \N__31407\
        );

    \I__6998\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31404\
        );

    \I__6997\ : Sp12to4
    port map (
            O => \N__31407\,
            I => \N__31401\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31398\
        );

    \I__6995\ : Odrv12
    port map (
            O => \N__31401\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__31398\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__6993\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31390\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__31390\,
            I => \VPP_VDDQ.un9_clk_100khz_10\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__31387\,
            I => \N__31383\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__31386\,
            I => \N__31380\
        );

    \I__6989\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31375\
        );

    \I__6988\ : InMux
    port map (
            O => \N__31380\,
            I => \N__31375\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__31375\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\
        );

    \I__6986\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31369\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__31369\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__31366\,
            I => \N__31362\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__31365\,
            I => \N__31359\
        );

    \I__6982\ : InMux
    port map (
            O => \N__31362\,
            I => \N__31356\
        );

    \I__6981\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31353\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__31356\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__31353\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31345\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__31345\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__6976\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31339\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31335\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31332\
        );

    \I__6973\ : Span4Mux_s1_h
    port map (
            O => \N__31335\,
            I => \N__31329\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__31332\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__6971\ : Odrv4
    port map (
            O => \N__31329\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__6970\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31321\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__31321\,
            I => \N__31318\
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__31318\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__6967\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31312\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__31312\,
            I => \N__31309\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__31309\,
            I => \VPP_VDDQ.un9_clk_100khz_1\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31303\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__31303\,
            I => \VPP_VDDQ.count_2_0_5\
        );

    \I__6962\ : CascadeMux
    port map (
            O => \N__31300\,
            I => \VPP_VDDQ.count_2_1_5_cascade_\
        );

    \I__6961\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31293\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31290\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__31293\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__31290\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__6957\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31282\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__31282\,
            I => \N__31279\
        );

    \I__6955\ : Span4Mux_v
    port map (
            O => \N__31279\,
            I => \N__31276\
        );

    \I__6954\ : Span4Mux_h
    port map (
            O => \N__31276\,
            I => \N__31273\
        );

    \I__6953\ : Span4Mux_h
    port map (
            O => \N__31273\,
            I => \N__31270\
        );

    \I__6952\ : Odrv4
    port map (
            O => \N__31270\,
            I => vr_ready_vccin
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__6950\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31258\
        );

    \I__6949\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31258\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__31255\,
            I => \N__31250\
        );

    \I__6946\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31245\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31245\
        );

    \I__6944\ : Span4Mux_h
    port map (
            O => \N__31250\,
            I => \N__31240\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__31245\,
            I => \N__31240\
        );

    \I__6942\ : Odrv4
    port map (
            O => \N__31240\,
            I => \PCH_PWRGD.N_174\
        );

    \I__6941\ : IoInMux
    port map (
            O => \N__31237\,
            I => \N__31233\
        );

    \I__6940\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31230\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__31233\,
            I => \N__31227\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31224\
        );

    \I__6937\ : Span4Mux_s0_h
    port map (
            O => \N__31227\,
            I => \N__31221\
        );

    \I__6936\ : Span12Mux_s3_h
    port map (
            O => \N__31224\,
            I => \N__31218\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__31221\,
            I => \N__31215\
        );

    \I__6934\ : Odrv12
    port map (
            O => \N__31218\,
            I => dsw_pwrok
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__31215\,
            I => dsw_pwrok
        );

    \I__6932\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31207\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__31207\,
            I => \N__31204\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__31204\,
            I => \N__31201\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__31201\,
            I => vccst_cpu_ok
        );

    \I__6928\ : CascadeMux
    port map (
            O => \N__31198\,
            I => \N__31195\
        );

    \I__6927\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31192\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__31192\,
            I => v5s_ok
        );

    \I__6925\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31186\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__31186\,
            I => \N__31183\
        );

    \I__6923\ : Span12Mux_v
    port map (
            O => \N__31183\,
            I => \N__31180\
        );

    \I__6922\ : Odrv12
    port map (
            O => \N__31180\,
            I => v33s_ok
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__31177\,
            I => \N__31173\
        );

    \I__6920\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31168\
        );

    \I__6919\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31168\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31160\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__31167\,
            I => \N__31155\
        );

    \I__6916\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31150\
        );

    \I__6915\ : CascadeMux
    port map (
            O => \N__31165\,
            I => \N__31142\
        );

    \I__6914\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31134\
        );

    \I__6913\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31134\
        );

    \I__6912\ : Span4Mux_s3_v
    port map (
            O => \N__31160\,
            I => \N__31129\
        );

    \I__6911\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31124\
        );

    \I__6910\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31124\
        );

    \I__6909\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31121\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__31154\,
            I => \N__31117\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__31153\,
            I => \N__31111\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31105\
        );

    \I__6905\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31102\
        );

    \I__6904\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31099\
        );

    \I__6903\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31090\
        );

    \I__6902\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31090\
        );

    \I__6901\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31090\
        );

    \I__6900\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31090\
        );

    \I__6899\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31085\
        );

    \I__6898\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31085\
        );

    \I__6897\ : InMux
    port map (
            O => \N__31139\,
            I => \N__31082\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31079\
        );

    \I__6895\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31076\
        );

    \I__6894\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31073\
        );

    \I__6893\ : Span4Mux_h
    port map (
            O => \N__31129\,
            I => \N__31068\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__31124\,
            I => \N__31068\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__31121\,
            I => \N__31065\
        );

    \I__6890\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31060\
        );

    \I__6889\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31060\
        );

    \I__6888\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31055\
        );

    \I__6887\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31055\
        );

    \I__6886\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31050\
        );

    \I__6885\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31050\
        );

    \I__6884\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31045\
        );

    \I__6883\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31045\
        );

    \I__6882\ : CascadeMux
    port map (
            O => \N__31108\,
            I => \N__31042\
        );

    \I__6881\ : Span4Mux_v
    port map (
            O => \N__31105\,
            I => \N__31039\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__31102\,
            I => \N__31032\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__31099\,
            I => \N__31032\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31032\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31029\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31019\
        );

    \I__6875\ : Span4Mux_h
    port map (
            O => \N__31079\,
            I => \N__31019\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__31076\,
            I => \N__31019\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31016\
        );

    \I__6872\ : Span4Mux_h
    port map (
            O => \N__31068\,
            I => \N__31013\
        );

    \I__6871\ : Span4Mux_h
    port map (
            O => \N__31065\,
            I => \N__31006\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__31006\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__31055\,
            I => \N__31006\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__31050\,
            I => \N__31001\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__31045\,
            I => \N__31001\
        );

    \I__6866\ : InMux
    port map (
            O => \N__31042\,
            I => \N__30998\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__31039\,
            I => \N__30991\
        );

    \I__6864\ : Span4Mux_v
    port map (
            O => \N__31032\,
            I => \N__30991\
        );

    \I__6863\ : Span4Mux_s3_h
    port map (
            O => \N__31029\,
            I => \N__30991\
        );

    \I__6862\ : InMux
    port map (
            O => \N__31028\,
            I => \N__30984\
        );

    \I__6861\ : InMux
    port map (
            O => \N__31027\,
            I => \N__30984\
        );

    \I__6860\ : InMux
    port map (
            O => \N__31026\,
            I => \N__30984\
        );

    \I__6859\ : Span4Mux_v
    port map (
            O => \N__31019\,
            I => \N__30981\
        );

    \I__6858\ : Span4Mux_v
    port map (
            O => \N__31016\,
            I => \N__30972\
        );

    \I__6857\ : Span4Mux_v
    port map (
            O => \N__31013\,
            I => \N__30972\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__31006\,
            I => \N__30972\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__31001\,
            I => \N__30972\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__30998\,
            I => slp_s3n_signal
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__30991\,
            I => slp_s3n_signal
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__30984\,
            I => slp_s3n_signal
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__30981\,
            I => slp_s3n_signal
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__30972\,
            I => slp_s3n_signal
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__30961\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\
        );

    \I__6848\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30955\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__30955\,
            I => \N__30952\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__30952\,
            I => \N__30947\
        );

    \I__6845\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30942\
        );

    \I__6844\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30942\
        );

    \I__6843\ : Span4Mux_s0_h
    port map (
            O => \N__30947\,
            I => \N__30935\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30932\
        );

    \I__6841\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30923\
        );

    \I__6840\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30923\
        );

    \I__6839\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30923\
        );

    \I__6838\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30923\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__30935\,
            I => rsmrst_pwrgd_signal
        );

    \I__6836\ : Odrv12
    port map (
            O => \N__30932\,
            I => rsmrst_pwrgd_signal
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__30923\,
            I => rsmrst_pwrgd_signal
        );

    \I__6834\ : IoInMux
    port map (
            O => \N__30916\,
            I => \N__30913\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30910\
        );

    \I__6832\ : IoSpan4Mux
    port map (
            O => \N__30910\,
            I => \N__30907\
        );

    \I__6831\ : Span4Mux_s3_v
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__30904\,
            I => \N__30901\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__30901\,
            I => vccin_en
        );

    \I__6828\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30895\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__30895\,
            I => \VPP_VDDQ.un1_count_2_1_axb_6\
        );

    \I__6826\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30888\
        );

    \I__6825\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30885\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__30888\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__30885\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__6822\ : InMux
    port map (
            O => \N__30880\,
            I => \N__30874\
        );

    \I__6821\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30874\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__30874\,
            I => \N__30871\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__30871\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__6818\ : InMux
    port map (
            O => \N__30868\,
            I => \N__30865\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__30865\,
            I => \VPP_VDDQ.un9_clk_100khz_9\
        );

    \I__6816\ : CascadeMux
    port map (
            O => \N__30862\,
            I => \VPP_VDDQ.un9_clk_100khz_0_cascade_\
        );

    \I__6815\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__30856\,
            I => \N__30853\
        );

    \I__6813\ : Odrv4
    port map (
            O => \N__30853\,
            I => \VPP_VDDQ.un9_clk_100khz_13\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__30850\,
            I => \N__30847\
        );

    \I__6811\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30843\
        );

    \I__6810\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30840\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__30843\,
            I => \N__30837\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__30840\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\
        );

    \I__6807\ : Odrv12
    port map (
            O => \N__30837\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\
        );

    \I__6806\ : CascadeMux
    port map (
            O => \N__30832\,
            I => \VPP_VDDQ.N_1_i_cascade_\
        );

    \I__6805\ : CascadeMux
    port map (
            O => \N__30829\,
            I => \N__30826\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30820\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30820\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__30820\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__6801\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30814\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__30814\,
            I => \VPP_VDDQ.N_361_0\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__30811\,
            I => \N__30804\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30800\
        );

    \I__6797\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30797\
        );

    \I__6796\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30794\
        );

    \I__6795\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30789\
        );

    \I__6794\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30789\
        );

    \I__6793\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30786\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__30800\,
            I => \N__30775\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__30797\,
            I => \N__30772\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30769\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__30789\,
            I => \N__30766\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__30786\,
            I => \N__30763\
        );

    \I__6787\ : CEMux
    port map (
            O => \N__30785\,
            I => \N__30736\
        );

    \I__6786\ : CEMux
    port map (
            O => \N__30784\,
            I => \N__30736\
        );

    \I__6785\ : CEMux
    port map (
            O => \N__30783\,
            I => \N__30736\
        );

    \I__6784\ : CEMux
    port map (
            O => \N__30782\,
            I => \N__30736\
        );

    \I__6783\ : CEMux
    port map (
            O => \N__30781\,
            I => \N__30736\
        );

    \I__6782\ : CEMux
    port map (
            O => \N__30780\,
            I => \N__30736\
        );

    \I__6781\ : CEMux
    port map (
            O => \N__30779\,
            I => \N__30736\
        );

    \I__6780\ : CEMux
    port map (
            O => \N__30778\,
            I => \N__30736\
        );

    \I__6779\ : Glb2LocalMux
    port map (
            O => \N__30775\,
            I => \N__30736\
        );

    \I__6778\ : Glb2LocalMux
    port map (
            O => \N__30772\,
            I => \N__30736\
        );

    \I__6777\ : Glb2LocalMux
    port map (
            O => \N__30769\,
            I => \N__30736\
        );

    \I__6776\ : Glb2LocalMux
    port map (
            O => \N__30766\,
            I => \N__30736\
        );

    \I__6775\ : Glb2LocalMux
    port map (
            O => \N__30763\,
            I => \N__30736\
        );

    \I__6774\ : GlobalMux
    port map (
            O => \N__30736\,
            I => \N__30733\
        );

    \I__6773\ : gio2CtrlBuf
    port map (
            O => \N__30733\,
            I => \N_570_g\
        );

    \I__6772\ : CascadeMux
    port map (
            O => \N__30730\,
            I => \N__30727\
        );

    \I__6771\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30721\
        );

    \I__6770\ : InMux
    port map (
            O => \N__30726\,
            I => \N__30721\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__30721\,
            I => \VPP_VDDQ.N_2192_i\
        );

    \I__6768\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30713\
        );

    \I__6767\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30708\
        );

    \I__6766\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30708\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__30713\,
            I => \VPP_VDDQ.N_62\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__30708\,
            I => \VPP_VDDQ.N_62\
        );

    \I__6763\ : SRMux
    port map (
            O => \N__30703\,
            I => \N__30700\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__30700\,
            I => \N__30697\
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__30697\,
            I => \VPP_VDDQ.N_62_i\
        );

    \I__6760\ : CascadeMux
    port map (
            O => \N__30694\,
            I => \VPP_VDDQ.count_2_1_14_cascade_\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__30691\,
            I => \VPP_VDDQ.count_2_1_4_cascade_\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__30688\,
            I => \N__30684\
        );

    \I__6757\ : CascadeMux
    port map (
            O => \N__30687\,
            I => \N__30681\
        );

    \I__6756\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30676\
        );

    \I__6755\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30676\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30673\
        );

    \I__6753\ : Span4Mux_s0_h
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__30670\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\
        );

    \I__6751\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30664\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__30664\,
            I => \VPP_VDDQ.count_2_0_4\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__30661\,
            I => \N__30657\
        );

    \I__6748\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30652\
        );

    \I__6747\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30652\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__30652\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\
        );

    \I__6745\ : InMux
    port map (
            O => \N__30649\,
            I => \N__30646\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__30646\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__6743\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30640\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__30640\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__6741\ : IoInMux
    port map (
            O => \N__30637\,
            I => \N__30633\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__30636\,
            I => \N__30627\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30624\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__30632\,
            I => \N__30621\
        );

    \I__6737\ : CascadeMux
    port map (
            O => \N__30631\,
            I => \N__30617\
        );

    \I__6736\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30607\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30607\
        );

    \I__6734\ : Span4Mux_s0_h
    port map (
            O => \N__30624\,
            I => \N__30596\
        );

    \I__6733\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30589\
        );

    \I__6732\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30589\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30617\,
            I => \N__30589\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30580\
        );

    \I__6729\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30580\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30580\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30580\
        );

    \I__6726\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30571\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30607\,
            I => \N__30568\
        );

    \I__6724\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30565\
        );

    \I__6723\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30558\
        );

    \I__6722\ : InMux
    port map (
            O => \N__30604\,
            I => \N__30558\
        );

    \I__6721\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30558\
        );

    \I__6720\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30549\
        );

    \I__6719\ : InMux
    port map (
            O => \N__30601\,
            I => \N__30549\
        );

    \I__6718\ : InMux
    port map (
            O => \N__30600\,
            I => \N__30549\
        );

    \I__6717\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30549\
        );

    \I__6716\ : Span4Mux_v
    port map (
            O => \N__30596\,
            I => \N__30539\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__30589\,
            I => \N__30539\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__30580\,
            I => \N__30539\
        );

    \I__6713\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30532\
        );

    \I__6712\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30532\
        );

    \I__6711\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30532\
        );

    \I__6710\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30526\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30526\
        );

    \I__6708\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30523\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30520\
        );

    \I__6706\ : Span4Mux_s2_h
    port map (
            O => \N__30568\,
            I => \N__30511\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30511\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__30558\,
            I => \N__30511\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30511\
        );

    \I__6702\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30508\
        );

    \I__6701\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30503\
        );

    \I__6700\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30503\
        );

    \I__6699\ : Span4Mux_v
    port map (
            O => \N__30539\,
            I => \N__30498\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30498\
        );

    \I__6697\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30495\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30492\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__30523\,
            I => \N__30485\
        );

    \I__6694\ : Span4Mux_v
    port map (
            O => \N__30520\,
            I => \N__30485\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__30511\,
            I => \N__30482\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__30508\,
            I => \N__30477\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__30503\,
            I => \N__30477\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__30498\,
            I => \N__30474\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30469\
        );

    \I__6688\ : Span4Mux_s3_h
    port map (
            O => \N__30492\,
            I => \N__30469\
        );

    \I__6687\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30466\
        );

    \I__6686\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30462\
        );

    \I__6685\ : Span4Mux_v
    port map (
            O => \N__30485\,
            I => \N__30457\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__30482\,
            I => \N__30457\
        );

    \I__6683\ : Span4Mux_s2_h
    port map (
            O => \N__30477\,
            I => \N__30454\
        );

    \I__6682\ : Span4Mux_h
    port map (
            O => \N__30474\,
            I => \N__30447\
        );

    \I__6681\ : Span4Mux_v
    port map (
            O => \N__30469\,
            I => \N__30447\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30447\
        );

    \I__6679\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30444\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__30462\,
            I => suswarn_n
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__30457\,
            I => suswarn_n
        );

    \I__6676\ : Odrv4
    port map (
            O => \N__30454\,
            I => suswarn_n
        );

    \I__6675\ : Odrv4
    port map (
            O => \N__30447\,
            I => suswarn_n
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__30444\,
            I => suswarn_n
        );

    \I__6673\ : CascadeMux
    port map (
            O => \N__30433\,
            I => \VPP_VDDQ.N_361_0_cascade_\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__30430\,
            I => \VPP_VDDQ.N_62_cascade_\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__30427\,
            I => \VPP_VDDQ.delayed_vddq_ok_en_cascade_\
        );

    \I__6670\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30421\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__30421\,
            I => \N__30418\
        );

    \I__6668\ : Span12Mux_s11_h
    port map (
            O => \N__30418\,
            I => \N__30415\
        );

    \I__6667\ : Odrv12
    port map (
            O => \N__30415\,
            I => \VPP_VDDQ_delayed_vddq_ok\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__30412\,
            I => \N__30407\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__30411\,
            I => \N__30403\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30396\
        );

    \I__6663\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30389\
        );

    \I__6662\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30389\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30389\
        );

    \I__6660\ : InMux
    port map (
            O => \N__30402\,
            I => \N__30380\
        );

    \I__6659\ : InMux
    port map (
            O => \N__30401\,
            I => \N__30380\
        );

    \I__6658\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30380\
        );

    \I__6657\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30380\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__30396\,
            I => \N__30375\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30375\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__30380\,
            I => \N__30372\
        );

    \I__6653\ : Span4Mux_v
    port map (
            O => \N__30375\,
            I => \N__30365\
        );

    \I__6652\ : Span4Mux_v
    port map (
            O => \N__30372\,
            I => \N__30365\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30360\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30370\,
            I => \N__30360\
        );

    \I__6649\ : Span4Mux_v
    port map (
            O => \N__30365\,
            I => \N__30353\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__30360\,
            I => \N__30353\
        );

    \I__6647\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30348\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30348\
        );

    \I__6645\ : Span4Mux_v
    port map (
            O => \N__30353\,
            I => \N__30345\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__30348\,
            I => \N__30342\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__30345\,
            I => vddq_ok
        );

    \I__6642\ : Odrv12
    port map (
            O => \N__30342\,
            I => vddq_ok
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \N__30334\
        );

    \I__6640\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__30331\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__6638\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30322\
        );

    \I__6637\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30322\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__30322\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__6635\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30316\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__30316\,
            I => \VPP_VDDQ.curr_state_7_0\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__30313\,
            I => \VPP_VDDQ.curr_state_7_0_cascade_\
        );

    \I__6632\ : InMux
    port map (
            O => \N__30310\,
            I => \N__30307\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__30307\,
            I => \N__30304\
        );

    \I__6630\ : Span4Mux_s2_v
    port map (
            O => \N__30304\,
            I => \N__30300\
        );

    \I__6629\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30297\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__30300\,
            I => \N_246\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__30297\,
            I => \N_246\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__30292\,
            I => \N_246_cascade_\
        );

    \I__6625\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30285\
        );

    \I__6624\ : InMux
    port map (
            O => \N__30288\,
            I => \N__30282\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__30285\,
            I => \N_381\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__30282\,
            I => \N_381\
        );

    \I__6621\ : InMux
    port map (
            O => \N__30277\,
            I => \N__30266\
        );

    \I__6620\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30266\
        );

    \I__6619\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30266\
        );

    \I__6618\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30261\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30261\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__30266\,
            I => \N__30257\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30254\
        );

    \I__6614\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30251\
        );

    \I__6613\ : Span4Mux_s2_h
    port map (
            O => \N__30257\,
            I => \N__30248\
        );

    \I__6612\ : Span12Mux_s3_h
    port map (
            O => \N__30254\,
            I => \N__30245\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__30251\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__30248\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6609\ : Odrv12
    port map (
            O => \N__30245\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__6608\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30234\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__30237\,
            I => \N__30230\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__30234\,
            I => \N__30225\
        );

    \I__6605\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30222\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30219\
        );

    \I__6603\ : CascadeMux
    port map (
            O => \N__30229\,
            I => \N__30215\
        );

    \I__6602\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30209\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__30225\,
            I => \N__30206\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__30222\,
            I => \N__30201\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__30219\,
            I => \N__30201\
        );

    \I__6598\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30194\
        );

    \I__6597\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30194\
        );

    \I__6596\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30194\
        );

    \I__6595\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30191\
        );

    \I__6594\ : IoInMux
    port map (
            O => \N__30212\,
            I => \N__30185\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__30209\,
            I => \N__30178\
        );

    \I__6592\ : Span4Mux_h
    port map (
            O => \N__30206\,
            I => \N__30178\
        );

    \I__6591\ : Span4Mux_v
    port map (
            O => \N__30201\,
            I => \N__30178\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__30194\,
            I => \N__30175\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__30191\,
            I => \N__30172\
        );

    \I__6588\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30169\
        );

    \I__6587\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30166\
        );

    \I__6586\ : CascadeMux
    port map (
            O => \N__30188\,
            I => \N__30161\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30156\
        );

    \I__6584\ : Span4Mux_v
    port map (
            O => \N__30178\,
            I => \N__30153\
        );

    \I__6583\ : Span4Mux_s2_h
    port map (
            O => \N__30175\,
            I => \N__30150\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__30172\,
            I => \N__30144\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30144\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__30166\,
            I => \N__30141\
        );

    \I__6579\ : InMux
    port map (
            O => \N__30165\,
            I => \N__30136\
        );

    \I__6578\ : InMux
    port map (
            O => \N__30164\,
            I => \N__30136\
        );

    \I__6577\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30129\
        );

    \I__6576\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30129\
        );

    \I__6575\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30129\
        );

    \I__6574\ : Span12Mux_s8_h
    port map (
            O => \N__30156\,
            I => \N__30126\
        );

    \I__6573\ : Span4Mux_s0_h
    port map (
            O => \N__30153\,
            I => \N__30123\
        );

    \I__6572\ : Span4Mux_v
    port map (
            O => \N__30150\,
            I => \N__30120\
        );

    \I__6571\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30117\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__30144\,
            I => \N__30108\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__30141\,
            I => \N__30108\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__30136\,
            I => \N__30108\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__30129\,
            I => \N__30108\
        );

    \I__6566\ : Odrv12
    port map (
            O => \N__30126\,
            I => vccst_en
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__30123\,
            I => vccst_en
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__30120\,
            I => vccst_en
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__30117\,
            I => vccst_en
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__30108\,
            I => vccst_en
        );

    \I__6561\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30089\
        );

    \I__6560\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30089\
        );

    \I__6559\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30084\
        );

    \I__6558\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30084\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__30089\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__30084\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__6555\ : CascadeMux
    port map (
            O => \N__30079\,
            I => \VPP_VDDQ.un6_count_10_cascade_\
        );

    \I__6554\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30073\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__30073\,
            I => \N__30069\
        );

    \I__6552\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30066\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__30069\,
            I => \VPP_VDDQ_un6_count\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__30066\,
            I => \VPP_VDDQ_un6_count\
        );

    \I__6549\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30058\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__30058\,
            I => \VPP_VDDQ.un6_count_8\
        );

    \I__6547\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30052\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__30052\,
            I => \N__30045\
        );

    \I__6545\ : InMux
    port map (
            O => \N__30051\,
            I => \N__30042\
        );

    \I__6544\ : InMux
    port map (
            O => \N__30050\,
            I => \N__30039\
        );

    \I__6543\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30032\
        );

    \I__6542\ : InMux
    port map (
            O => \N__30048\,
            I => \N__30032\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__30045\,
            I => \N__30027\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__30042\,
            I => \N__30027\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__30039\,
            I => \N__30024\
        );

    \I__6538\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30021\
        );

    \I__6537\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30018\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30013\
        );

    \I__6535\ : Span4Mux_h
    port map (
            O => \N__30027\,
            I => \N__30013\
        );

    \I__6534\ : Odrv4
    port map (
            O => \N__30024\,
            I => \POWERLED.N_396\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__30021\,
            I => \POWERLED.N_396\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__30018\,
            I => \POWERLED.N_396\
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__30013\,
            I => \POWERLED.N_396\
        );

    \I__6530\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29999\
        );

    \I__6529\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29996\
        );

    \I__6528\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29978\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__29999\,
            I => \N__29973\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__29996\,
            I => \N__29973\
        );

    \I__6525\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29970\
        );

    \I__6524\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29967\
        );

    \I__6523\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29958\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29958\
        );

    \I__6521\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29958\
        );

    \I__6520\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29958\
        );

    \I__6519\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29953\
        );

    \I__6518\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29953\
        );

    \I__6517\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29948\
        );

    \I__6516\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29948\
        );

    \I__6515\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29945\
        );

    \I__6514\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29940\
        );

    \I__6513\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29936\
        );

    \I__6512\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29931\
        );

    \I__6511\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29931\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__29978\,
            I => \N__29928\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__29973\,
            I => \N__29923\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29923\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__29967\,
            I => \N__29918\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29918\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__29953\,
            I => \N__29908\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__29948\,
            I => \N__29908\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__29945\,
            I => \N__29905\
        );

    \I__6502\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29900\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29900\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29897\
        );

    \I__6499\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29893\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__29936\,
            I => \N__29890\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29887\
        );

    \I__6496\ : Span4Mux_v
    port map (
            O => \N__29928\,
            I => \N__29880\
        );

    \I__6495\ : Span4Mux_v
    port map (
            O => \N__29923\,
            I => \N__29880\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__29918\,
            I => \N__29880\
        );

    \I__6493\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29875\
        );

    \I__6492\ : InMux
    port map (
            O => \N__29916\,
            I => \N__29875\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29915\,
            I => \N__29872\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29867\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29867\
        );

    \I__6488\ : Span4Mux_h
    port map (
            O => \N__29908\,
            I => \N__29864\
        );

    \I__6487\ : Span4Mux_v
    port map (
            O => \N__29905\,
            I => \N__29857\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29857\
        );

    \I__6485\ : Span4Mux_h
    port map (
            O => \N__29897\,
            I => \N__29857\
        );

    \I__6484\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29854\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__29893\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6482\ : Odrv4
    port map (
            O => \N__29890\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6481\ : Odrv12
    port map (
            O => \N__29887\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6480\ : Odrv4
    port map (
            O => \N__29880\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__29875\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__29872\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__29867\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__29864\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__29857\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__29854\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__29833\,
            I => \POWERLED.count_clk_en_2_cascade_\
        );

    \I__6472\ : CascadeMux
    port map (
            O => \N__29830\,
            I => \N__29822\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__29829\,
            I => \N__29817\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__29828\,
            I => \N__29813\
        );

    \I__6469\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29803\
        );

    \I__6468\ : IoInMux
    port map (
            O => \N__29826\,
            I => \N__29800\
        );

    \I__6467\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29797\
        );

    \I__6466\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29790\
        );

    \I__6465\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29790\
        );

    \I__6464\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29790\
        );

    \I__6463\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29781\
        );

    \I__6462\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29781\
        );

    \I__6461\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29781\
        );

    \I__6460\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29781\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__29811\,
            I => \N__29775\
        );

    \I__6458\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29763\
        );

    \I__6457\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29763\
        );

    \I__6456\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29763\
        );

    \I__6455\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29763\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__29806\,
            I => \N__29760\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29755\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__29800\,
            I => \N__29752\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__29797\,
            I => \N__29745\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__29790\,
            I => \N__29745\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__29781\,
            I => \N__29745\
        );

    \I__6448\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29738\
        );

    \I__6447\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29738\
        );

    \I__6446\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29735\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29728\
        );

    \I__6444\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29728\
        );

    \I__6443\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29728\
        );

    \I__6442\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29725\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__29763\,
            I => \N__29722\
        );

    \I__6440\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29717\
        );

    \I__6439\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29717\
        );

    \I__6438\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29714\
        );

    \I__6437\ : Span4Mux_v
    port map (
            O => \N__29755\,
            I => \N__29708\
        );

    \I__6436\ : Span4Mux_s3_h
    port map (
            O => \N__29752\,
            I => \N__29705\
        );

    \I__6435\ : Span4Mux_v
    port map (
            O => \N__29745\,
            I => \N__29702\
        );

    \I__6434\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29697\
        );

    \I__6433\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29697\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29738\,
            I => \N__29694\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29735\,
            I => \N__29689\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__29728\,
            I => \N__29689\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__29725\,
            I => \N__29682\
        );

    \I__6428\ : Span4Mux_h
    port map (
            O => \N__29722\,
            I => \N__29682\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__29717\,
            I => \N__29682\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29679\
        );

    \I__6425\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29675\
        );

    \I__6424\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29672\
        );

    \I__6423\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29669\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__29708\,
            I => \N__29664\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__29705\,
            I => \N__29664\
        );

    \I__6420\ : Span4Mux_v
    port map (
            O => \N__29702\,
            I => \N__29661\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__29697\,
            I => \N__29658\
        );

    \I__6418\ : Span4Mux_v
    port map (
            O => \N__29694\,
            I => \N__29649\
        );

    \I__6417\ : Span4Mux_h
    port map (
            O => \N__29689\,
            I => \N__29649\
        );

    \I__6416\ : Span4Mux_v
    port map (
            O => \N__29682\,
            I => \N__29649\
        );

    \I__6415\ : Span4Mux_h
    port map (
            O => \N__29679\,
            I => \N__29649\
        );

    \I__6414\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29646\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__29675\,
            I => \N__29643\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__29672\,
            I => \G_155\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__29669\,
            I => \G_155\
        );

    \I__6410\ : Odrv4
    port map (
            O => \N__29664\,
            I => \G_155\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__29661\,
            I => \G_155\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__29658\,
            I => \G_155\
        );

    \I__6407\ : Odrv4
    port map (
            O => \N__29649\,
            I => \G_155\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__29646\,
            I => \G_155\
        );

    \I__6405\ : Odrv12
    port map (
            O => \N__29643\,
            I => \G_155\
        );

    \I__6404\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29622\
        );

    \I__6403\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29617\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29614\
        );

    \I__6401\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29611\
        );

    \I__6400\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29608\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__29617\,
            I => \N__29605\
        );

    \I__6398\ : Span4Mux_h
    port map (
            O => \N__29614\,
            I => \N__29602\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__29611\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__29608\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__29605\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__29602\,
            I => \POWERLED.func_state_RNI_2Z0Z_1\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__29593\,
            I => \N__29584\
        );

    \I__6392\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29575\
        );

    \I__6391\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29575\
        );

    \I__6390\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29575\
        );

    \I__6389\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29570\
        );

    \I__6388\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29567\
        );

    \I__6387\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29564\
        );

    \I__6386\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29557\
        );

    \I__6385\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29557\
        );

    \I__6384\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29557\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__29575\,
            I => \N__29554\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__29574\,
            I => \N__29551\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__29573\,
            I => \N__29548\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29545\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29536\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__29564\,
            I => \N__29536\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__29557\,
            I => \N__29536\
        );

    \I__6376\ : Span4Mux_s3_h
    port map (
            O => \N__29554\,
            I => \N__29536\
        );

    \I__6375\ : InMux
    port map (
            O => \N__29551\,
            I => \N__29533\
        );

    \I__6374\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29530\
        );

    \I__6373\ : Span4Mux_v
    port map (
            O => \N__29545\,
            I => \N__29525\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__29536\,
            I => \N__29525\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__29533\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__29530\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__29525\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6368\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29515\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__29515\,
            I => \POWERLED.N_176\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__29512\,
            I => \POWERLED.N_176_cascade_\
        );

    \I__6365\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29501\
        );

    \I__6363\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29496\
        );

    \I__6362\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29496\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__29501\,
            I => \N__29491\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__29496\,
            I => \N__29491\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__29491\,
            I => \POWERLED.N_2218_i\
        );

    \I__6358\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29485\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__29485\,
            I => \N__29482\
        );

    \I__6356\ : Span4Mux_v
    port map (
            O => \N__29482\,
            I => \N__29475\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__29481\,
            I => \N__29470\
        );

    \I__6354\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29466\
        );

    \I__6353\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29461\
        );

    \I__6352\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29461\
        );

    \I__6351\ : IoSpan4Mux
    port map (
            O => \N__29475\,
            I => \N__29455\
        );

    \I__6350\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29452\
        );

    \I__6349\ : CascadeMux
    port map (
            O => \N__29473\,
            I => \N__29448\
        );

    \I__6348\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29442\
        );

    \I__6347\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29442\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__29466\,
            I => \N__29439\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__29461\,
            I => \N__29436\
        );

    \I__6344\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29433\
        );

    \I__6343\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29430\
        );

    \I__6342\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29427\
        );

    \I__6341\ : Span4Mux_s3_h
    port map (
            O => \N__29455\,
            I => \N__29419\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__29452\,
            I => \N__29419\
        );

    \I__6339\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29412\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29412\
        );

    \I__6337\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29412\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29409\
        );

    \I__6335\ : Span4Mux_h
    port map (
            O => \N__29439\,
            I => \N__29398\
        );

    \I__6334\ : Span4Mux_s3_v
    port map (
            O => \N__29436\,
            I => \N__29398\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__29433\,
            I => \N__29398\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29398\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29398\
        );

    \I__6330\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29393\
        );

    \I__6329\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29393\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29389\
        );

    \I__6327\ : Span4Mux_h
    port map (
            O => \N__29419\,
            I => \N__29384\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29384\
        );

    \I__6325\ : Span4Mux_v
    port map (
            O => \N__29409\,
            I => \N__29375\
        );

    \I__6324\ : Span4Mux_v
    port map (
            O => \N__29398\,
            I => \N__29375\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29375\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__29392\,
            I => \N__29372\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29389\,
            I => \N__29366\
        );

    \I__6320\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29366\
        );

    \I__6319\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29361\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29361\
        );

    \I__6317\ : Sp12to4
    port map (
            O => \N__29375\,
            I => \N__29358\
        );

    \I__6316\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29353\
        );

    \I__6315\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29353\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__29366\,
            I => \POWERLED.N_2216_i\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__29361\,
            I => \POWERLED.N_2216_i\
        );

    \I__6312\ : Odrv12
    port map (
            O => \N__29358\,
            I => \POWERLED.N_2216_i\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__29353\,
            I => \POWERLED.N_2216_i\
        );

    \I__6310\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29341\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__29341\,
            I => \N__29338\
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__29338\,
            I => \POWERLED.N_27\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__29335\,
            I => \N__29326\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \N__29323\
        );

    \I__6305\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29319\
        );

    \I__6304\ : InMux
    port map (
            O => \N__29332\,
            I => \N__29308\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29308\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__29330\,
            I => \N__29298\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__29329\,
            I => \N__29295\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29291\
        );

    \I__6299\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29288\
        );

    \I__6298\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29285\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__29319\,
            I => \N__29282\
        );

    \I__6296\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29279\
        );

    \I__6295\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29272\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29272\
        );

    \I__6293\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29272\
        );

    \I__6292\ : InMux
    port map (
            O => \N__29314\,
            I => \N__29269\
        );

    \I__6291\ : InMux
    port map (
            O => \N__29313\,
            I => \N__29266\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29263\
        );

    \I__6289\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29256\
        );

    \I__6288\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29256\
        );

    \I__6287\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29256\
        );

    \I__6286\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29253\
        );

    \I__6285\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29250\
        );

    \I__6284\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29247\
        );

    \I__6283\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29241\
        );

    \I__6282\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29241\
        );

    \I__6281\ : InMux
    port map (
            O => \N__29295\,
            I => \N__29236\
        );

    \I__6280\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29236\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__29291\,
            I => \N__29229\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29288\,
            I => \N__29229\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29229\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__29282\,
            I => \N__29224\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29224\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__29272\,
            I => \N__29220\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__29269\,
            I => \N__29215\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__29266\,
            I => \N__29215\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__29263\,
            I => \N__29210\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29210\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29203\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29203\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__29247\,
            I => \N__29203\
        );

    \I__6266\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29199\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__29241\,
            I => \N__29196\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29193\
        );

    \I__6263\ : Span4Mux_v
    port map (
            O => \N__29229\,
            I => \N__29188\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__29224\,
            I => \N__29188\
        );

    \I__6261\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29185\
        );

    \I__6260\ : Span4Mux_h
    port map (
            O => \N__29220\,
            I => \N__29176\
        );

    \I__6259\ : Span4Mux_v
    port map (
            O => \N__29215\,
            I => \N__29176\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__29210\,
            I => \N__29176\
        );

    \I__6257\ : Span4Mux_v
    port map (
            O => \N__29203\,
            I => \N__29176\
        );

    \I__6256\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29173\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__29199\,
            I => \N__29166\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__29196\,
            I => \N__29166\
        );

    \I__6253\ : Span4Mux_s2_h
    port map (
            O => \N__29193\,
            I => \N__29166\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__29188\,
            I => \POWERLED.func_state\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__29185\,
            I => \POWERLED.func_state\
        );

    \I__6250\ : Odrv4
    port map (
            O => \N__29176\,
            I => \POWERLED.func_state\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__29173\,
            I => \POWERLED.func_state\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__29166\,
            I => \POWERLED.func_state\
        );

    \I__6247\ : InMux
    port map (
            O => \N__29155\,
            I => \N__29152\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__29152\,
            I => \N__29149\
        );

    \I__6245\ : Span4Mux_s1_h
    port map (
            O => \N__29149\,
            I => \N__29146\
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__29146\,
            I => \POWERLED.N_219\
        );

    \I__6243\ : IoInMux
    port map (
            O => \N__29143\,
            I => \N__29140\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__29140\,
            I => \N__29137\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__29137\,
            I => vpp_en
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__29134\,
            I => \VPP_VDDQ.N_64_cascade_\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__29131\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\
        );

    \I__6238\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29122\
        );

    \I__6237\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29122\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__29122\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__29119\,
            I => \POWERLED.count_clk_RNIZ0Z_1_cascade_\
        );

    \I__6234\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29110\
        );

    \I__6233\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29110\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__29110\,
            I => \N__29106\
        );

    \I__6231\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29103\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__29106\,
            I => \N__29100\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__29103\,
            I => \POWERLED.count_clk_RNI_0Z0Z_1\
        );

    \I__6228\ : Odrv4
    port map (
            O => \N__29100\,
            I => \POWERLED.count_clk_RNI_0Z0Z_1\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__29095\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_a2_0_0_cascade_\
        );

    \I__6226\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29089\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29086\
        );

    \I__6224\ : Span4Mux_s1_h
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__6223\ : Span4Mux_v
    port map (
            O => \N__29083\,
            I => \N__29080\
        );

    \I__6222\ : Odrv4
    port map (
            O => \N__29080\,
            I => \POWERLED.N_285\
        );

    \I__6221\ : InMux
    port map (
            O => \N__29077\,
            I => \N__29074\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__29074\,
            I => \POWERLED.N_177\
        );

    \I__6219\ : CascadeMux
    port map (
            O => \N__29071\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_1_cascade_\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__29068\,
            I => \N__29063\
        );

    \I__6217\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29055\
        );

    \I__6216\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29055\
        );

    \I__6215\ : InMux
    port map (
            O => \N__29063\,
            I => \N__29052\
        );

    \I__6214\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29044\
        );

    \I__6213\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29044\
        );

    \I__6212\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29041\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__29055\,
            I => \N__29037\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__29052\,
            I => \N__29034\
        );

    \I__6209\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29031\
        );

    \I__6208\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29026\
        );

    \I__6207\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29026\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__29044\,
            I => \N__29021\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__29041\,
            I => \N__29021\
        );

    \I__6204\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29018\
        );

    \I__6203\ : Span4Mux_v
    port map (
            O => \N__29037\,
            I => \N__29011\
        );

    \I__6202\ : Span4Mux_h
    port map (
            O => \N__29034\,
            I => \N__29011\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__29031\,
            I => \N__29011\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__29026\,
            I => \N__29008\
        );

    \I__6199\ : Span4Mux_v
    port map (
            O => \N__29021\,
            I => \N__29003\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__29018\,
            I => \N__29003\
        );

    \I__6197\ : Span4Mux_v
    port map (
            O => \N__29011\,
            I => \N__29000\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__29008\,
            I => \N__28995\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__29003\,
            I => \N__28995\
        );

    \I__6194\ : Span4Mux_v
    port map (
            O => \N__29000\,
            I => \N__28992\
        );

    \I__6193\ : Span4Mux_v
    port map (
            O => \N__28995\,
            I => \N__28989\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__28992\,
            I => gpio_fpga_soc_4
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__28989\,
            I => gpio_fpga_soc_4
        );

    \I__6190\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28974\
        );

    \I__6189\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28974\
        );

    \I__6188\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28971\
        );

    \I__6187\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28966\
        );

    \I__6186\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28966\
        );

    \I__6185\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28963\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28950\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28950\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28945\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28945\
        );

    \I__6180\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28942\
        );

    \I__6179\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28932\
        );

    \I__6178\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28932\
        );

    \I__6177\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28932\
        );

    \I__6176\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28932\
        );

    \I__6175\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28927\
        );

    \I__6174\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28927\
        );

    \I__6173\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28924\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__28950\,
            I => \N__28917\
        );

    \I__6171\ : Span4Mux_h
    port map (
            O => \N__28945\,
            I => \N__28917\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28917\
        );

    \I__6169\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28914\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__28932\,
            I => \N__28905\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28902\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__28924\,
            I => \N__28898\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__28917\,
            I => \N__28893\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__28914\,
            I => \N__28893\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28886\
        );

    \I__6162\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28886\
        );

    \I__6161\ : InMux
    port map (
            O => \N__28911\,
            I => \N__28886\
        );

    \I__6160\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28882\
        );

    \I__6159\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28879\
        );

    \I__6158\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28876\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__28905\,
            I => \N__28871\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__28902\,
            I => \N__28871\
        );

    \I__6155\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28868\
        );

    \I__6154\ : Span4Mux_v
    port map (
            O => \N__28898\,
            I => \N__28861\
        );

    \I__6153\ : Span4Mux_v
    port map (
            O => \N__28893\,
            I => \N__28861\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28861\
        );

    \I__6151\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28858\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__28882\,
            I => \N__28847\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__28879\,
            I => \N__28847\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__28876\,
            I => \N__28847\
        );

    \I__6147\ : Sp12to4
    port map (
            O => \N__28871\,
            I => \N__28847\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__28868\,
            I => \N__28847\
        );

    \I__6145\ : Span4Mux_h
    port map (
            O => \N__28861\,
            I => \N__28842\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28842\
        );

    \I__6143\ : Span12Mux_s8_h
    port map (
            O => \N__28847\,
            I => \N__28839\
        );

    \I__6142\ : IoSpan4Mux
    port map (
            O => \N__28842\,
            I => \N__28836\
        );

    \I__6141\ : Odrv12
    port map (
            O => \N__28839\,
            I => slp_s4n
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__28836\,
            I => slp_s4n
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__28831\,
            I => \POWERLED.un1_func_state25_4_i_a2_0_cascade_\
        );

    \I__6138\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28824\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__28827\,
            I => \N__28821\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28817\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28814\
        );

    \I__6134\ : CascadeMux
    port map (
            O => \N__28820\,
            I => \N__28811\
        );

    \I__6133\ : Span4Mux_s3_h
    port map (
            O => \N__28817\,
            I => \N__28808\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28805\
        );

    \I__6131\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28802\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__28808\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__28805\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28802\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0\
        );

    \I__6127\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28792\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__28792\,
            I => \POWERLED.N_291\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \POWERLED.count_clk_en_0_cascade_\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__28786\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__28783\,
            I => \POWERLED.count_clkZ0Z_0_cascade_\
        );

    \I__6122\ : CascadeMux
    port map (
            O => \N__28780\,
            I => \POWERLED.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__6121\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28774\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__28774\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__6119\ : CascadeMux
    port map (
            O => \N__28771\,
            I => \N__28768\
        );

    \I__6118\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28765\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__28765\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28759\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__28759\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__6114\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28750\
        );

    \I__6113\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28750\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__6111\ : Span4Mux_h
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__28744\,
            I => \POWERLED.count_clk_RNIZ0Z_1\
        );

    \I__6109\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28738\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__28738\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__6107\ : CascadeMux
    port map (
            O => \N__28735\,
            I => \POWERLED.count_clkZ0Z_14_cascade_\
        );

    \I__6106\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28729\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__28729\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28723\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__28723\,
            I => \POWERLED.count_clk_0_14\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__28720\,
            I => \VPP_VDDQ.count_2_1_7_cascade_\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28713\
        );

    \I__6100\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28710\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__28713\,
            I => \N__28707\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__28710\,
            I => \N__28704\
        );

    \I__6097\ : Span4Mux_v
    port map (
            O => \N__28707\,
            I => \N__28701\
        );

    \I__6096\ : Span4Mux_s2_h
    port map (
            O => \N__28704\,
            I => \N__28698\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__28701\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__28698\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__28693\,
            I => \VPP_VDDQ.un9_clk_100khz_7_cascade_\
        );

    \I__6092\ : InMux
    port map (
            O => \N__28690\,
            I => \N__28686\
        );

    \I__6091\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28683\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__28686\,
            I => \N__28678\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__28683\,
            I => \N__28678\
        );

    \I__6088\ : Span4Mux_v
    port map (
            O => \N__28678\,
            I => \N__28675\
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__28675\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__6086\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28669\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__28669\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__6084\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28663\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28660\
        );

    \I__6082\ : Odrv4
    port map (
            O => \N__28660\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__6081\ : InMux
    port map (
            O => \N__28657\,
            I => \N__28651\
        );

    \I__6080\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28651\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__28648\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\
        );

    \I__6077\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28639\
        );

    \I__6076\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28639\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__28639\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__28636\,
            I => \VPP_VDDQ.count_2_1_0_cascade_\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__28633\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28627\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__28627\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28624\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28614\
        );

    \I__6067\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28611\
        );

    \I__6066\ : Span4Mux_s3_h
    port map (
            O => \N__28614\,
            I => \N__28608\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__28611\,
            I => \N__28605\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__28608\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__6063\ : Odrv12
    port map (
            O => \N__28605\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__28600\,
            I => \N__28596\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__28599\,
            I => \N__28593\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28588\
        );

    \I__6059\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28588\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__28588\,
            I => \N__28585\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__28585\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\
        );

    \I__6056\ : InMux
    port map (
            O => \N__28582\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__28579\,
            I => \N__28575\
        );

    \I__6054\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28570\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28570\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28570\,
            I => \N__28567\
        );

    \I__6051\ : Span4Mux_v
    port map (
            O => \N__28567\,
            I => \N__28564\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__28564\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\
        );

    \I__6049\ : InMux
    port map (
            O => \N__28561\,
            I => \bfn_11_7_0_\
        );

    \I__6048\ : CascadeMux
    port map (
            O => \N__28558\,
            I => \N__28554\
        );

    \I__6047\ : CascadeMux
    port map (
            O => \N__28557\,
            I => \N__28551\
        );

    \I__6046\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28548\
        );

    \I__6045\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28545\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28542\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28539\
        );

    \I__6042\ : Span4Mux_v
    port map (
            O => \N__28542\,
            I => \N__28536\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__28539\,
            I => \N__28533\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__28536\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__28533\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\
        );

    \I__6038\ : InMux
    port map (
            O => \N__28528\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__6037\ : InMux
    port map (
            O => \N__28525\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28522\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28519\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28516\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__6033\ : InMux
    port map (
            O => \N__28513\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__28510\,
            I => \N__28506\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28501\
        );

    \I__6030\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28501\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__28501\,
            I => \N__28498\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__28498\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__28495\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\
        );

    \I__6026\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__28489\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__6024\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28483\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__28483\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__6022\ : InMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__28477\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__28474\,
            I => \N__28470\
        );

    \I__6019\ : InMux
    port map (
            O => \N__28473\,
            I => \N__28465\
        );

    \I__6018\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28465\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__28465\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\
        );

    \I__6016\ : InMux
    port map (
            O => \N__28462\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__6015\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28455\
        );

    \I__6014\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28452\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__28455\,
            I => \N__28449\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__28452\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__28449\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__6010\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28440\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28437\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__28440\,
            I => \N__28434\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__28437\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__6006\ : Odrv4
    port map (
            O => \N__28434\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__6005\ : InMux
    port map (
            O => \N__28429\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__6004\ : InMux
    port map (
            O => \N__28426\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__6003\ : InMux
    port map (
            O => \N__28423\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__6002\ : InMux
    port map (
            O => \N__28420\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__28417\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__6000\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28411\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__28411\,
            I => \VPP_VDDQ.curr_state_2_0_1\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__28408\,
            I => \VPP_VDDQ.N_55_cascade_\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__28405\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__28402\,
            I => \VPP_VDDQ.count_2_1_3_cascade_\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__28399\,
            I => \VPP_VDDQ.count_2_1_2_cascade_\
        );

    \I__5994\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28393\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__28393\,
            I => \VPP_VDDQ.count_2_0_2\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__28390\,
            I => \VPP_VDDQ.count_2Z0Z_2_cascade_\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__28387\,
            I => \G_1939_cascade_\
        );

    \I__5990\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28380\
        );

    \I__5989\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28377\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__28380\,
            I => \N__28373\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__28377\,
            I => \N__28370\
        );

    \I__5986\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28367\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__28373\,
            I => \N__28362\
        );

    \I__5984\ : Span4Mux_s2_h
    port map (
            O => \N__28370\,
            I => \N__28362\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__28367\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__28362\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__5981\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28354\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__28354\,
            I => \N__28350\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28347\
        );

    \I__5978\ : Span4Mux_s2_v
    port map (
            O => \N__28350\,
            I => \N__28344\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__28347\,
            I => \N_218\
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__28344\,
            I => \N_218\
        );

    \I__5975\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__28336\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__5973\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28327\
        );

    \I__5972\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28327\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__28327\,
            I => \N__28323\
        );

    \I__5970\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28320\
        );

    \I__5969\ : Span4Mux_h
    port map (
            O => \N__28323\,
            I => \N__28317\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__28320\,
            I => \G_1939\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__28317\,
            I => \G_1939\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__28312\,
            I => \N_218_cascade_\
        );

    \I__5965\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28306\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__28306\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__28303\,
            I => \PCH_PWRGD.curr_state_0_1_cascade_\
        );

    \I__5962\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28294\
        );

    \I__5961\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28294\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__28294\,
            I => \N__28291\
        );

    \I__5959\ : Span4Mux_s2_v
    port map (
            O => \N__28291\,
            I => \N__28287\
        );

    \I__5958\ : InMux
    port map (
            O => \N__28290\,
            I => \N__28284\
        );

    \I__5957\ : Odrv4
    port map (
            O => \N__28287\,
            I => \PCH_PWRGD.N_2190_i\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__28284\,
            I => \PCH_PWRGD.N_2190_i\
        );

    \I__5955\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28275\
        );

    \I__5954\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28272\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__28275\,
            I => \N__28267\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__28272\,
            I => \N__28264\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28261\
        );

    \I__5950\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28258\
        );

    \I__5949\ : Span4Mux_s3_v
    port map (
            O => \N__28267\,
            I => \N__28253\
        );

    \I__5948\ : Span4Mux_s3_v
    port map (
            O => \N__28264\,
            I => \N__28253\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__28261\,
            I => \PCH_PWRGD.N_2171_i\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__28258\,
            I => \PCH_PWRGD.N_2171_i\
        );

    \I__5945\ : Odrv4
    port map (
            O => \N__28253\,
            I => \PCH_PWRGD.N_2171_i\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__28246\,
            I => \PCH_PWRGD.N_2190_i_cascade_\
        );

    \I__5943\ : SRMux
    port map (
            O => \N__28243\,
            I => \N__28236\
        );

    \I__5942\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28229\
        );

    \I__5941\ : SRMux
    port map (
            O => \N__28241\,
            I => \N__28229\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__28240\,
            I => \N__28219\
        );

    \I__5939\ : CascadeMux
    port map (
            O => \N__28239\,
            I => \N__28213\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__28236\,
            I => \N__28200\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__28235\,
            I => \N__28197\
        );

    \I__5936\ : CascadeMux
    port map (
            O => \N__28234\,
            I => \N__28194\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__28229\,
            I => \N__28190\
        );

    \I__5934\ : SRMux
    port map (
            O => \N__28228\,
            I => \N__28187\
        );

    \I__5933\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28182\
        );

    \I__5932\ : SRMux
    port map (
            O => \N__28226\,
            I => \N__28182\
        );

    \I__5931\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28179\
        );

    \I__5930\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28174\
        );

    \I__5929\ : InMux
    port map (
            O => \N__28223\,
            I => \N__28174\
        );

    \I__5928\ : InMux
    port map (
            O => \N__28222\,
            I => \N__28171\
        );

    \I__5927\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28163\
        );

    \I__5926\ : InMux
    port map (
            O => \N__28218\,
            I => \N__28160\
        );

    \I__5925\ : SRMux
    port map (
            O => \N__28217\,
            I => \N__28151\
        );

    \I__5924\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28151\
        );

    \I__5923\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28151\
        );

    \I__5922\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28151\
        );

    \I__5921\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28140\
        );

    \I__5920\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28140\
        );

    \I__5919\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28140\
        );

    \I__5918\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28140\
        );

    \I__5917\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28140\
        );

    \I__5916\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28131\
        );

    \I__5915\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28131\
        );

    \I__5914\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28131\
        );

    \I__5913\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28131\
        );

    \I__5912\ : Span4Mux_s3_v
    port map (
            O => \N__28200\,
            I => \N__28128\
        );

    \I__5911\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28121\
        );

    \I__5910\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28121\
        );

    \I__5909\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28121\
        );

    \I__5908\ : Span4Mux_v
    port map (
            O => \N__28190\,
            I => \N__28114\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__28187\,
            I => \N__28114\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__28182\,
            I => \N__28114\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__28179\,
            I => \N__28107\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__28174\,
            I => \N__28107\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28107\
        );

    \I__5902\ : SRMux
    port map (
            O => \N__28170\,
            I => \N__28098\
        );

    \I__5901\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28098\
        );

    \I__5900\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28098\
        );

    \I__5899\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28098\
        );

    \I__5898\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28095\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__28163\,
            I => \N__28084\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__28160\,
            I => \N__28084\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28084\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__28140\,
            I => \N__28084\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__28131\,
            I => \N__28084\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__28128\,
            I => \N__28080\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__28121\,
            I => \N__28075\
        );

    \I__5890\ : Span4Mux_h
    port map (
            O => \N__28114\,
            I => \N__28075\
        );

    \I__5889\ : Span4Mux_s2_v
    port map (
            O => \N__28107\,
            I => \N__28072\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__28098\,
            I => \N__28069\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__28095\,
            I => \N__28064\
        );

    \I__5886\ : Span4Mux_s2_v
    port map (
            O => \N__28084\,
            I => \N__28064\
        );

    \I__5885\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28061\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__28080\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__28075\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__28072\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__28069\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__5880\ : Odrv4
    port map (
            O => \N__28064\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__28061\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__5878\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28045\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__28045\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__28042\,
            I => \VPP_VDDQ.N_53_cascade_\
        );

    \I__5875\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28036\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__28036\,
            I => \PCH_PWRGD.count_rst_7\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__28033\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__5872\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28027\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__28027\,
            I => \PCH_PWRGD.count_1_i_a2_5_0\
        );

    \I__5870\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28018\
        );

    \I__5869\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28018\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__28018\,
            I => \N__28015\
        );

    \I__5867\ : Span4Mux_s3_h
    port map (
            O => \N__28015\,
            I => \N__28012\
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__28012\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__28009\,
            I => \N__28006\
        );

    \I__5864\ : InMux
    port map (
            O => \N__28006\,
            I => \N__28003\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__28003\,
            I => \N__27998\
        );

    \I__5862\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27993\
        );

    \I__5861\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27993\
        );

    \I__5860\ : Span4Mux_s1_v
    port map (
            O => \N__27998\,
            I => \N__27990\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__27993\,
            I => \PCH_PWRGD.un2_count_1_axb_7\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__27990\,
            I => \PCH_PWRGD.un2_count_1_axb_7\
        );

    \I__5857\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27979\
        );

    \I__5856\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27979\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__27979\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__5854\ : CascadeMux
    port map (
            O => \N__27976\,
            I => \PCH_PWRGD.count_rst_9_cascade_\
        );

    \I__5853\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27970\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__27970\,
            I => \N__27967\
        );

    \I__5851\ : Span4Mux_s1_v
    port map (
            O => \N__27967\,
            I => \N__27962\
        );

    \I__5850\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27957\
        );

    \I__5849\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27957\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__27962\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__27957\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__5846\ : CascadeMux
    port map (
            O => \N__27952\,
            I => \N__27949\
        );

    \I__5845\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27943\
        );

    \I__5844\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27943\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__27943\,
            I => \N__27940\
        );

    \I__5842\ : Span4Mux_v
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__27937\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__27934\,
            I => \PCH_PWRGD.countZ0Z_5_cascade_\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27928\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__27928\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__5837\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27922\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__27922\,
            I => \N__27918\
        );

    \I__5835\ : InMux
    port map (
            O => \N__27921\,
            I => \N__27915\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__27918\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__27915\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__27910\,
            I => \N__27906\
        );

    \I__5831\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27902\
        );

    \I__5830\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27899\
        );

    \I__5829\ : CascadeMux
    port map (
            O => \N__27905\,
            I => \N__27895\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27890\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27890\
        );

    \I__5826\ : CascadeMux
    port map (
            O => \N__27898\,
            I => \N__27887\
        );

    \I__5825\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27884\
        );

    \I__5824\ : Span4Mux_s2_v
    port map (
            O => \N__27890\,
            I => \N__27881\
        );

    \I__5823\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27878\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__27884\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__27881\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__27878\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__5819\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27868\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__27862\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__5815\ : CEMux
    port map (
            O => \N__27859\,
            I => \N__27853\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__27858\,
            I => \N__27846\
        );

    \I__5813\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27839\
        );

    \I__5812\ : CEMux
    port map (
            O => \N__27856\,
            I => \N__27839\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27853\,
            I => \N__27835\
        );

    \I__5810\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27822\
        );

    \I__5809\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27822\
        );

    \I__5808\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27822\
        );

    \I__5807\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27822\
        );

    \I__5806\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27815\
        );

    \I__5805\ : CEMux
    port map (
            O => \N__27845\,
            I => \N__27815\
        );

    \I__5804\ : CEMux
    port map (
            O => \N__27844\,
            I => \N__27812\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__27839\,
            I => \N__27799\
        );

    \I__5802\ : CEMux
    port map (
            O => \N__27838\,
            I => \N__27796\
        );

    \I__5801\ : Span4Mux_s1_v
    port map (
            O => \N__27835\,
            I => \N__27793\
        );

    \I__5800\ : CEMux
    port map (
            O => \N__27834\,
            I => \N__27784\
        );

    \I__5799\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27784\
        );

    \I__5798\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27784\
        );

    \I__5797\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27784\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27781\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27776\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27773\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27770\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__27812\,
            I => \N__27767\
        );

    \I__5791\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27764\
        );

    \I__5790\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27755\
        );

    \I__5789\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27755\
        );

    \I__5788\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27755\
        );

    \I__5787\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27755\
        );

    \I__5786\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27750\
        );

    \I__5785\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27750\
        );

    \I__5784\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27743\
        );

    \I__5783\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27743\
        );

    \I__5782\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27743\
        );

    \I__5781\ : Span4Mux_s1_h
    port map (
            O => \N__27799\,
            I => \N__27732\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27732\
        );

    \I__5779\ : Span4Mux_s1_h
    port map (
            O => \N__27793\,
            I => \N__27732\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27732\
        );

    \I__5777\ : Span4Mux_s1_v
    port map (
            O => \N__27781\,
            I => \N__27732\
        );

    \I__5776\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27727\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27779\,
            I => \N__27727\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__27776\,
            I => \N__27722\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__27773\,
            I => \N__27722\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__27770\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__27767\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__27764\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__27755\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__27750\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__27743\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__27732\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__27727\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5764\ : Odrv12
    port map (
            O => \N__27722\,
            I => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27686\
        );

    \I__5762\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27686\
        );

    \I__5761\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27674\
        );

    \I__5760\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27674\
        );

    \I__5759\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27674\
        );

    \I__5758\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27674\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27697\,
            I => \N__27674\
        );

    \I__5756\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27671\
        );

    \I__5755\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27659\
        );

    \I__5754\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27659\
        );

    \I__5753\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27659\
        );

    \I__5752\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27659\
        );

    \I__5751\ : InMux
    port map (
            O => \N__27691\,
            I => \N__27659\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27656\
        );

    \I__5749\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27653\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__27674\,
            I => \N__27648\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27671\,
            I => \N__27648\
        );

    \I__5746\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27645\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27659\,
            I => \N__27642\
        );

    \I__5744\ : Span4Mux_s2_v
    port map (
            O => \N__27656\,
            I => \N__27633\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__27653\,
            I => \N__27633\
        );

    \I__5742\ : Span4Mux_s2_v
    port map (
            O => \N__27648\,
            I => \N__27633\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27633\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__27642\,
            I => \PCH_PWRGD.N_364\
        );

    \I__5739\ : Odrv4
    port map (
            O => \N__27633\,
            I => \PCH_PWRGD.N_364\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__27628\,
            I => \N__27625\
        );

    \I__5737\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27621\
        );

    \I__5736\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27618\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27615\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__27618\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__5733\ : Odrv12
    port map (
            O => \N__27615\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__27610\,
            I => \PCH_PWRGD.un2_count_1_axb_1_cascade_\
        );

    \I__5731\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27600\
        );

    \I__5730\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27600\
        );

    \I__5729\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27597\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27594\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__27597\,
            I => \N__27591\
        );

    \I__5726\ : Span4Mux_s2_h
    port map (
            O => \N__27594\,
            I => \N__27588\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__27591\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__27588\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27583\,
            I => \N__27580\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__27580\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27571\
        );

    \I__5720\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27571\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__27571\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__27568\,
            I => \PCH_PWRGD.count_rst_13_cascade_\
        );

    \I__5717\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27562\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__27562\,
            I => \N__27559\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__27559\,
            I => \PCH_PWRGD.count_1_i_a2_6_0\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__27556\,
            I => \PCH_PWRGD.count_1_i_a2_3_0_cascade_\
        );

    \I__5713\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27546\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27546\
        );

    \I__5711\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27543\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__27546\,
            I => \N__27540\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__27543\,
            I => \N__27537\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__27540\,
            I => \N__27534\
        );

    \I__5707\ : Span4Mux_h
    port map (
            O => \N__27537\,
            I => \N__27531\
        );

    \I__5706\ : Odrv4
    port map (
            O => \N__27534\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__27531\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__27526\,
            I => \N__27522\
        );

    \I__5703\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27519\
        );

    \I__5702\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27516\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__27519\,
            I => \N__27513\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__27516\,
            I => \N__27508\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__27513\,
            I => \N__27508\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__27508\,
            I => \PCH_PWRGD.un2_count_1_axb_9\
        );

    \I__5697\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27502\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__27502\,
            I => \N__27498\
        );

    \I__5695\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27495\
        );

    \I__5694\ : Span4Mux_s1_v
    port map (
            O => \N__27498\,
            I => \N__27492\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__27495\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__27492\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__27487\,
            I => \PCH_PWRGD.un2_count_1_axb_9_cascade_\
        );

    \I__5690\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27481\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__27481\,
            I => \PCH_PWRGD.count_rst_5\
        );

    \I__5688\ : InMux
    port map (
            O => \N__27478\,
            I => \N__27472\
        );

    \I__5687\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27472\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__27472\,
            I => \N__27469\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__27469\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__5684\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27461\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__27465\,
            I => \N__27458\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__27464\,
            I => \N__27455\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27452\
        );

    \I__5680\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27449\
        );

    \I__5679\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27446\
        );

    \I__5678\ : Odrv12
    port map (
            O => \N__27452\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__27449\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__27446\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__27439\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__5674\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27433\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__27433\,
            I => \PCH_PWRGD.count_1_i_a2_4_0\
        );

    \I__5672\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27425\
        );

    \I__5671\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27416\
        );

    \I__5670\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27413\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__27425\,
            I => \N__27408\
        );

    \I__5668\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27403\
        );

    \I__5667\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27403\
        );

    \I__5666\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27400\
        );

    \I__5665\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27397\
        );

    \I__5664\ : InMux
    port map (
            O => \N__27420\,
            I => \N__27392\
        );

    \I__5663\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27392\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27387\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__27413\,
            I => \N__27387\
        );

    \I__5660\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27384\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__27411\,
            I => \N__27381\
        );

    \I__5658\ : Span4Mux_v
    port map (
            O => \N__27408\,
            I => \N__27378\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__27403\,
            I => \N__27375\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27366\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__27397\,
            I => \N__27366\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__27392\,
            I => \N__27366\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__27387\,
            I => \N__27366\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27384\,
            I => \N__27363\
        );

    \I__5651\ : InMux
    port map (
            O => \N__27381\,
            I => \N__27360\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__27378\,
            I => \POWERLED.func_state_RNIZ0Z_1\
        );

    \I__5649\ : Odrv4
    port map (
            O => \N__27375\,
            I => \POWERLED.func_state_RNIZ0Z_1\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__27366\,
            I => \POWERLED.func_state_RNIZ0Z_1\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__27363\,
            I => \POWERLED.func_state_RNIZ0Z_1\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__27360\,
            I => \POWERLED.func_state_RNIZ0Z_1\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__27349\,
            I => \N__27342\
        );

    \I__5644\ : CascadeMux
    port map (
            O => \N__27348\,
            I => \N__27336\
        );

    \I__5643\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27326\
        );

    \I__5642\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27326\
        );

    \I__5641\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27326\
        );

    \I__5640\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27323\
        );

    \I__5639\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27320\
        );

    \I__5638\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27316\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__27339\,
            I => \N__27312\
        );

    \I__5636\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27307\
        );

    \I__5635\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27307\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__27334\,
            I => \N__27304\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__27333\,
            I => \N__27299\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27292\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27292\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27292\
        );

    \I__5629\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27289\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__27316\,
            I => \N__27286\
        );

    \I__5627\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27281\
        );

    \I__5626\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27281\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__27307\,
            I => \N__27278\
        );

    \I__5624\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27274\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27269\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27302\,
            I => \N__27269\
        );

    \I__5621\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27266\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__27292\,
            I => \N__27259\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27259\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__27286\,
            I => \N__27254\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27254\
        );

    \I__5616\ : Span4Mux_v
    port map (
            O => \N__27278\,
            I => \N__27251\
        );

    \I__5615\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27248\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__27274\,
            I => \N__27243\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__27269\,
            I => \N__27243\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27240\
        );

    \I__5611\ : InMux
    port map (
            O => \N__27265\,
            I => \N__27237\
        );

    \I__5610\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27234\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__27259\,
            I => \N__27231\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__27254\,
            I => \N__27228\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__27251\,
            I => \N__27223\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__27248\,
            I => \N__27223\
        );

    \I__5605\ : Span4Mux_v
    port map (
            O => \N__27243\,
            I => \N__27216\
        );

    \I__5604\ : Span4Mux_h
    port map (
            O => \N__27240\,
            I => \N__27216\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__27237\,
            I => \N__27216\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__27234\,
            I => \N__27213\
        );

    \I__5601\ : IoSpan4Mux
    port map (
            O => \N__27231\,
            I => \N__27210\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__27228\,
            I => \N__27207\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__27223\,
            I => \N__27204\
        );

    \I__5598\ : IoSpan4Mux
    port map (
            O => \N__27216\,
            I => \N__27201\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__27213\,
            I => \N__27198\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__27210\,
            I => slp_s3n
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__27207\,
            I => slp_s3n
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__27204\,
            I => slp_s3n
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__27201\,
            I => slp_s3n
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__27198\,
            I => slp_s3n
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__27187\,
            I => \POWERLED.un1_clk_100khz_51_and_i_a2_6_0_cascade_\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__27184\,
            I => \POWERLED.un1_clk_100khz_51_and_i_a2_6_sx_cascade_\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__27181\,
            I => \POWERLED.func_state_RNIPUGO_0Z0Z_1_cascade_\
        );

    \I__5588\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27175\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__27175\,
            I => \POWERLED.N_309_N\
        );

    \I__5586\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__27169\,
            I => \POWERLED.count_clk_RNI2O4A1Z0Z_10\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__27166\,
            I => \POWERLED.un1_clk_100khz_51_and_i_o2_4_1_cascade_\
        );

    \I__5583\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27155\
        );

    \I__5582\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27155\
        );

    \I__5581\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27146\
        );

    \I__5580\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27146\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__27155\,
            I => \N__27137\
        );

    \I__5578\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27134\
        );

    \I__5577\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27129\
        );

    \I__5576\ : InMux
    port map (
            O => \N__27152\,
            I => \N__27129\
        );

    \I__5575\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27126\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27123\
        );

    \I__5573\ : CascadeMux
    port map (
            O => \N__27145\,
            I => \N__27120\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__27144\,
            I => \N__27114\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__27143\,
            I => \N__27111\
        );

    \I__5570\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27105\
        );

    \I__5569\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27105\
        );

    \I__5568\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27102\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__27137\,
            I => \N__27097\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27097\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__27129\,
            I => \N__27094\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__27126\,
            I => \N__27089\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__27123\,
            I => \N__27089\
        );

    \I__5562\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27086\
        );

    \I__5561\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27079\
        );

    \I__5560\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27079\
        );

    \I__5559\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27079\
        );

    \I__5558\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27073\
        );

    \I__5557\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27073\
        );

    \I__5556\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27070\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__27105\,
            I => \N__27066\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__27102\,
            I => \N__27055\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__27097\,
            I => \N__27055\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__27094\,
            I => \N__27055\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__27089\,
            I => \N__27055\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__27086\,
            I => \N__27055\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__27079\,
            I => \N__27050\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__27078\,
            I => \N__27047\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__27073\,
            I => \N__27044\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__27070\,
            I => \N__27041\
        );

    \I__5545\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27038\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__27066\,
            I => \N__27035\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__27055\,
            I => \N__27032\
        );

    \I__5542\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27027\
        );

    \I__5541\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27027\
        );

    \I__5540\ : Span12Mux_s6_h
    port map (
            O => \N__27050\,
            I => \N__27024\
        );

    \I__5539\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27021\
        );

    \I__5538\ : Span4Mux_v
    port map (
            O => \N__27044\,
            I => \N__27014\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__27041\,
            I => \N__27014\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27014\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__27035\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__27032\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__27027\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5532\ : Odrv12
    port map (
            O => \N__27024\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__27021\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__27014\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5529\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26998\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26995\
        );

    \I__5527\ : Odrv12
    port map (
            O => \N__26995\,
            I => \POWERLED.N_145_N\
        );

    \I__5526\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26989\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__26989\,
            I => \POWERLED.un1_clk_100khz_51_and_i_a2_5_0\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__26986\,
            I => \POWERLED.un1_clk_100khz_51_and_i_a2_5_0_cascade_\
        );

    \I__5523\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26974\
        );

    \I__5522\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26974\
        );

    \I__5521\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26974\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__5519\ : Span4Mux_v
    port map (
            O => \N__26971\,
            I => \N__26966\
        );

    \I__5518\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26963\
        );

    \I__5517\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26960\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__26966\,
            I => \RSMRSTn_fast\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__26963\,
            I => \RSMRSTn_fast\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__26960\,
            I => \RSMRSTn_fast\
        );

    \I__5513\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__26950\,
            I => \POWERLED.func_state_RNIPUGOZ0Z_1\
        );

    \I__5511\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26943\
        );

    \I__5510\ : InMux
    port map (
            O => \N__26946\,
            I => \N__26939\
        );

    \I__5509\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26934\
        );

    \I__5508\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26934\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__26939\,
            I => \POWERLED.N_340\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__26934\,
            I => \POWERLED.N_340\
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__26929\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_\
        );

    \I__5504\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26923\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__26923\,
            I => \POWERLED.N_284\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26896\
        );

    \I__5501\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26896\
        );

    \I__5500\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26896\
        );

    \I__5499\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26896\
        );

    \I__5498\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26887\
        );

    \I__5497\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26887\
        );

    \I__5496\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26887\
        );

    \I__5495\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26887\
        );

    \I__5494\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26880\
        );

    \I__5493\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26880\
        );

    \I__5492\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26880\
        );

    \I__5491\ : InMux
    port map (
            O => \N__26909\,
            I => \N__26875\
        );

    \I__5490\ : InMux
    port map (
            O => \N__26908\,
            I => \N__26875\
        );

    \I__5489\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26868\
        );

    \I__5488\ : InMux
    port map (
            O => \N__26906\,
            I => \N__26868\
        );

    \I__5487\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26868\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__26896\,
            I => \N__26865\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__26887\,
            I => \N__26856\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__26880\,
            I => \N__26856\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__26875\,
            I => \N__26853\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26848\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__26865\,
            I => \N__26848\
        );

    \I__5480\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26839\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26839\
        );

    \I__5478\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26839\
        );

    \I__5477\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26839\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__26856\,
            I => \N__26836\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__26853\,
            I => \N__26833\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__26848\,
            I => \N__26828\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26828\
        );

    \I__5472\ : Span4Mux_h
    port map (
            O => \N__26836\,
            I => \N__26825\
        );

    \I__5471\ : Span4Mux_v
    port map (
            O => \N__26833\,
            I => \N__26820\
        );

    \I__5470\ : Span4Mux_v
    port map (
            O => \N__26828\,
            I => \N__26820\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__26825\,
            I => \POWERLED.func_state_RNIBQDB2Z0Z_0\
        );

    \I__5468\ : Odrv4
    port map (
            O => \N__26820\,
            I => \POWERLED.func_state_RNIBQDB2Z0Z_0\
        );

    \I__5467\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26809\
        );

    \I__5466\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26809\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__26809\,
            I => \N__26806\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__26806\,
            I => \POWERLED.N_340_N\
        );

    \I__5463\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26799\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__26802\,
            I => \N__26796\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26793\
        );

    \I__5460\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26790\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__26793\,
            I => \POWERLED.func_state_RNI_1Z0Z_0\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__26790\,
            I => \POWERLED.func_state_RNI_1Z0Z_0\
        );

    \I__5457\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26782\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__26782\,
            I => \POWERLED.un1_func_state25_6_0_o_N_294_N\
        );

    \I__5455\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26776\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26773\
        );

    \I__5453\ : Odrv12
    port map (
            O => \N__26773\,
            I => \POWERLED.func_state_1_m2_am_1_1\
        );

    \I__5452\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26760\
        );

    \I__5451\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26760\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__26768\,
            I => \N__26756\
        );

    \I__5449\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26752\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26749\
        );

    \I__5447\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26746\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26743\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__26759\,
            I => \N__26738\
        );

    \I__5444\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26733\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26733\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__26752\,
            I => \N__26728\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26728\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26725\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__26743\,
            I => \N__26722\
        );

    \I__5438\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26717\
        );

    \I__5437\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26717\
        );

    \I__5436\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26712\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__26733\,
            I => \N__26701\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__26728\,
            I => \N__26701\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__26725\,
            I => \N__26701\
        );

    \I__5432\ : Span4Mux_h
    port map (
            O => \N__26722\,
            I => \N__26701\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26701\
        );

    \I__5430\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26695\
        );

    \I__5429\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26695\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__26712\,
            I => \N__26686\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__26701\,
            I => \N__26683\
        );

    \I__5426\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26679\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__26695\,
            I => \N__26674\
        );

    \I__5424\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26667\
        );

    \I__5423\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26667\
        );

    \I__5422\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26667\
        );

    \I__5421\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26660\
        );

    \I__5420\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26660\
        );

    \I__5419\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26660\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__26686\,
            I => \N__26655\
        );

    \I__5417\ : Span4Mux_s3_h
    port map (
            O => \N__26683\,
            I => \N__26655\
        );

    \I__5416\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26652\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__26679\,
            I => \N__26649\
        );

    \I__5414\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26644\
        );

    \I__5413\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26644\
        );

    \I__5412\ : Sp12to4
    port map (
            O => \N__26674\,
            I => \N__26639\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__26667\,
            I => \N__26639\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__26660\,
            I => \POWERLED.func_N_5_mux_0\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__26655\,
            I => \POWERLED.func_N_5_mux_0\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__26652\,
            I => \POWERLED.func_N_5_mux_0\
        );

    \I__5407\ : Odrv12
    port map (
            O => \N__26649\,
            I => \POWERLED.func_N_5_mux_0\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__26644\,
            I => \POWERLED.func_N_5_mux_0\
        );

    \I__5405\ : Odrv12
    port map (
            O => \N__26639\,
            I => \POWERLED.func_N_5_mux_0\
        );

    \I__5404\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26620\
        );

    \I__5402\ : Odrv12
    port map (
            O => \N__26620\,
            I => \POWERLED.func_state_RNIBL3Q3Z0Z_1\
        );

    \I__5401\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26614\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__26614\,
            I => \N__26611\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__26608\,
            I => \POWERLED.func_state_1_m2s2_i_a2_0_0\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__26605\,
            I => \N__26596\
        );

    \I__5396\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26591\
        );

    \I__5395\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26588\
        );

    \I__5394\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26583\
        );

    \I__5393\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26583\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__26600\,
            I => \N__26580\
        );

    \I__5391\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26571\
        );

    \I__5390\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26566\
        );

    \I__5389\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26566\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26563\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26560\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26555\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__26583\,
            I => \N__26555\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26552\
        );

    \I__5383\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26549\
        );

    \I__5382\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26546\
        );

    \I__5381\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26540\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26540\
        );

    \I__5379\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26535\
        );

    \I__5378\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26535\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__26571\,
            I => \N__26532\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26566\,
            I => \N__26527\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__26563\,
            I => \N__26527\
        );

    \I__5374\ : Span4Mux_s3_h
    port map (
            O => \N__26560\,
            I => \N__26522\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__26555\,
            I => \N__26522\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__26552\,
            I => \N__26517\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26517\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__26546\,
            I => \N__26513\
        );

    \I__5369\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26510\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__26540\,
            I => \N__26505\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__26535\,
            I => \N__26505\
        );

    \I__5366\ : Span12Mux_s10_v
    port map (
            O => \N__26532\,
            I => \N__26502\
        );

    \I__5365\ : Span4Mux_v
    port map (
            O => \N__26527\,
            I => \N__26499\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__26522\,
            I => \N__26494\
        );

    \I__5363\ : Span4Mux_v
    port map (
            O => \N__26517\,
            I => \N__26494\
        );

    \I__5362\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26491\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__26513\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__26510\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5359\ : Odrv4
    port map (
            O => \N__26505\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5358\ : Odrv12
    port map (
            O => \N__26502\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__26499\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__26494\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__26491\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5354\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26471\
        );

    \I__5353\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26463\
        );

    \I__5352\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26463\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26471\,
            I => \N__26460\
        );

    \I__5350\ : InMux
    port map (
            O => \N__26470\,
            I => \N__26457\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26469\,
            I => \N__26451\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26451\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26448\
        );

    \I__5346\ : Span4Mux_v
    port map (
            O => \N__26460\,
            I => \N__26445\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__26457\,
            I => \N__26442\
        );

    \I__5344\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26439\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__26451\,
            I => \N__26432\
        );

    \I__5342\ : Span4Mux_v
    port map (
            O => \N__26448\,
            I => \N__26432\
        );

    \I__5341\ : Span4Mux_v
    port map (
            O => \N__26445\,
            I => \N__26432\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__26442\,
            I => \N__26427\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__26439\,
            I => \N__26427\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__26432\,
            I => \func_state_RNI_7_1\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__26427\,
            I => \func_state_RNI_7_1\
        );

    \I__5336\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26419\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__26419\,
            I => \N__26416\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__26416\,
            I => \N_7\
        );

    \I__5333\ : IoInMux
    port map (
            O => \N__26413\,
            I => \N__26408\
        );

    \I__5332\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26405\
        );

    \I__5331\ : CascadeMux
    port map (
            O => \N__26411\,
            I => \N__26401\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__26408\,
            I => \N__26398\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__26405\,
            I => \N__26394\
        );

    \I__5328\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26391\
        );

    \I__5327\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26388\
        );

    \I__5326\ : IoSpan4Mux
    port map (
            O => \N__26398\,
            I => \N__26383\
        );

    \I__5325\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26380\
        );

    \I__5324\ : Span4Mux_h
    port map (
            O => \N__26394\,
            I => \N__26373\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__26391\,
            I => \N__26373\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26373\
        );

    \I__5321\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26370\
        );

    \I__5320\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26367\
        );

    \I__5319\ : Span4Mux_s1_v
    port map (
            O => \N__26383\,
            I => \N__26362\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__26380\,
            I => \N__26362\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__26373\,
            I => \N__26359\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26356\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__26367\,
            I => \N__26348\
        );

    \I__5314\ : Span4Mux_h
    port map (
            O => \N__26362\,
            I => \N__26341\
        );

    \I__5313\ : Span4Mux_s3_h
    port map (
            O => \N__26359\,
            I => \N__26341\
        );

    \I__5312\ : Span4Mux_s1_v
    port map (
            O => \N__26356\,
            I => \N__26341\
        );

    \I__5311\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26338\
        );

    \I__5310\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26333\
        );

    \I__5309\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26333\
        );

    \I__5308\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26328\
        );

    \I__5307\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26328\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__26348\,
            I => \N__26325\
        );

    \I__5305\ : Sp12to4
    port map (
            O => \N__26341\,
            I => \N__26318\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__26338\,
            I => \N__26318\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__26333\,
            I => \N__26318\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26328\,
            I => rsmrstn
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__26325\,
            I => rsmrstn
        );

    \I__5300\ : Odrv12
    port map (
            O => \N__26318\,
            I => rsmrstn
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__26311\,
            I => \G_34_0_a4_0_2_cascade_\
        );

    \I__5298\ : CascadeMux
    port map (
            O => \N__26308\,
            I => \N__26305\
        );

    \I__5297\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26299\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26299\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__26299\,
            I => \POWERLED_un1_dutycycle_172_m3_0_0\
        );

    \I__5294\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26290\
        );

    \I__5293\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26290\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__26290\,
            I => \POWERLED.N_8_0\
        );

    \I__5291\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26282\
        );

    \I__5290\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26277\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26277\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__26282\,
            I => \N__26274\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__26277\,
            I => \N__26271\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__26274\,
            I => \N__26268\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__26271\,
            I => \POWERLED.un1_dutycycle_172_m1_ns_1\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__26268\,
            I => \POWERLED.un1_dutycycle_172_m1_ns_1\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__26263\,
            I => \N__26260\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26254\
        );

    \I__5281\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26254\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__5279\ : Span4Mux_v
    port map (
            O => \N__26251\,
            I => \N__26246\
        );

    \I__5278\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26243\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__26249\,
            I => \N__26240\
        );

    \I__5276\ : Sp12to4
    port map (
            O => \N__26246\,
            I => \N__26234\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__26243\,
            I => \N__26234\
        );

    \I__5274\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26231\
        );

    \I__5273\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26228\
        );

    \I__5272\ : Span12Mux_s5_h
    port map (
            O => \N__26234\,
            I => \N__26223\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__26231\,
            I => \N__26223\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__26228\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_3\
        );

    \I__5269\ : Odrv12
    port map (
            O => \N__26223\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_3\
        );

    \I__5268\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26215\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__26215\,
            I => \N_11\
        );

    \I__5266\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26206\
        );

    \I__5265\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26203\
        );

    \I__5264\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26200\
        );

    \I__5263\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26196\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__26206\,
            I => \N__26193\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26190\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__26200\,
            I => \N__26187\
        );

    \I__5259\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26184\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__26196\,
            I => \N__26181\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__26193\,
            I => \N__26178\
        );

    \I__5256\ : Span12Mux_s10_v
    port map (
            O => \N__26190\,
            I => \N__26175\
        );

    \I__5255\ : Odrv12
    port map (
            O => \N__26187\,
            I => \POWERLED.N_319_0\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__26184\,
            I => \POWERLED.N_319_0\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__26181\,
            I => \POWERLED.N_319_0\
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__26178\,
            I => \POWERLED.N_319_0\
        );

    \I__5251\ : Odrv12
    port map (
            O => \N__26175\,
            I => \POWERLED.N_319_0\
        );

    \I__5250\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26158\
        );

    \I__5249\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26158\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__26157\,
            I => \N__26148\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__26156\,
            I => \N__26144\
        );

    \I__5245\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26141\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__26152\,
            I => \N__26138\
        );

    \I__5243\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26135\
        );

    \I__5242\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26130\
        );

    \I__5241\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26130\
        );

    \I__5240\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26127\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__26141\,
            I => \N__26124\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__26138\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__26135\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__26130\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__26127\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5234\ : Odrv12
    port map (
            O => \N__26124\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5233\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26110\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__26110\,
            I => \POWERLED.N_297\
        );

    \I__5231\ : InMux
    port map (
            O => \N__26107\,
            I => \N__26104\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__26104\,
            I => \N__26101\
        );

    \I__5229\ : Odrv4
    port map (
            O => \N__26101\,
            I => \POWERLED.un1_func_state25_6_0_a2_1\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__26098\,
            I => \POWERLED.un1_func_state25_6_0_o_N_296_N_cascade_\
        );

    \I__5227\ : CascadeMux
    port map (
            O => \N__26095\,
            I => \POWERLED.un1_func_state25_6_0_1_cascade_\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__26092\,
            I => \N__26089\
        );

    \I__5225\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26086\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__26086\,
            I => \N__26083\
        );

    \I__5223\ : Span4Mux_h
    port map (
            O => \N__26083\,
            I => \N__26080\
        );

    \I__5222\ : Span4Mux_v
    port map (
            O => \N__26080\,
            I => \N__26077\
        );

    \I__5221\ : Odrv4
    port map (
            O => \N__26077\,
            I => \POWERLED.un1_func_state25_6_0_2\
        );

    \I__5220\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26071\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26065\
        );

    \I__5218\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26060\
        );

    \I__5217\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26060\
        );

    \I__5216\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26057\
        );

    \I__5215\ : Odrv12
    port map (
            O => \N__26065\,
            I => \RSMRSTn_rep1\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__26060\,
            I => \RSMRSTn_rep1\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__26057\,
            I => \RSMRSTn_rep1\
        );

    \I__5212\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26043\
        );

    \I__5211\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26038\
        );

    \I__5210\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26038\
        );

    \I__5209\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26031\
        );

    \I__5208\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26031\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__26043\,
            I => \N__26026\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__26038\,
            I => \N__26026\
        );

    \I__5205\ : InMux
    port map (
            O => \N__26037\,
            I => \N__26021\
        );

    \I__5204\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26021\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__26031\,
            I => \N__26018\
        );

    \I__5202\ : Span4Mux_v
    port map (
            O => \N__26026\,
            I => \N__26013\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26013\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__26018\,
            I => \N__26010\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__26013\,
            I => \N__26007\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__26010\,
            I => \POWERLED.N_4_0_3\
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__26007\,
            I => \POWERLED.N_4_0_3\
        );

    \I__5196\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25998\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__26001\,
            I => \N__25993\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__25998\,
            I => \N__25990\
        );

    \I__5193\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25987\
        );

    \I__5192\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25984\
        );

    \I__5191\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25981\
        );

    \I__5190\ : Span4Mux_v
    port map (
            O => \N__25990\,
            I => \N__25978\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25975\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25970\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__25981\,
            I => \N__25970\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__25978\,
            I => \POWERLED.func_state_RNIOGRSZ0Z_0\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__25975\,
            I => \POWERLED.func_state_RNIOGRSZ0Z_0\
        );

    \I__5184\ : Odrv4
    port map (
            O => \N__25970\,
            I => \POWERLED.func_state_RNIOGRSZ0Z_0\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__25963\,
            I => \N__25959\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__25962\,
            I => \N__25956\
        );

    \I__5181\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25953\
        );

    \I__5180\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25950\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__25953\,
            I => \N__25947\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25942\
        );

    \I__5177\ : Span4Mux_h
    port map (
            O => \N__25947\,
            I => \N__25942\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__25942\,
            I => \POWERLED.func_state_1_ss0_i_0_o2_1\
        );

    \I__5175\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25935\
        );

    \I__5174\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25932\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25927\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__25932\,
            I => \N__25927\
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__25927\,
            I => \POWERLED.N_76\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__25924\,
            I => \POWERLED.func_state_RNI91IA4Z0Z_1_cascade_\
        );

    \I__5169\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25918\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__25918\,
            I => \POWERLED.func_state_1_m2_1\
        );

    \I__5167\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25909\
        );

    \I__5166\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25909\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__25909\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \POWERLED.func_state_1_m2_1_cascade_\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__25903\,
            I => \N__25900\
        );

    \I__5162\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25897\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__25897\,
            I => \N__25891\
        );

    \I__5160\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25888\
        );

    \I__5159\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25883\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25883\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__25891\,
            I => \N__25876\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__25888\,
            I => \N__25876\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__25883\,
            I => \N__25876\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__25876\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__25873\,
            I => \N__25869\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__25872\,
            I => \N__25866\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25857\
        );

    \I__5150\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25854\
        );

    \I__5149\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25849\
        );

    \I__5148\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25849\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25843\
        );

    \I__5146\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25843\
        );

    \I__5145\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25840\
        );

    \I__5144\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25837\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__25857\,
            I => \N__25830\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25830\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__25849\,
            I => \N__25830\
        );

    \I__5140\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25827\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__25843\,
            I => \N__25824\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__25840\,
            I => \N__25821\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__25837\,
            I => \N__25818\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__25830\,
            I => \N__25814\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__25827\,
            I => \N__25809\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__25824\,
            I => \N__25809\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__25821\,
            I => \N__25804\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__25818\,
            I => \N__25804\
        );

    \I__5131\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25801\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__25814\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__25809\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__25804\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__25801\,
            I => \POWERLED.un1_N_3_mux_0\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__25792\,
            I => \N_4_1_cascade_\
        );

    \I__5125\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25786\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__25786\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25780\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__25780\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__5121\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25774\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__25774\,
            I => \N__25771\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__25768\,
            I => \N__25765\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__25762\,
            I => \POWERLED.count_off_0_5\
        );

    \I__5115\ : InMux
    port map (
            O => \N__25759\,
            I => \N__25756\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__25756\,
            I => \N__25752\
        );

    \I__5113\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25749\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__25752\,
            I => \N__25746\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__25749\,
            I => \N__25743\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__25746\,
            I => \N__25740\
        );

    \I__5109\ : Odrv12
    port map (
            O => \N__25743\,
            I => \POWERLED.count_off_1_5\
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__25740\,
            I => \POWERLED.count_off_1_5\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25731\
        );

    \I__5106\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25728\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25725\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__25728\,
            I => \N__25722\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__25725\,
            I => \N__25719\
        );

    \I__5102\ : Sp12to4
    port map (
            O => \N__25722\,
            I => \N__25716\
        );

    \I__5101\ : Span4Mux_v
    port map (
            O => \N__25719\,
            I => \N__25713\
        );

    \I__5100\ : Odrv12
    port map (
            O => \N__25716\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__25713\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__5098\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__25705\,
            I => \N__25702\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__5095\ : Span4Mux_h
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__5094\ : Span4Mux_v
    port map (
            O => \N__25696\,
            I => \N__25693\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__25693\,
            I => \POWERLED.count_off_0_6\
        );

    \I__5092\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25686\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25683\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25680\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__25683\,
            I => \N__25677\
        );

    \I__5088\ : Span12Mux_s6_h
    port map (
            O => \N__25680\,
            I => \N__25674\
        );

    \I__5087\ : Odrv12
    port map (
            O => \N__25677\,
            I => \POWERLED.count_off_1_6\
        );

    \I__5086\ : Odrv12
    port map (
            O => \N__25674\,
            I => \POWERLED.count_off_1_6\
        );

    \I__5085\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25665\
        );

    \I__5084\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25662\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25659\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__25662\,
            I => \N__25656\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__25659\,
            I => \N__25653\
        );

    \I__5080\ : Span12Mux_s8_v
    port map (
            O => \N__25656\,
            I => \N__25650\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__25653\,
            I => \N__25647\
        );

    \I__5078\ : Odrv12
    port map (
            O => \N__25650\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__25647\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__25639\,
            I => \N__25636\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__25636\,
            I => \N__25633\
        );

    \I__5073\ : Span4Mux_h
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__5072\ : Span4Mux_v
    port map (
            O => \N__25630\,
            I => \N__25627\
        );

    \I__5071\ : Odrv4
    port map (
            O => \N__25627\,
            I => \POWERLED.count_off_0_2\
        );

    \I__5070\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25617\
        );

    \I__5068\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25614\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__25617\,
            I => \N__25611\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__25614\,
            I => \N__25608\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__25611\,
            I => \N__25605\
        );

    \I__5064\ : Span4Mux_h
    port map (
            O => \N__25608\,
            I => \N__25602\
        );

    \I__5063\ : Odrv4
    port map (
            O => \N__25605\,
            I => \POWERLED.count_off_1_2\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__25602\,
            I => \POWERLED.count_off_1_2\
        );

    \I__5061\ : CEMux
    port map (
            O => \N__25597\,
            I => \N__25593\
        );

    \I__5060\ : CEMux
    port map (
            O => \N__25596\,
            I => \N__25587\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__25593\,
            I => \N__25584\
        );

    \I__5058\ : CEMux
    port map (
            O => \N__25592\,
            I => \N__25580\
        );

    \I__5057\ : CascadeMux
    port map (
            O => \N__25591\,
            I => \N__25575\
        );

    \I__5056\ : CEMux
    port map (
            O => \N__25590\,
            I => \N__25571\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__25587\,
            I => \N__25565\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__25584\,
            I => \N__25562\
        );

    \I__5053\ : CEMux
    port map (
            O => \N__25583\,
            I => \N__25559\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__25580\,
            I => \N__25554\
        );

    \I__5051\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25541\
        );

    \I__5050\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25541\
        );

    \I__5049\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25541\
        );

    \I__5048\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25541\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__25571\,
            I => \N__25538\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25531\
        );

    \I__5045\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25531\
        );

    \I__5044\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25531\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__25565\,
            I => \N__25528\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__25562\,
            I => \N__25523\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25523\
        );

    \I__5040\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25518\
        );

    \I__5039\ : CEMux
    port map (
            O => \N__25557\,
            I => \N__25518\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__25554\,
            I => \N__25514\
        );

    \I__5037\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25505\
        );

    \I__5036\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25505\
        );

    \I__5035\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25505\
        );

    \I__5034\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25505\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25502\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__25538\,
            I => \N__25497\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__25531\,
            I => \N__25497\
        );

    \I__5030\ : Span4Mux_h
    port map (
            O => \N__25528\,
            I => \N__25492\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__25523\,
            I => \N__25489\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__25518\,
            I => \N__25486\
        );

    \I__5027\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25483\
        );

    \I__5026\ : Span4Mux_s3_h
    port map (
            O => \N__25514\,
            I => \N__25474\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__25505\,
            I => \N__25474\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__25502\,
            I => \N__25474\
        );

    \I__5023\ : Span4Mux_v
    port map (
            O => \N__25497\,
            I => \N__25474\
        );

    \I__5022\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25469\
        );

    \I__5021\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25469\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__25492\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__25489\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0\
        );

    \I__5018\ : Odrv4
    port map (
            O => \N__25486\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__25483\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__25474\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__25469\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0\
        );

    \I__5014\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25452\
        );

    \I__5013\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25449\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__25452\,
            I => \N__25446\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25441\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__25446\,
            I => \N__25441\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__25441\,
            I => \N__25438\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__25438\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__5007\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__25432\,
            I => \N__25428\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__25431\,
            I => \N__25423\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__25428\,
            I => \N__25419\
        );

    \I__5003\ : InMux
    port map (
            O => \N__25427\,
            I => \N__25416\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25413\
        );

    \I__5001\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25408\
        );

    \I__5000\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25408\
        );

    \I__4999\ : Sp12to4
    port map (
            O => \N__25419\,
            I => \N__25400\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__25416\,
            I => \N__25400\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25413\,
            I => \N__25395\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25395\
        );

    \I__4995\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25390\
        );

    \I__4994\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25390\
        );

    \I__4993\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25387\
        );

    \I__4992\ : Odrv12
    port map (
            O => \N__25400\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__25395\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__25390\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__25387\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4988\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25372\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__25377\,
            I => \N__25367\
        );

    \I__4986\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25362\
        );

    \I__4985\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25359\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__25372\,
            I => \N__25356\
        );

    \I__4983\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25353\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__25370\,
            I => \N__25350\
        );

    \I__4981\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25345\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25345\
        );

    \I__4979\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25342\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__25362\,
            I => \N__25338\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__25359\,
            I => \N__25331\
        );

    \I__4976\ : Span4Mux_h
    port map (
            O => \N__25356\,
            I => \N__25331\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__25353\,
            I => \N__25331\
        );

    \I__4974\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25328\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25323\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25323\
        );

    \I__4971\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25320\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__25338\,
            I => \N__25313\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__25331\,
            I => \N__25313\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__25328\,
            I => \N__25313\
        );

    \I__4967\ : Odrv12
    port map (
            O => \N__25323\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__25320\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__25313\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4964\ : InMux
    port map (
            O => \N__25306\,
            I => \N__25302\
        );

    \I__4963\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25299\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__25302\,
            I => \N__25296\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__25299\,
            I => \N__25293\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__25296\,
            I => \N__25290\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__25293\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_13\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__25290\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_13\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25282\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__25282\,
            I => \N__25279\
        );

    \I__4955\ : Span4Mux_h
    port map (
            O => \N__25279\,
            I => \N__25276\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__25276\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_15\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__25273\,
            I => \N__25263\
        );

    \I__4952\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25252\
        );

    \I__4951\ : InMux
    port map (
            O => \N__25271\,
            I => \N__25252\
        );

    \I__4950\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25252\
        );

    \I__4949\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25252\
        );

    \I__4948\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25252\
        );

    \I__4947\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25247\
        );

    \I__4946\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25247\
        );

    \I__4945\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25244\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__25252\,
            I => \N__25241\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__25247\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__25244\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4941\ : Odrv12
    port map (
            O => \N__25241\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__25234\,
            I => \N__25229\
        );

    \I__4939\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25222\
        );

    \I__4938\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25222\
        );

    \I__4937\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25222\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__25222\,
            I => \N__25217\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__25221\,
            I => \N__25214\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__25220\,
            I => \N__25211\
        );

    \I__4933\ : Span4Mux_s3_v
    port map (
            O => \N__25217\,
            I => \N__25204\
        );

    \I__4932\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25191\
        );

    \I__4931\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25191\
        );

    \I__4930\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25191\
        );

    \I__4929\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25191\
        );

    \I__4928\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25191\
        );

    \I__4927\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25191\
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__25204\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__25191\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__4924\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__25183\,
            I => \POWERLED.N_301\
        );

    \I__4922\ : SRMux
    port map (
            O => \N__25180\,
            I => \N__25177\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25174\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__25174\,
            I => \N__25169\
        );

    \I__4919\ : SRMux
    port map (
            O => \N__25173\,
            I => \N__25166\
        );

    \I__4918\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25162\
        );

    \I__4917\ : Span4Mux_s2_v
    port map (
            O => \N__25169\,
            I => \N__25157\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25157\
        );

    \I__4915\ : SRMux
    port map (
            O => \N__25165\,
            I => \N__25154\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__25162\,
            I => \N__25151\
        );

    \I__4913\ : Sp12to4
    port map (
            O => \N__25157\,
            I => \N__25148\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__25154\,
            I => \N__25145\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__25151\,
            I => \N__25142\
        );

    \I__4910\ : Odrv12
    port map (
            O => \N__25148\,
            I => \G_11\
        );

    \I__4909\ : Odrv12
    port map (
            O => \N__25145\,
            I => \G_11\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__25142\,
            I => \G_11\
        );

    \I__4907\ : CEMux
    port map (
            O => \N__25135\,
            I => \N__25132\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__25126\,
            I => \RSMRST_PWRGD.N_29_2\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__25123\,
            I => \N__25114\
        );

    \I__4902\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25111\
        );

    \I__4901\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25107\
        );

    \I__4900\ : CascadeMux
    port map (
            O => \N__25120\,
            I => \N__25103\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__25119\,
            I => \N__25100\
        );

    \I__4898\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25093\
        );

    \I__4897\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25090\
        );

    \I__4896\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25087\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__25111\,
            I => \N__25084\
        );

    \I__4894\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25081\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__25107\,
            I => \N__25078\
        );

    \I__4892\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25075\
        );

    \I__4891\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25062\
        );

    \I__4890\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25062\
        );

    \I__4889\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25062\
        );

    \I__4888\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25062\
        );

    \I__4887\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25062\
        );

    \I__4886\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25062\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__25093\,
            I => \N__25051\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__25090\,
            I => \N__25051\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__25087\,
            I => \N__25051\
        );

    \I__4882\ : Span4Mux_s3_v
    port map (
            O => \N__25084\,
            I => \N__25051\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25051\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__25078\,
            I => \N__25048\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__25075\,
            I => \N__25043\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__25062\,
            I => \N__25043\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__25051\,
            I => \N__25040\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__25048\,
            I => \N__25035\
        );

    \I__4875\ : Span4Mux_s2_v
    port map (
            O => \N__25043\,
            I => \N__25035\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__25040\,
            I => \N__25032\
        );

    \I__4873\ : Odrv4
    port map (
            O => \N__25035\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__25032\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__25027\,
            I => \N__25023\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__25026\,
            I => \N__25020\
        );

    \I__4869\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25013\
        );

    \I__4868\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25013\
        );

    \I__4867\ : InMux
    port map (
            O => \N__25019\,
            I => \N__25010\
        );

    \I__4866\ : InMux
    port map (
            O => \N__25018\,
            I => \N__25007\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__25013\,
            I => \N__25004\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__25010\,
            I => \N__25001\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__25007\,
            I => \N__24998\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__25004\,
            I => \N__24995\
        );

    \I__4861\ : Span4Mux_h
    port map (
            O => \N__25001\,
            I => \N__24992\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__24998\,
            I => \N__24988\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__24995\,
            I => \N__24985\
        );

    \I__4858\ : Span4Mux_s2_h
    port map (
            O => \N__24992\,
            I => \N__24982\
        );

    \I__4857\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24979\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__24988\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__24985\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__24982\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__24979\,
            I => \POWERLED.dutycycle_N_3_mux_0\
        );

    \I__4852\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24967\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__24967\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__4850\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__24961\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__24958\,
            I => \VPP_VDDQ.count_2_1_9_cascade_\
        );

    \I__4847\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__24952\,
            I => \VPP_VDDQ.count_2_0_10\
        );

    \I__4845\ : IoInMux
    port map (
            O => \N__24949\,
            I => \N__24946\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__4843\ : IoSpan4Mux
    port map (
            O => \N__24943\,
            I => \N__24939\
        );

    \I__4842\ : IoInMux
    port map (
            O => \N__24942\,
            I => \N__24936\
        );

    \I__4841\ : IoSpan4Mux
    port map (
            O => \N__24939\,
            I => \N__24930\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__24936\,
            I => \N__24930\
        );

    \I__4839\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24927\
        );

    \I__4838\ : IoSpan4Mux
    port map (
            O => \N__24930\,
            I => \N__24924\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24921\
        );

    \I__4836\ : Span4Mux_s3_h
    port map (
            O => \N__24924\,
            I => \N__24918\
        );

    \I__4835\ : Span4Mux_h
    port map (
            O => \N__24921\,
            I => \N__24915\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__24918\,
            I => \N__24912\
        );

    \I__4833\ : Span4Mux_v
    port map (
            O => \N__24915\,
            I => \N__24909\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__24912\,
            I => \N__24904\
        );

    \I__4831\ : Span4Mux_v
    port map (
            O => \N__24909\,
            I => \N__24904\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__24904\,
            I => v33a_ok
        );

    \I__4829\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24898\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__24898\,
            I => \N__24895\
        );

    \I__4827\ : Span4Mux_v
    port map (
            O => \N__24895\,
            I => \N__24892\
        );

    \I__4826\ : Sp12to4
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__4825\ : Odrv12
    port map (
            O => \N__24889\,
            I => v5a_ok
        );

    \I__4824\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__24883\,
            I => \N__24879\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__24882\,
            I => \N__24876\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__24879\,
            I => \N__24873\
        );

    \I__4820\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24870\
        );

    \I__4819\ : Span4Mux_h
    port map (
            O => \N__24873\,
            I => \N__24867\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__24870\,
            I => \N__24864\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__24867\,
            I => slp_susn
        );

    \I__4816\ : Odrv12
    port map (
            O => \N__24864\,
            I => slp_susn
        );

    \I__4815\ : IoInMux
    port map (
            O => \N__24859\,
            I => \N__24856\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__24856\,
            I => \N__24852\
        );

    \I__4813\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24849\
        );

    \I__4812\ : Span4Mux_s2_h
    port map (
            O => \N__24852\,
            I => \N__24846\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24843\
        );

    \I__4810\ : Sp12to4
    port map (
            O => \N__24846\,
            I => \N__24838\
        );

    \I__4809\ : Sp12to4
    port map (
            O => \N__24843\,
            I => \N__24838\
        );

    \I__4808\ : Span12Mux_s11_v
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__4807\ : Odrv12
    port map (
            O => \N__24835\,
            I => v1p8a_ok
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__24832\,
            I => \rsmrst_pwrgd_signal_cascade_\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__24829\,
            I => \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\
        );

    \I__4804\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24822\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__24825\,
            I => \N__24819\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__24822\,
            I => \N__24815\
        );

    \I__4801\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24810\
        );

    \I__4800\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24810\
        );

    \I__4799\ : Odrv12
    port map (
            O => \N__24815\,
            I => \N_382\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__24810\,
            I => \N_382\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__24805\,
            I => \N__24801\
        );

    \I__4796\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24798\
        );

    \I__4795\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24795\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__24798\,
            I => \N__24792\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24789\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__24792\,
            I => \N__24784\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__24789\,
            I => \N__24784\
        );

    \I__4790\ : Odrv4
    port map (
            O => \N__24784\,
            I => \RSMRST_PWRGD.N_254_i\
        );

    \I__4789\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24777\
        );

    \I__4788\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24774\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__24777\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__24774\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__4785\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24765\
        );

    \I__4784\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24762\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__24765\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__24762\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__24757\,
            I => \N__24754\
        );

    \I__4780\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24751\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__24751\,
            I => \N__24748\
        );

    \I__4778\ : Span4Mux_h
    port map (
            O => \N__24748\,
            I => \N__24745\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__24745\,
            I => \RSMRST_PWRGD.m4_0_a2_0\
        );

    \I__4776\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24738\
        );

    \I__4775\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24735\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__24738\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__24735\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24727\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__24727\,
            I => \RSMRST_PWRGD.m4_0_a2_12\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__24724\,
            I => \VPP_VDDQ.count_2_1_10_cascade_\
        );

    \I__4769\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24715\
        );

    \I__4768\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24715\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24712\
        );

    \I__4766\ : Span4Mux_h
    port map (
            O => \N__24712\,
            I => \N__24707\
        );

    \I__4765\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24704\
        );

    \I__4764\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24701\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__24707\,
            I => \PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__24704\,
            I => \PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__24701\,
            I => \PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0\
        );

    \I__4760\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__24691\,
            I => \PCH_PWRGD.curr_state_0_0\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__24688\,
            I => \PCH_PWRGD.m4_0_cascade_\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__24685\,
            I => \VPP_VDDQ.count_2_1_8_cascade_\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__24682\,
            I => \PCH_PWRGD.countZ0Z_0_cascade_\
        );

    \I__4755\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24673\
        );

    \I__4754\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24673\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__24673\,
            I => \PCH_PWRGD.N_2173_i\
        );

    \I__4752\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24666\
        );

    \I__4751\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24663\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__24666\,
            I => \PCH_PWRGD.count_1_i_a2_11_0\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__24663\,
            I => \PCH_PWRGD.count_1_i_a2_11_0\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__24658\,
            I => \PCH_PWRGD.N_2173_i_cascade_\
        );

    \I__4747\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24651\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24648\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__24651\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__24648\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__4743\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24639\
        );

    \I__4742\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24636\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__24639\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__24636\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__4739\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24627\
        );

    \I__4738\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24624\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__24627\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__24624\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__24619\,
            I => \RSMRST_PWRGD.m4_0_a2_11_cascade_\
        );

    \I__4734\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24612\
        );

    \I__4733\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24609\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__24612\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__24609\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24600\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24597\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__24600\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24597\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__24592\,
            I => \N__24588\
        );

    \I__4725\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24585\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24582\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__24585\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__24582\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__4721\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24573\
        );

    \I__4720\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24570\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__24573\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__24570\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__4717\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__24562\,
            I => \RSMRST_PWRGD.m4_0_a2_10\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24555\
        );

    \I__4714\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24552\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__24555\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__24552\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__4711\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24543\
        );

    \I__4710\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24540\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__24543\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__24540\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__24535\,
            I => \N__24531\
        );

    \I__4706\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24528\
        );

    \I__4705\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24525\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__24528\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__24525\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__4702\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24516\
        );

    \I__4701\ : InMux
    port map (
            O => \N__24519\,
            I => \N__24513\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__24516\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__24513\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24505\,
            I => \RSMRST_PWRGD.m4_0_a2_9\
        );

    \I__4696\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24499\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__24499\,
            I => \N__24496\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__24496\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__4693\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24487\
        );

    \I__4692\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24487\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__24487\,
            I => \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\
        );

    \I__4690\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__24481\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__4688\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24472\
        );

    \I__4687\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24472\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__24472\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__24469\,
            I => \PCH_PWRGD.countZ0Z_6_cascade_\
        );

    \I__4684\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24461\
        );

    \I__4683\ : InMux
    port map (
            O => \N__24465\,
            I => \N__24456\
        );

    \I__4682\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24456\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__24461\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__24456\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__4679\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24448\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__24448\,
            I => \N__24445\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__24445\,
            I => \PCH_PWRGD.count_1_i_a2_1_0\
        );

    \I__4676\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__24439\,
            I => \N__24435\
        );

    \I__4674\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24432\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__24435\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__24432\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__24427\,
            I => \PCH_PWRGD.count_1_i_a2_0_0_cascade_\
        );

    \I__4670\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__24421\,
            I => \N__24418\
        );

    \I__4668\ : Span4Mux_v
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__24415\,
            I => \PCH_PWRGD.count_1_i_a2_2_0\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__24412\,
            I => \PCH_PWRGD.count_1_i_a2_11_0_cascade_\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__24409\,
            I => \PCH_PWRGD.count_rst_3_cascade_\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__24406\,
            I => \N_253_cascade_\
        );

    \I__4663\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__24400\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__4661\ : InMux
    port map (
            O => \N__24397\,
            I => \N__24394\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__24394\,
            I => \PCH_PWRGD.count_RNIM6A821Z0Z_1\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__24391\,
            I => \PCH_PWRGD.countZ0Z_3_cascade_\
        );

    \I__4658\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24382\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24382\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__24382\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__4655\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__24376\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__24373\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__24370\,
            I => \PCH_PWRGD.countZ0Z_8_cascade_\
        );

    \I__4651\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24361\
        );

    \I__4650\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24361\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__24361\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__4648\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__24355\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__4646\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24349\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__24349\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24343\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__24343\,
            I => \N__24339\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24336\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__24339\,
            I => \POWERLED.dutycycle_RNIZ0Z_6\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__24336\,
            I => \POWERLED.dutycycle_RNIZ0Z_6\
        );

    \I__4639\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24327\
        );

    \I__4638\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24324\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24327\,
            I => \N__24319\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__24324\,
            I => \N__24319\
        );

    \I__4635\ : Span12Mux_s10_v
    port map (
            O => \N__24319\,
            I => \N__24316\
        );

    \I__4634\ : Odrv12
    port map (
            O => \N__24316\,
            I => \POWERLED.un1_dutycycle_172_m3s4_1\
        );

    \I__4633\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24307\
        );

    \I__4632\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24307\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__24307\,
            I => \N__24302\
        );

    \I__4630\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24297\
        );

    \I__4629\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24297\
        );

    \I__4628\ : Odrv12
    port map (
            O => \N__24302\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_6\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__24297\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_6\
        );

    \I__4626\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24289\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__24289\,
            I => \POWERLED.N_239\
        );

    \I__4624\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24279\
        );

    \I__4622\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24276\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__24279\,
            I => \N__24273\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24270\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__24273\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__4618\ : Odrv12
    port map (
            O => \N__24270\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__24265\,
            I => \N__24262\
        );

    \I__4616\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24256\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__24256\,
            I => \POWERLED.N_271\
        );

    \I__4613\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24250\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__4611\ : Span4Mux_v
    port map (
            O => \N__24247\,
            I => \N__24243\
        );

    \I__4610\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24240\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__24243\,
            I => \POWERLED.N_366\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__24240\,
            I => \POWERLED.N_366\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \N__24230\
        );

    \I__4606\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24221\
        );

    \I__4605\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24221\
        );

    \I__4604\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24221\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__24229\,
            I => \N__24218\
        );

    \I__4602\ : InMux
    port map (
            O => \N__24228\,
            I => \N__24214\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__24221\,
            I => \N__24211\
        );

    \I__4600\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24208\
        );

    \I__4599\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24205\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24202\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__24211\,
            I => \N__24197\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__24208\,
            I => \N__24197\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__24205\,
            I => \POWERLED.N_331\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__24202\,
            I => \POWERLED.N_331\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__24197\,
            I => \POWERLED.N_331\
        );

    \I__4592\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24187\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__24187\,
            I => \POWERLED.N_272\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__24184\,
            I => \N__24181\
        );

    \I__4589\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24178\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__24178\,
            I => \N__24175\
        );

    \I__4587\ : Odrv12
    port map (
            O => \N__24175\,
            I => \POWERLED.dutycycle_N_3_mux_0_0\
        );

    \I__4586\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24169\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24166\
        );

    \I__4584\ : Odrv12
    port map (
            O => \N__24166\,
            I => \PCH_PWRGD.count_rst_10\
        );

    \I__4583\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24160\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__24160\,
            I => \N__24156\
        );

    \I__4581\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24153\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__24156\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__24153\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__4578\ : CascadeMux
    port map (
            O => \N__24148\,
            I => \PCH_PWRGD.count_rst_11_cascade_\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__24145\,
            I => \N__24142\
        );

    \I__4576\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24135\
        );

    \I__4575\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24135\
        );

    \I__4574\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24132\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__24135\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__24132\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__24127\,
            I => \POWERLED.count_off_1_sqmuxa_cascade_\
        );

    \I__4570\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24121\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__24121\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_6\
        );

    \I__4568\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24115\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24111\
        );

    \I__4566\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24108\
        );

    \I__4565\ : Span4Mux_h
    port map (
            O => \N__24111\,
            I => \N__24105\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24102\
        );

    \I__4563\ : Span4Mux_h
    port map (
            O => \N__24105\,
            I => \N__24099\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__24102\,
            I => \N__24096\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__24099\,
            I => \N__24093\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__24096\,
            I => \POWERLED.N_325\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__24093\,
            I => \POWERLED.N_325\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__24088\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_6_cascade_\
        );

    \I__4557\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24079\
        );

    \I__4556\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24074\
        );

    \I__4555\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24074\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__24082\,
            I => \N__24071\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__24079\,
            I => \N__24066\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24066\
        );

    \I__4551\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24063\
        );

    \I__4550\ : Span4Mux_v
    port map (
            O => \N__24066\,
            I => \N__24060\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24057\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__24060\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__24057\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__4546\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24048\
        );

    \I__4545\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24045\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__24048\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_0\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__24045\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_0\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__24040\,
            I => \N__24037\
        );

    \I__4541\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24033\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24030\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__24033\,
            I => \N__24027\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24024\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__24027\,
            I => \POWERLED.dutycycle_RNINH5P1Z0Z_2\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__24024\,
            I => \POWERLED.dutycycle_RNINH5P1Z0Z_2\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__24019\,
            I => \N__24015\
        );

    \I__4534\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24010\
        );

    \I__4533\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24010\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24010\,
            I => \N__24006\
        );

    \I__4531\ : InMux
    port map (
            O => \N__24009\,
            I => \N__24003\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__24006\,
            I => \POWERLED.dutycycle_RNI4G9K2Z0Z_5\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__24003\,
            I => \POWERLED.dutycycle_RNI4G9K2Z0Z_5\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__23998\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__23995\,
            I => \POWERLED.dutycycle_RNO_2Z0Z_5_cascade_\
        );

    \I__4526\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23989\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23986\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__23986\,
            I => \POWERLED.N_240\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__23983\,
            I => \N__23979\
        );

    \I__4522\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23976\
        );

    \I__4521\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23973\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__23976\,
            I => \N__23968\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N__23968\
        );

    \I__4518\ : Span4Mux_h
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__23965\,
            I => \N__23962\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__23962\,
            I => \POWERLED.dutycycle_eena_13\
        );

    \I__4515\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23956\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23956\,
            I => \N__23953\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__23950\,
            I => \POWERLED.un2_count_clk_17_0_0\
        );

    \I__4511\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23944\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__23944\,
            I => \POWERLED.g3\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__23941\,
            I => \POWERLED.un1_dutycycle_172_m3_1_0_cascade_\
        );

    \I__4508\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23935\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__23935\,
            I => \POWERLED.dutycycle_RNO_3Z0Z_5\
        );

    \I__4506\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23927\
        );

    \I__4505\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23922\
        );

    \I__4504\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23922\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__23927\,
            I => \POWERLED.dutycycle_1_0_5\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__23922\,
            I => \POWERLED.dutycycle_1_0_5\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__23917\,
            I => \N__23914\
        );

    \I__4500\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23911\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__23911\,
            I => \POWERLED.dutycycle_fb_15_1_1\
        );

    \I__4498\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23905\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23902\
        );

    \I__4496\ : Span4Mux_v
    port map (
            O => \N__23902\,
            I => \N__23899\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__23899\,
            I => \POWERLED.g2_0\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23893\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__4492\ : Odrv12
    port map (
            O => \N__23890\,
            I => \POWERLED.N_398_0\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__23884\,
            I => \POWERLED.g0_1_0\
        );

    \I__4489\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23876\
        );

    \I__4488\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23870\
        );

    \I__4487\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23870\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23867\
        );

    \I__4485\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23864\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__23870\,
            I => \N__23859\
        );

    \I__4483\ : Span4Mux_v
    port map (
            O => \N__23867\,
            I => \N__23859\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23856\
        );

    \I__4481\ : Span4Mux_v
    port map (
            O => \N__23859\,
            I => \N__23851\
        );

    \I__4480\ : Span4Mux_v
    port map (
            O => \N__23856\,
            I => \N__23851\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__23851\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_10\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23845\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__23839\,
            I => \POWERLED.func_state_1_m2s2_i_a3_0\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__23836\,
            I => \N__23833\
        );

    \I__4473\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23823\
        );

    \I__4471\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23820\
        );

    \I__4470\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23813\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23813\
        );

    \I__4468\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23813\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__23823\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__23820\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__23813\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4464\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__23803\,
            I => \N__23800\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__23800\,
            I => \POWERLED.dutycycle_fb_14_a4_1\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__23797\,
            I => \N__23793\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__23796\,
            I => \N__23787\
        );

    \I__4459\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23783\
        );

    \I__4458\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23778\
        );

    \I__4457\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23778\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__23790\,
            I => \N__23775\
        );

    \I__4455\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23770\
        );

    \I__4454\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23770\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23765\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__23778\,
            I => \N__23765\
        );

    \I__4451\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23762\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__23770\,
            I => \N__23752\
        );

    \I__4449\ : Span4Mux_v
    port map (
            O => \N__23765\,
            I => \N__23752\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__23762\,
            I => \N__23749\
        );

    \I__4447\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23746\
        );

    \I__4446\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23741\
        );

    \I__4445\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23741\
        );

    \I__4444\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23738\
        );

    \I__4443\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23735\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__23752\,
            I => \N__23730\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__23749\,
            I => \N__23730\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__23746\,
            I => \POWERLED.dutycycle\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__23741\,
            I => \POWERLED.dutycycle\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__23738\,
            I => \POWERLED.dutycycle\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__23735\,
            I => \POWERLED.dutycycle\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__23730\,
            I => \POWERLED.dutycycle\
        );

    \I__4435\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23716\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__23716\,
            I => \POWERLED.count_off_1_sqmuxa\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__23713\,
            I => \POWERLED.g0_9_1_cascade_\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__23710\,
            I => \POWERLED.dutycycle_fb_15_4_0_cascade_\
        );

    \I__4431\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23704\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__23704\,
            I => \POWERLED.dutycycle_fb_15_0\
        );

    \I__4429\ : CascadeMux
    port map (
            O => \N__23701\,
            I => \POWERLED.dutycycle_en_14_cascade_\
        );

    \I__4428\ : SRMux
    port map (
            O => \N__23698\,
            I => \N__23692\
        );

    \I__4427\ : SRMux
    port map (
            O => \N__23697\,
            I => \N__23689\
        );

    \I__4426\ : SRMux
    port map (
            O => \N__23696\,
            I => \N__23686\
        );

    \I__4425\ : SRMux
    port map (
            O => \N__23695\,
            I => \N__23682\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__23692\,
            I => \N__23677\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__23689\,
            I => \N__23677\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__23686\,
            I => \N__23674\
        );

    \I__4421\ : SRMux
    port map (
            O => \N__23685\,
            I => \N__23671\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__23682\,
            I => \N__23665\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__23677\,
            I => \N__23661\
        );

    \I__4418\ : Span4Mux_v
    port map (
            O => \N__23674\,
            I => \N__23656\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__23671\,
            I => \N__23656\
        );

    \I__4416\ : SRMux
    port map (
            O => \N__23670\,
            I => \N__23653\
        );

    \I__4415\ : SRMux
    port map (
            O => \N__23669\,
            I => \N__23650\
        );

    \I__4414\ : SRMux
    port map (
            O => \N__23668\,
            I => \N__23647\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__23665\,
            I => \N__23643\
        );

    \I__4412\ : SRMux
    port map (
            O => \N__23664\,
            I => \N__23640\
        );

    \I__4411\ : Span4Mux_v
    port map (
            O => \N__23661\,
            I => \N__23637\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__23656\,
            I => \N__23634\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__23653\,
            I => \N__23631\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23628\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23625\
        );

    \I__4406\ : SRMux
    port map (
            O => \N__23646\,
            I => \N__23622\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__23643\,
            I => \N__23617\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23617\
        );

    \I__4403\ : Sp12to4
    port map (
            O => \N__23637\,
            I => \N__23612\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__23634\,
            I => \N__23607\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__23631\,
            I => \N__23607\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__23628\,
            I => \N__23600\
        );

    \I__4399\ : Span4Mux_h
    port map (
            O => \N__23625\,
            I => \N__23600\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__23622\,
            I => \N__23600\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__23617\,
            I => \N__23597\
        );

    \I__4396\ : SRMux
    port map (
            O => \N__23616\,
            I => \N__23594\
        );

    \I__4395\ : SRMux
    port map (
            O => \N__23615\,
            I => \N__23591\
        );

    \I__4394\ : Odrv12
    port map (
            O => \N__23612\,
            I => \POWERLED.func_m2_0_a2_isoZ0\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__23607\,
            I => \POWERLED.func_m2_0_a2_isoZ0\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__23600\,
            I => \POWERLED.func_m2_0_a2_isoZ0\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__23597\,
            I => \POWERLED.func_m2_0_a2_isoZ0\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__23594\,
            I => \POWERLED.func_m2_0_a2_isoZ0\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__23591\,
            I => \POWERLED.func_m2_0_a2_isoZ0\
        );

    \I__4388\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23569\
        );

    \I__4387\ : InMux
    port map (
            O => \N__23577\,
            I => \N__23569\
        );

    \I__4386\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23569\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__23569\,
            I => \POWERLED.dutycycle_eena_14_0Z0Z_0\
        );

    \I__4384\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23563\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__23563\,
            I => \N__23560\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__23560\,
            I => \POWERLED.dutycycle_fb_15_1\
        );

    \I__4381\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23554\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__23554\,
            I => \POWERLED.g1_0\
        );

    \I__4379\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23548\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__23548\,
            I => \N__23545\
        );

    \I__4377\ : Odrv12
    port map (
            O => \N__23545\,
            I => \POWERLED.g1\
        );

    \I__4376\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23539\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__23539\,
            I => \POWERLED.dutycycle_fb_15_2_0\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__23536\,
            I => \N__23529\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23524\
        );

    \I__4372\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23524\
        );

    \I__4371\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23521\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23518\
        );

    \I__4369\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23515\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__23524\,
            I => \SUSWARN_N_rep1\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__23521\,
            I => \SUSWARN_N_rep1\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__23518\,
            I => \SUSWARN_N_rep1\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__23515\,
            I => \SUSWARN_N_rep1\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__23506\,
            I => \POWERLED.N_340_cascade_\
        );

    \I__4363\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__23500\,
            I => \N__23497\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__23497\,
            I => \POWERLED.func_state_RNIRAVV2Z0Z_0\
        );

    \I__4360\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23488\
        );

    \I__4358\ : Span4Mux_v
    port map (
            O => \N__23488\,
            I => \N__23485\
        );

    \I__4357\ : Sp12to4
    port map (
            O => \N__23485\,
            I => \N__23482\
        );

    \I__4356\ : Odrv12
    port map (
            O => \N__23482\,
            I => \POWERLED.m18_e_5\
        );

    \I__4355\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23476\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__23476\,
            I => \POWERLED.m18_e_6\
        );

    \I__4353\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23470\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__23470\,
            I => \POWERLED.func_m2_0_a2Z0Z_0\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__23467\,
            I => \POWERLED.func_m2_0_a2Z0Z_0_cascade_\
        );

    \I__4350\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23452\
        );

    \I__4349\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23452\
        );

    \I__4348\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23449\
        );

    \I__4347\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23444\
        );

    \I__4346\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23444\
        );

    \I__4345\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23441\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23438\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__23457\,
            I => \N__23435\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23432\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__23449\,
            I => \N__23427\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23427\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23422\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23422\
        );

    \I__4337\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23419\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__23432\,
            I => \N__23416\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__23427\,
            I => \N__23413\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__23422\,
            I => \N__23408\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23408\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__23416\,
            I => \POWERLED.count_clk_RNI2O4A1_0Z0Z_10\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__23413\,
            I => \POWERLED.count_clk_RNI2O4A1_0Z0Z_10\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__23408\,
            I => \POWERLED.count_clk_RNI2O4A1_0Z0Z_10\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__23401\,
            I => \POWERLED.func_state_RNI91IA4_0Z0Z_1_cascade_\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23398\,
            I => \N__23395\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__23395\,
            I => \POWERLED.func_state_1_m2_0\
        );

    \I__4326\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23386\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23386\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__23386\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__23383\,
            I => \POWERLED.func_state_1_m2_0_cascade_\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__23380\,
            I => \N__23377\
        );

    \I__4321\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23366\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23366\
        );

    \I__4319\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23361\
        );

    \I__4318\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23361\
        );

    \I__4317\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23358\
        );

    \I__4316\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23353\
        );

    \I__4315\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23353\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__23366\,
            I => \N__23350\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__23361\,
            I => \N__23347\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__23358\,
            I => \N__23342\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23339\
        );

    \I__4310\ : Span4Mux_h
    port map (
            O => \N__23350\,
            I => \N__23336\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__23347\,
            I => \N__23333\
        );

    \I__4308\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23330\
        );

    \I__4307\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23327\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__23342\,
            I => \POWERLED.N_335\
        );

    \I__4305\ : Odrv12
    port map (
            O => \N__23339\,
            I => \POWERLED.N_335\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__23336\,
            I => \POWERLED.N_335\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__23333\,
            I => \POWERLED.N_335\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__23330\,
            I => \POWERLED.N_335\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__23327\,
            I => \POWERLED.N_335\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__23314\,
            I => \POWERLED.func_state_RNI2O4A1Z0Z_1_cascade_\
        );

    \I__4299\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23305\
        );

    \I__4298\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23305\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__23305\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__23302\,
            I => \N__23299\
        );

    \I__4295\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__4294\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23293\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__23293\,
            I => \POWERLED.dutycycle_en_9\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__23290\,
            I => \POWERLED.func_state_RNI2O4A1_1Z0Z_1_cascade_\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__4290\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23281\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__23281\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\
        );

    \I__4288\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23275\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__23275\,
            I => \N__23270\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__23274\,
            I => \N__23262\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__23273\,
            I => \N__23257\
        );

    \I__4284\ : Span4Mux_v
    port map (
            O => \N__23270\,
            I => \N__23254\
        );

    \I__4283\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23251\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__23268\,
            I => \N__23248\
        );

    \I__4281\ : InMux
    port map (
            O => \N__23267\,
            I => \N__23244\
        );

    \I__4280\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23241\
        );

    \I__4279\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23230\
        );

    \I__4278\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23230\
        );

    \I__4277\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23230\
        );

    \I__4276\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23230\
        );

    \I__4275\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23230\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__23254\,
            I => \N__23224\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23224\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23219\
        );

    \I__4271\ : InMux
    port map (
            O => \N__23247\,
            I => \N__23219\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__23244\,
            I => \N__23214\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__23241\,
            I => \N__23214\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__23230\,
            I => \N__23211\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__23229\,
            I => \N__23208\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__23224\,
            I => \N__23205\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23202\
        );

    \I__4264\ : Span4Mux_h
    port map (
            O => \N__23214\,
            I => \N__23199\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__23211\,
            I => \N__23196\
        );

    \I__4262\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23193\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__23205\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4260\ : Odrv12
    port map (
            O => \N__23202\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__23199\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__23196\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__23193\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__23182\,
            I => \POWERLED.dutycycleZ0Z_11_cascade_\
        );

    \I__4255\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__23176\,
            I => \POWERLED.un1_clk_100khz_42_and_i_0_0\
        );

    \I__4253\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23167\
        );

    \I__4252\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23167\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__23167\,
            I => \N__23163\
        );

    \I__4250\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23159\
        );

    \I__4249\ : Span12Mux_s7_h
    port map (
            O => \N__23163\,
            I => \N__23156\
        );

    \I__4248\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23153\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__23159\,
            I => \POWERLED.func_state_RNI2O4A1Z0Z_1\
        );

    \I__4246\ : Odrv12
    port map (
            O => \N__23156\,
            I => \POWERLED.func_state_RNI2O4A1Z0Z_1\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__23153\,
            I => \POWERLED.func_state_RNI2O4A1Z0Z_1\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__23146\,
            I => \POWERLED.un1_clk_100khz_47_and_i_0_0_cascade_\
        );

    \I__4243\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23137\
        );

    \I__4242\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23137\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__23137\,
            I => \N__23133\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__23136\,
            I => \N__23130\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__23133\,
            I => \N__23126\
        );

    \I__4238\ : InMux
    port map (
            O => \N__23130\,
            I => \N__23121\
        );

    \I__4237\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23121\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__23126\,
            I => \POWERLED.N_399_N\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__23121\,
            I => \POWERLED.N_399_N\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__23116\,
            I => \N__23112\
        );

    \I__4233\ : InMux
    port map (
            O => \N__23115\,
            I => \N__23109\
        );

    \I__4232\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23106\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__23101\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__23106\,
            I => \N__23101\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__23098\,
            I => \POWERLED.dutycycle_en_11\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \POWERLED.N_2216_i_cascade_\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__23092\,
            I => \POWERLED.func_state_1_m2s2_i_1_cascade_\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__23089\,
            I => \N__23085\
        );

    \I__4224\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23080\
        );

    \I__4223\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23080\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__23077\,
            I => \POWERLED.N_160\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__23074\,
            I => \N__23065\
        );

    \I__4219\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23060\
        );

    \I__4218\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23060\
        );

    \I__4217\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23057\
        );

    \I__4216\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23052\
        );

    \I__4215\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23052\
        );

    \I__4214\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23047\
        );

    \I__4213\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23047\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__23060\,
            I => \N__23044\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23037\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23037\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__23047\,
            I => \N__23037\
        );

    \I__4208\ : Span4Mux_h
    port map (
            O => \N__23044\,
            I => \N__23032\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__23037\,
            I => \N__23032\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__23032\,
            I => \POWERLED.N_3_0\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__23029\,
            I => \slp_s3n_signal_cascade_\
        );

    \I__4204\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23020\
        );

    \I__4203\ : InMux
    port map (
            O => \N__23025\,
            I => \N__23020\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__23020\,
            I => \POWERLED.N_183\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__23017\,
            I => \POWERLED.func_state_RNIZ0Z_1_cascade_\
        );

    \I__4200\ : InMux
    port map (
            O => \N__23014\,
            I => \N__22994\
        );

    \I__4199\ : InMux
    port map (
            O => \N__23013\,
            I => \N__22994\
        );

    \I__4198\ : InMux
    port map (
            O => \N__23012\,
            I => \N__22994\
        );

    \I__4197\ : InMux
    port map (
            O => \N__23011\,
            I => \N__22987\
        );

    \I__4196\ : InMux
    port map (
            O => \N__23010\,
            I => \N__22987\
        );

    \I__4195\ : InMux
    port map (
            O => \N__23009\,
            I => \N__22987\
        );

    \I__4194\ : InMux
    port map (
            O => \N__23008\,
            I => \N__22978\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23007\,
            I => \N__22978\
        );

    \I__4192\ : InMux
    port map (
            O => \N__23006\,
            I => \N__22978\
        );

    \I__4191\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22978\
        );

    \I__4190\ : InMux
    port map (
            O => \N__23004\,
            I => \N__22969\
        );

    \I__4189\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22969\
        );

    \I__4188\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22969\
        );

    \I__4187\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22969\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__22994\,
            I => \POWERLED.N_162_i\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__22987\,
            I => \POWERLED.N_162_i\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__22978\,
            I => \POWERLED.N_162_i\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__22969\,
            I => \POWERLED.N_162_i\
        );

    \I__4182\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__22957\,
            I => \POWERLED.count_off_0_1\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__4179\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__22948\,
            I => \POWERLED.count_off_RNIZ0Z_1\
        );

    \I__4177\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22942\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__22942\,
            I => \N__22938\
        );

    \I__4175\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22935\
        );

    \I__4174\ : Span4Mux_h
    port map (
            O => \N__22938\,
            I => \N__22932\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__22935\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__22932\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__22927\,
            I => \POWERLED.count_offZ0Z_1_cascade_\
        );

    \I__4170\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__22921\,
            I => \POWERLED.un34_clk_100khz_10\
        );

    \I__4168\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22912\
        );

    \I__4166\ : Span12Mux_v
    port map (
            O => \N__22912\,
            I => \N__22909\
        );

    \I__4165\ : Odrv12
    port map (
            O => \N__22909\,
            I => \POWERLED.un34_clk_100khz_8\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__22906\,
            I => \POWERLED.un34_clk_100khz_9_cascade_\
        );

    \I__4163\ : InMux
    port map (
            O => \N__22903\,
            I => \N__22900\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__22894\,
            I => \POWERLED.un34_clk_100khz_11\
        );

    \I__4159\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22888\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__22888\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__22885\,
            I => \POWERLED.N_220_cascade_\
        );

    \I__4156\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22878\
        );

    \I__4155\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22875\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__22878\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__22875\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__22870\,
            I => \POWERLED.N_304_cascade_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22867\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__4150\ : InMux
    port map (
            O => \N__22864\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__4149\ : InMux
    port map (
            O => \N__22861\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__4148\ : InMux
    port map (
            O => \N__22858\,
            I => \bfn_8_5_0_\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__22855\,
            I => \POWERLED.count_off_RNIBQDB2Z0Z_0_cascade_\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__22852\,
            I => \POWERLED.count_offZ0Z_0_cascade_\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__22849\,
            I => \POWERLED.count_off_RNIZ0Z_1_cascade_\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__4143\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22840\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__22840\,
            I => \N__22834\
        );

    \I__4141\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22831\
        );

    \I__4140\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22826\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22837\,
            I => \N__22826\
        );

    \I__4138\ : Span4Mux_h
    port map (
            O => \N__22834\,
            I => \N__22823\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__22831\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__22826\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__22823\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__4134\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22813\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__22813\,
            I => \POWERLED.count_off_0_0\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22810\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__4131\ : InMux
    port map (
            O => \N__22807\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__4130\ : InMux
    port map (
            O => \N__22804\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__4129\ : InMux
    port map (
            O => \N__22801\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22798\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22795\,
            I => \bfn_8_4_0_\
        );

    \I__4126\ : InMux
    port map (
            O => \N__22792\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__4125\ : InMux
    port map (
            O => \N__22789\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__4124\ : InMux
    port map (
            O => \N__22786\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__4123\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22777\
        );

    \I__4122\ : InMux
    port map (
            O => \N__22782\,
            I => \N__22777\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__22777\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__4120\ : InMux
    port map (
            O => \N__22774\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22768\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22768\,
            I => \PCH_PWRGD.un2_count_1_axb_13\
        );

    \I__4117\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22758\
        );

    \I__4116\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22758\
        );

    \I__4115\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22755\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__22758\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__22755\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__4112\ : InMux
    port map (
            O => \N__22750\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__4111\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__22744\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__4109\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22735\
        );

    \I__4108\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22735\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22732\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__22732\,
            I => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\
        );

    \I__4105\ : InMux
    port map (
            O => \N__22729\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__4104\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__22723\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__4102\ : InMux
    port map (
            O => \N__22720\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__4101\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22711\
        );

    \I__4100\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22711\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__22711\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22704\
        );

    \I__4097\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22701\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__22704\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__22701\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__4094\ : InMux
    port map (
            O => \N__22696\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__4093\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22689\
        );

    \I__4092\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22686\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__22689\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22686\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__4089\ : InMux
    port map (
            O => \N__22681\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__4088\ : InMux
    port map (
            O => \N__22678\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__22675\,
            I => \N__22672\
        );

    \I__4086\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22668\
        );

    \I__4085\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22665\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__22668\,
            I => \PCH_PWRGD.un2_count_1_axb_4\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__22665\,
            I => \PCH_PWRGD.un2_count_1_axb_4\
        );

    \I__4082\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22654\
        );

    \I__4081\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22654\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__22654\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22651\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__4078\ : InMux
    port map (
            O => \N__22648\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__4077\ : InMux
    port map (
            O => \N__22645\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__4076\ : InMux
    port map (
            O => \N__22642\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__4075\ : InMux
    port map (
            O => \N__22639\,
            I => \PCH_PWRGD.un2_count_1_cry_7\
        );

    \I__4074\ : InMux
    port map (
            O => \N__22636\,
            I => \bfn_8_2_0_\
        );

    \I__4073\ : InMux
    port map (
            O => \N__22633\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__4072\ : InMux
    port map (
            O => \N__22630\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__4071\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22624\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__22624\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__22621\,
            I => \N__22618\
        );

    \I__4068\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22615\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__22615\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__4066\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22609\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__22609\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \N__22603\
        );

    \I__4063\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22593\
        );

    \I__4062\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22593\
        );

    \I__4061\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22593\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22590\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__22593\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__22590\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__22585\,
            I => \N__22581\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22573\
        );

    \I__4055\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22573\
        );

    \I__4054\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22573\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__22573\,
            I => \G_2078\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__4051\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22564\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__22564\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__4049\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22558\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__22558\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__4047\ : InMux
    port map (
            O => \N__22555\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22549\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22546\
        );

    \I__4044\ : Span4Mux_v
    port map (
            O => \N__22546\,
            I => \N__22543\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__22540\,
            I => \POWERLED.un85_clk_100khz_0\
        );

    \I__4041\ : IoInMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__22534\,
            I => \G_9\
        );

    \I__4039\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__22528\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__4037\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22516\
        );

    \I__4036\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22516\
        );

    \I__4035\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22516\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__22516\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__4033\ : InMux
    port map (
            O => \N__22513\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__4031\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22504\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__22498\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__4027\ : InMux
    port map (
            O => \N__22495\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__4026\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22489\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__22489\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__4024\ : InMux
    port map (
            O => \N__22486\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__4022\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22477\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__22477\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__4020\ : InMux
    port map (
            O => \N__22474\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__4019\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__22468\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__4016\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22454\
        );

    \I__4015\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22454\
        );

    \I__4014\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22451\
        );

    \I__4013\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22448\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__22454\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__22451\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__22448\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__4009\ : InMux
    port map (
            O => \N__22441\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__22438\,
            I => \N__22434\
        );

    \I__4007\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22426\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22426\
        );

    \I__4005\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22426\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__22426\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__4002\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22417\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__22417\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__4000\ : InMux
    port map (
            O => \N__22414\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__3999\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__22408\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__3997\ : InMux
    port map (
            O => \N__22405\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \POWERLED.mult1_un159_sum_s_7_cascade_\
        );

    \I__3995\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22393\
        );

    \I__3993\ : Span4Mux_v
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__3992\ : Span4Mux_h
    port map (
            O => \N__22390\,
            I => \N__22387\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__22387\,
            I => \POWERLED.un85_clk_100khz_1\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__22384\,
            I => \N__22379\
        );

    \I__3989\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22373\
        );

    \I__3988\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22370\
        );

    \I__3987\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22367\
        );

    \I__3986\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22361\
        );

    \I__3985\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22361\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__22376\,
            I => \N__22358\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__22373\,
            I => \N__22353\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22350\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22347\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22344\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__22361\,
            I => \N__22339\
        );

    \I__3978\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22334\
        );

    \I__3977\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22334\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__22356\,
            I => \N__22331\
        );

    \I__3975\ : Span4Mux_v
    port map (
            O => \N__22353\,
            I => \N__22328\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__22350\,
            I => \N__22323\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__22347\,
            I => \N__22323\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22319\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22314\
        );

    \I__3970\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22314\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__22339\,
            I => \N__22309\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22309\
        );

    \I__3967\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22306\
        );

    \I__3966\ : Span4Mux_h
    port map (
            O => \N__22328\,
            I => \N__22301\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__22323\,
            I => \N__22301\
        );

    \I__3964\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22298\
        );

    \I__3963\ : Span12Mux_s4_v
    port map (
            O => \N__22319\,
            I => \N__22289\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__22314\,
            I => \N__22289\
        );

    \I__3961\ : Sp12to4
    port map (
            O => \N__22309\,
            I => \N__22289\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__22306\,
            I => \N__22289\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__22301\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__22298\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3957\ : Odrv12
    port map (
            O => \N__22289\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__3955\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22276\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__3953\ : Span12Mux_s8_h
    port map (
            O => \N__22273\,
            I => \N__22270\
        );

    \I__3952\ : Odrv12
    port map (
            O => \N__22270\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__3951\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22264\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__22264\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__3949\ : InMux
    port map (
            O => \N__22261\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__22258\,
            I => \N__22255\
        );

    \I__3947\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22252\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__22252\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__3945\ : InMux
    port map (
            O => \N__22249\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__3944\ : InMux
    port map (
            O => \N__22246\,
            I => \N__22243\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__22243\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__3942\ : InMux
    port map (
            O => \N__22240\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__3941\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__22234\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__3939\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__22228\,
            I => \N__22225\
        );

    \I__3937\ : Span4Mux_s2_v
    port map (
            O => \N__22225\,
            I => \N__22220\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__22224\,
            I => \N__22217\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__22223\,
            I => \N__22214\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__22220\,
            I => \N__22210\
        );

    \I__3933\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22207\
        );

    \I__3932\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22204\
        );

    \I__3931\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22201\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__22210\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__22207\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__22204\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__22201\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3926\ : InMux
    port map (
            O => \N__22192\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__3925\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__22186\,
            I => \N__22183\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__22183\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__22180\,
            I => \N__22176\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__22179\,
            I => \N__22172\
        );

    \I__3920\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22165\
        );

    \I__3919\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22165\
        );

    \I__3918\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22165\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__22165\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__3916\ : InMux
    port map (
            O => \N__22162\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__3915\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22156\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__22156\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__3913\ : InMux
    port map (
            O => \N__22153\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__22150\,
            I => \POWERLED.mult1_un152_sum_s_8_cascade_\
        );

    \I__3911\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22136\
        );

    \I__3910\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22133\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__22145\,
            I => \N__22130\
        );

    \I__3908\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22126\
        );

    \I__3907\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22121\
        );

    \I__3906\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22121\
        );

    \I__3905\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22118\
        );

    \I__3904\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22113\
        );

    \I__3903\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22113\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__22136\,
            I => \N__22107\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__22133\,
            I => \N__22107\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22130\,
            I => \N__22103\
        );

    \I__3899\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22100\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22095\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22095\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22090\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22087\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__22112\,
            I => \N__22083\
        );

    \I__3893\ : Sp12to4
    port map (
            O => \N__22107\,
            I => \N__22080\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__22106\,
            I => \N__22077\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22074\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22069\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__22095\,
            I => \N__22069\
        );

    \I__3888\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22064\
        );

    \I__3887\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22064\
        );

    \I__3886\ : Span4Mux_v
    port map (
            O => \N__22090\,
            I => \N__22059\
        );

    \I__3885\ : Span4Mux_s2_h
    port map (
            O => \N__22087\,
            I => \N__22059\
        );

    \I__3884\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22056\
        );

    \I__3883\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22053\
        );

    \I__3882\ : Span12Mux_v
    port map (
            O => \N__22080\,
            I => \N__22050\
        );

    \I__3881\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22047\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__22074\,
            I => \N__22044\
        );

    \I__3879\ : Span4Mux_v
    port map (
            O => \N__22069\,
            I => \N__22033\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__22064\,
            I => \N__22033\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__22059\,
            I => \N__22033\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__22056\,
            I => \N__22033\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__22053\,
            I => \N__22033\
        );

    \I__3874\ : Odrv12
    port map (
            O => \N__22050\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__22047\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__22044\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__22033\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__22024\,
            I => \G_155_cascade_\
        );

    \I__3869\ : InMux
    port map (
            O => \N__22021\,
            I => \N__22018\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__22018\,
            I => \POWERLED.N_73\
        );

    \I__3867\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22009\
        );

    \I__3866\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22009\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__22009\,
            I => \POWERLED.dutycycle_eena_1\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__22006\,
            I => \POWERLED.N_73_cascade_\
        );

    \I__3863\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21997\
        );

    \I__3862\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21997\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__21997\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__21994\,
            I => \N__21991\
        );

    \I__3859\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21988\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__21988\,
            I => \POWERLED.N_277\
        );

    \I__3857\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21982\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__21982\,
            I => \N__21979\
        );

    \I__3855\ : Odrv12
    port map (
            O => \N__21979\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\
        );

    \I__3854\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21973\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__21973\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_2\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__21970\,
            I => \POWERLED.dutycycle_1_0_iv_0_1_5_cascade_\
        );

    \I__3851\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21958\
        );

    \I__3850\ : InMux
    port map (
            O => \N__21966\,
            I => \N__21958\
        );

    \I__3849\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21958\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__21958\,
            I => \SUSWARN_N_fast\
        );

    \I__3847\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21946\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__21954\,
            I => \N__21943\
        );

    \I__3845\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21940\
        );

    \I__3844\ : InMux
    port map (
            O => \N__21952\,
            I => \N__21936\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__21951\,
            I => \N__21933\
        );

    \I__3842\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21930\
        );

    \I__3841\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21927\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__21946\,
            I => \N__21922\
        );

    \I__3839\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21919\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__21940\,
            I => \N__21916\
        );

    \I__3837\ : InMux
    port map (
            O => \N__21939\,
            I => \N__21913\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__21936\,
            I => \N__21910\
        );

    \I__3835\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21907\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21904\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__21927\,
            I => \N__21901\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__21926\,
            I => \N__21897\
        );

    \I__3831\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21885\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__21922\,
            I => \N__21880\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21880\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__21916\,
            I => \N__21875\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__21913\,
            I => \N__21875\
        );

    \I__3826\ : Span4Mux_v
    port map (
            O => \N__21910\,
            I => \N__21870\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__21907\,
            I => \N__21870\
        );

    \I__3824\ : Span4Mux_v
    port map (
            O => \N__21904\,
            I => \N__21865\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__21901\,
            I => \N__21865\
        );

    \I__3822\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21858\
        );

    \I__3821\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21858\
        );

    \I__3820\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21858\
        );

    \I__3819\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21847\
        );

    \I__3818\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21847\
        );

    \I__3817\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21847\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21847\
        );

    \I__3815\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21847\
        );

    \I__3814\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21840\
        );

    \I__3813\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21840\
        );

    \I__3812\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21840\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__21885\,
            I => \N__21835\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__21880\,
            I => \N__21835\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__21875\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__21870\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__21865\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__21858\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__21847\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__21840\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__21835\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3802\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__21817\,
            I => \POWERLED.m18_e_0\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__21814\,
            I => \N__21810\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__21813\,
            I => \N__21797\
        );

    \I__3798\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21793\
        );

    \I__3797\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21788\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21788\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21785\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__21806\,
            I => \N__21781\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21778\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__21804\,
            I => \N__21772\
        );

    \I__3791\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21767\
        );

    \I__3790\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21767\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__21801\,
            I => \N__21763\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \N__21759\
        );

    \I__3787\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21756\
        );

    \I__3786\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21753\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21750\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21747\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21744\
        );

    \I__3782\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21741\
        );

    \I__3781\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21738\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__21778\,
            I => \N__21735\
        );

    \I__3779\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21730\
        );

    \I__3778\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21730\
        );

    \I__3777\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21723\
        );

    \I__3776\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21723\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__21767\,
            I => \N__21720\
        );

    \I__3774\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21711\
        );

    \I__3773\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21711\
        );

    \I__3772\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21711\
        );

    \I__3771\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21711\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__21756\,
            I => \N__21708\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21705\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__21750\,
            I => \N__21694\
        );

    \I__3767\ : Span4Mux_v
    port map (
            O => \N__21747\,
            I => \N__21694\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__21744\,
            I => \N__21694\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21694\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21694\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__21735\,
            I => \N__21689\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__21730\,
            I => \N__21689\
        );

    \I__3761\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21684\
        );

    \I__3760\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21684\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21681\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__21720\,
            I => \N__21676\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__21711\,
            I => \N__21676\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__21708\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__21705\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__21694\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__21689\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__21684\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__21681\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__21676\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3749\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__21658\,
            I => \POWERLED.un1_dutycycle_94_cry_4_c_RNI919HZ0Z1\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__21655\,
            I => \POWERLED.dutycycle_1_0_5_cascade_\
        );

    \I__3746\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21648\
        );

    \I__3745\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21645\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__21648\,
            I => \POWERLED.func_state_RNIT69J5Z0Z_1\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__21645\,
            I => \POWERLED.func_state_RNIT69J5Z0Z_1\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__21640\,
            I => \POWERLED.N_366_cascade_\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__21637\,
            I => \POWERLED.dutycycle_RNI2O4A1Z0Z_6_cascade_\
        );

    \I__3740\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__21631\,
            I => \POWERLED.dutycycle_RNI2O4A1_2Z0Z_2\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__21628\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m1_cascade_\
        );

    \I__3737\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__21622\,
            I => \N__21617\
        );

    \I__3735\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21612\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21612\
        );

    \I__3733\ : Span4Mux_v
    port map (
            O => \N__21617\,
            I => \N__21607\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__21612\,
            I => \N__21607\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__21607\,
            I => \POWERLED.dutycycle_RNIZ0Z_5\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__21604\,
            I => \POWERLED.func_state_RNI_0Z0Z_0_cascade_\
        );

    \I__3729\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21598\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__21598\,
            I => \POWERLED.func_state_RNI68EU3Z0Z_1\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__3725\ : Span4Mux_h
    port map (
            O => \N__21589\,
            I => \N__21586\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__21586\,
            I => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21577\
        );

    \I__3722\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21577\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__21577\,
            I => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\
        );

    \I__3720\ : InMux
    port map (
            O => \N__21574\,
            I => \POWERLED.un1_dutycycle_94_cry_10\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21571\,
            I => \POWERLED.un1_dutycycle_94_cry_11\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21563\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21559\
        );

    \I__3716\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21556\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21552\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__21562\,
            I => \N__21548\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__21559\,
            I => \N__21544\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__21556\,
            I => \N__21541\
        );

    \I__3711\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21538\
        );

    \I__3710\ : Span4Mux_v
    port map (
            O => \N__21552\,
            I => \N__21535\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21530\
        );

    \I__3708\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21530\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__21547\,
            I => \N__21525\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__21544\,
            I => \N__21518\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__21541\,
            I => \N__21518\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__21538\,
            I => \N__21518\
        );

    \I__3703\ : Span4Mux_h
    port map (
            O => \N__21535\,
            I => \N__21513\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__21530\,
            I => \N__21513\
        );

    \I__3701\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21510\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21507\
        );

    \I__3699\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21504\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__21518\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__21513\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__21510\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__21507\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__21504\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3693\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21487\
        );

    \I__3692\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21487\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__21487\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21484\,
            I => \POWERLED.un1_dutycycle_94_cry_12\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21475\
        );

    \I__3688\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21475\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__21472\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__3685\ : InMux
    port map (
            O => \N__21469\,
            I => \POWERLED.un1_dutycycle_94_cry_13\
        );

    \I__3684\ : InMux
    port map (
            O => \N__21466\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__3683\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21457\
        );

    \I__3682\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21457\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21454\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__21454\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__3679\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21446\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__21450\,
            I => \N__21443\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__21449\,
            I => \N__21440\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__21446\,
            I => \N__21435\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21430\
        );

    \I__3674\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21427\
        );

    \I__3673\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21424\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__21438\,
            I => \N__21421\
        );

    \I__3671\ : Span4Mux_v
    port map (
            O => \N__21435\,
            I => \N__21418\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21415\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21412\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21409\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21404\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21404\
        );

    \I__3665\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21401\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__21418\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__21415\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__21412\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3661\ : Odrv12
    port map (
            O => \N__21409\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__21404\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__21401\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__21388\,
            I => \N__21382\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__21387\,
            I => \N__21377\
        );

    \I__3656\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21374\
        );

    \I__3655\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21369\
        );

    \I__3654\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21369\
        );

    \I__3653\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21362\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21362\
        );

    \I__3651\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21362\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__21374\,
            I => \N__21355\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__21369\,
            I => \N__21352\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21349\
        );

    \I__3647\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21340\
        );

    \I__3646\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21340\
        );

    \I__3645\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21340\
        );

    \I__3644\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21340\
        );

    \I__3643\ : Span4Mux_h
    port map (
            O => \N__21355\,
            I => \N__21335\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__21352\,
            I => \N__21335\
        );

    \I__3641\ : Odrv12
    port map (
            O => \N__21349\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__21340\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__21335\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21322\
        );

    \I__3637\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21322\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__21322\,
            I => \N__21319\
        );

    \I__3635\ : Odrv12
    port map (
            O => \N__21319\,
            I => \POWERLED.N_115_f0_1\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__21316\,
            I => \N__21311\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__21315\,
            I => \N__21308\
        );

    \I__3632\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21302\
        );

    \I__3631\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21302\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21293\
        );

    \I__3629\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21290\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__21302\,
            I => \N__21287\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__21301\,
            I => \N__21284\
        );

    \I__3626\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21281\
        );

    \I__3625\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21275\
        );

    \I__3624\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21268\
        );

    \I__3623\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21268\
        );

    \I__3622\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21268\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__21293\,
            I => \N__21264\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__21290\,
            I => \N__21259\
        );

    \I__3619\ : Span4Mux_v
    port map (
            O => \N__21287\,
            I => \N__21259\
        );

    \I__3618\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21256\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__21281\,
            I => \N__21253\
        );

    \I__3616\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21250\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__21279\,
            I => \N__21246\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \N__21243\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__21275\,
            I => \N__21237\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21234\
        );

    \I__3611\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21231\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__21264\,
            I => \N__21228\
        );

    \I__3609\ : Span4Mux_h
    port map (
            O => \N__21259\,
            I => \N__21223\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__21256\,
            I => \N__21223\
        );

    \I__3607\ : Span4Mux_h
    port map (
            O => \N__21253\,
            I => \N__21218\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21218\
        );

    \I__3605\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21213\
        );

    \I__3604\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21213\
        );

    \I__3603\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21204\
        );

    \I__3602\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21204\
        );

    \I__3601\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21204\
        );

    \I__3600\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21204\
        );

    \I__3599\ : Span4Mux_h
    port map (
            O => \N__21237\,
            I => \N__21199\
        );

    \I__3598\ : Span4Mux_v
    port map (
            O => \N__21234\,
            I => \N__21199\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__21231\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__21228\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__21223\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__21218\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__21213\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__21204\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__21199\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3590\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21178\
        );

    \I__3589\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21178\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21175\
        );

    \I__3587\ : Span4Mux_h
    port map (
            O => \N__21175\,
            I => \N__21172\
        );

    \I__3586\ : Odrv4
    port map (
            O => \N__21172\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI765BZ0Z1\
        );

    \I__3585\ : InMux
    port map (
            O => \N__21169\,
            I => \POWERLED.un1_dutycycle_94_cry_2\
        );

    \I__3584\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21163\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N__21159\
        );

    \I__3582\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21156\
        );

    \I__3581\ : Sp12to4
    port map (
            O => \N__21159\,
            I => \N__21151\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21151\
        );

    \I__3579\ : Odrv12
    port map (
            O => \N__21151\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI886BZ0Z1\
        );

    \I__3578\ : InMux
    port map (
            O => \N__21148\,
            I => \POWERLED.un1_dutycycle_94_cry_3\
        );

    \I__3577\ : InMux
    port map (
            O => \N__21145\,
            I => \POWERLED.un1_dutycycle_94_cry_4_cZ0\
        );

    \I__3576\ : InMux
    port map (
            O => \N__21142\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3575\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21132\
        );

    \I__3574\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21132\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__21137\,
            I => \N__21126\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__21118\
        );

    \I__3571\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21115\
        );

    \I__3570\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21110\
        );

    \I__3569\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21110\
        );

    \I__3568\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21095\
        );

    \I__3567\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21095\
        );

    \I__3566\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21095\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__21123\,
            I => \N__21092\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__21122\,
            I => \N__21089\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__21121\,
            I => \N__21086\
        );

    \I__3562\ : Span4Mux_h
    port map (
            O => \N__21118\,
            I => \N__21083\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__21115\,
            I => \N__21078\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__21110\,
            I => \N__21078\
        );

    \I__3559\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21073\
        );

    \I__3558\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21073\
        );

    \I__3557\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21068\
        );

    \I__3556\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21068\
        );

    \I__3555\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21054\
        );

    \I__3554\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21054\
        );

    \I__3553\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21054\
        );

    \I__3552\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21051\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21048\
        );

    \I__3550\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21045\
        );

    \I__3549\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21040\
        );

    \I__3548\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21040\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__21083\,
            I => \N__21035\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__21078\,
            I => \N__21035\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21030\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21030\
        );

    \I__3543\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21023\
        );

    \I__3542\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21023\
        );

    \I__3541\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21023\
        );

    \I__3540\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21016\
        );

    \I__3539\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21016\
        );

    \I__3538\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21016\
        );

    \I__3537\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21013\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__21054\,
            I => \N__21010\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21003\
        );

    \I__3534\ : Span4Mux_s3_h
    port map (
            O => \N__21048\,
            I => \N__21003\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__21045\,
            I => \N__21003\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__21040\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__21035\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__21030\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__21023\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__21016\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__21013\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__21010\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__21003\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__3524\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20980\
        );

    \I__3523\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20980\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__20980\,
            I => \N__20977\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__20977\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4AZ0Z1\
        );

    \I__3520\ : InMux
    port map (
            O => \N__20974\,
            I => \POWERLED.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__20971\,
            I => \N__20965\
        );

    \I__3518\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20959\
        );

    \I__3517\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20952\
        );

    \I__3516\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20952\
        );

    \I__3515\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20952\
        );

    \I__3514\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20944\
        );

    \I__3513\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20944\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__20962\,
            I => \N__20934\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__20959\,
            I => \N__20928\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20925\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__20951\,
            I => \N__20921\
        );

    \I__3508\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20914\
        );

    \I__3507\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20914\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20910\
        );

    \I__3505\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20907\
        );

    \I__3504\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20898\
        );

    \I__3503\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20898\
        );

    \I__3502\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20898\
        );

    \I__3501\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20898\
        );

    \I__3500\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20895\
        );

    \I__3499\ : InMux
    port map (
            O => \N__20937\,
            I => \N__20892\
        );

    \I__3498\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20889\
        );

    \I__3497\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20882\
        );

    \I__3496\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20882\
        );

    \I__3495\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20882\
        );

    \I__3494\ : Span4Mux_h
    port map (
            O => \N__20928\,
            I => \N__20877\
        );

    \I__3493\ : Span4Mux_s3_h
    port map (
            O => \N__20925\,
            I => \N__20877\
        );

    \I__3492\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20868\
        );

    \I__3491\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20868\
        );

    \I__3490\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20868\
        );

    \I__3489\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20868\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20865\
        );

    \I__3487\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20862\
        );

    \I__3486\ : Span4Mux_h
    port map (
            O => \N__20910\,
            I => \N__20859\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__20907\,
            I => \N__20854\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__20898\,
            I => \N__20854\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__20895\,
            I => \N__20847\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__20892\,
            I => \N__20847\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20847\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__20882\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__20877\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__20868\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__20865\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__20862\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__20859\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3474\ : Odrv12
    port map (
            O => \N__20854\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3473\ : Odrv12
    port map (
            O => \N__20847\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20824\
        );

    \I__3471\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20824\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__3469\ : Odrv12
    port map (
            O => \N__20821\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNICGABZ0Z1\
        );

    \I__3468\ : InMux
    port map (
            O => \N__20818\,
            I => \bfn_7_8_0_\
        );

    \I__3467\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20802\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__20814\,
            I => \N__20799\
        );

    \I__3465\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20794\
        );

    \I__3464\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20794\
        );

    \I__3463\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20785\
        );

    \I__3462\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20785\
        );

    \I__3461\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20785\
        );

    \I__3460\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20785\
        );

    \I__3459\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20780\
        );

    \I__3458\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20780\
        );

    \I__3457\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20777\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__20802\,
            I => \N__20768\
        );

    \I__3455\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20765\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__20794\,
            I => \N__20759\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__20785\,
            I => \N__20756\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20751\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__20777\,
            I => \N__20751\
        );

    \I__3450\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20746\
        );

    \I__3449\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20746\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__20774\,
            I => \N__20743\
        );

    \I__3447\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20740\
        );

    \I__3446\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20735\
        );

    \I__3445\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20735\
        );

    \I__3444\ : Span4Mux_h
    port map (
            O => \N__20768\,
            I => \N__20732\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20729\
        );

    \I__3442\ : InMux
    port map (
            O => \N__20764\,
            I => \N__20722\
        );

    \I__3441\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20722\
        );

    \I__3440\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20722\
        );

    \I__3439\ : Span4Mux_v
    port map (
            O => \N__20759\,
            I => \N__20713\
        );

    \I__3438\ : Span4Mux_s3_h
    port map (
            O => \N__20756\,
            I => \N__20713\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__20751\,
            I => \N__20713\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20713\
        );

    \I__3435\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20710\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__20740\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__20735\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__20732\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__20729\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__20722\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__20713\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__20710\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3427\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20689\
        );

    \I__3426\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20689\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__20689\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\
        );

    \I__3424\ : InMux
    port map (
            O => \N__20686\,
            I => \POWERLED.un1_dutycycle_94_cry_8_cZ0\
        );

    \I__3423\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20677\
        );

    \I__3422\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20677\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__20677\,
            I => \N__20674\
        );

    \I__3420\ : Span4Mux_v
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__20671\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCBZ0Z1\
        );

    \I__3418\ : InMux
    port map (
            O => \N__20668\,
            I => \POWERLED.un1_dutycycle_94_cry_9\
        );

    \I__3417\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20659\
        );

    \I__3416\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20659\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20656\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__20656\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__20653\,
            I => \POWERLED.dutycycleZ1Z_6_cascade_\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_0_cascade_\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__3410\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20641\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__20641\,
            I => \POWERLED.un1_dutycycle_96_0_a3_0\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__20632\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_0\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__20629\,
            I => \POWERLED.un2_count_clk_17_0_cascade_\
        );

    \I__3404\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20623\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__20623\,
            I => \N__20620\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__20620\,
            I => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\
        );

    \I__3401\ : InMux
    port map (
            O => \N__20617\,
            I => \POWERLED.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__3400\ : InMux
    port map (
            O => \N__20614\,
            I => \POWERLED.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__20611\,
            I => \POWERLED.func_state_RNISKPU6Z0Z_0_cascade_\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20602\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20602\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__20602\,
            I => \POWERLED.count_off_1_13\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20596\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__20596\,
            I => \POWERLED.count_off_0_13\
        );

    \I__3393\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20587\
        );

    \I__3392\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20587\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__20587\,
            I => \POWERLED.count_off_1_14\
        );

    \I__3390\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__20581\,
            I => \POWERLED.count_off_0_14\
        );

    \I__3388\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20574\
        );

    \I__3387\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20571\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20574\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__20571\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2\
        );

    \I__3384\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20563\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__20563\,
            I => \POWERLED.count_off_0_15\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20557\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__20557\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__3380\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20550\
        );

    \I__3379\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20547\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__20550\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__20547\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__20542\,
            I => \POWERLED.count_offZ0Z_15_cascade_\
        );

    \I__3375\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20535\
        );

    \I__3374\ : InMux
    port map (
            O => \N__20538\,
            I => \N__20532\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__20535\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__20532\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__20527\,
            I => \POWERLED.dutycycleZ0Z_1_cascade_\
        );

    \I__3370\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20521\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__20521\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__20518\,
            I => \POWERLED.dutycycle_eena_cascade_\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__20515\,
            I => \N__20511\
        );

    \I__3366\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20508\
        );

    \I__3365\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20505\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__20508\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__20505\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__20500\,
            I => \POWERLED.dutycycle_1_0_1_cascade_\
        );

    \I__3361\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20494\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__20494\,
            I => \POWERLED.dutycycle_eena_0\
        );

    \I__3359\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20488\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__20488\,
            I => \POWERLED.dutycycle_1_0_1\
        );

    \I__3357\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20479\
        );

    \I__3356\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20479\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__20479\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__20476\,
            I => \POWERLED.dutycycle_eena_0_cascade_\
        );

    \I__3353\ : InMux
    port map (
            O => \N__20473\,
            I => \N__20467\
        );

    \I__3352\ : InMux
    port map (
            O => \N__20472\,
            I => \N__20467\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__20467\,
            I => \POWERLED.dutycycle_1_0_0\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__3349\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__20458\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__3347\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__3346\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20449\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__20449\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__20446\,
            I => \PCH_PWRGD.countZ0Z_14_cascade_\
        );

    \I__3343\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__20440\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__3341\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20431\
        );

    \I__3340\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20431\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__20431\,
            I => \N__20427\
        );

    \I__3338\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20424\
        );

    \I__3337\ : Span4Mux_s3_h
    port map (
            O => \N__20427\,
            I => \N__20419\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__20424\,
            I => \N__20419\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__20419\,
            I => \PCH_PWRGD_delayed_vccin_ok\
        );

    \I__3334\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__20413\,
            I => \PCH_PWRGD.N_250_0\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__20410\,
            I => \PCH_PWRGD.N_250_0_cascade_\
        );

    \I__3331\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__3330\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20401\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__20401\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__3328\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__20395\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__3326\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20386\
        );

    \I__3325\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20386\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__20386\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__20383\,
            I => \PCH_PWRGD.countZ0Z_15_cascade_\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__20380\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__20377\,
            I => \PCH_PWRGD.un2_count_1_axb_4_cascade_\
        );

    \I__3320\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__20371\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20368\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__20365\,
            I => \N__20362\
        );

    \I__3316\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20359\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__20359\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__3314\ : InMux
    port map (
            O => \N__20356\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__20353\,
            I => \N__20350\
        );

    \I__3312\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20347\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__20347\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__3310\ : InMux
    port map (
            O => \N__20344\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20338\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__20338\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__3307\ : InMux
    port map (
            O => \N__20335\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__20332\,
            I => \POWERLED.mult1_un145_sum_s_8_cascade_\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__20329\,
            I => \N__20325\
        );

    \I__3304\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20318\
        );

    \I__3303\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20318\
        );

    \I__3302\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20315\
        );

    \I__3301\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20312\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__20318\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__20315\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__20312\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__20305\,
            I => \N__20301\
        );

    \I__3296\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20293\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20293\
        );

    \I__3294\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20293\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__20293\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20287\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20284\
        );

    \I__3290\ : Span4Mux_s3_v
    port map (
            O => \N__20284\,
            I => \N__20280\
        );

    \I__3289\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20277\
        );

    \I__3288\ : Span4Mux_v
    port map (
            O => \N__20280\,
            I => \N__20274\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__20277\,
            I => \N__20271\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__20274\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__3285\ : Odrv12
    port map (
            O => \N__20271\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__3283\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20260\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__20260\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20254\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__20254\,
            I => \N__20251\
        );

    \I__3279\ : Span4Mux_h
    port map (
            O => \N__20251\,
            I => \N__20247\
        );

    \I__3278\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20244\
        );

    \I__3277\ : Sp12to4
    port map (
            O => \N__20247\,
            I => \N__20239\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20239\
        );

    \I__3275\ : Odrv12
    port map (
            O => \N__20239\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__20236\,
            I => \N__20233\
        );

    \I__3273\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20230\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__20230\,
            I => \N__20227\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__20224\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__20221\,
            I => \N__20217\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__20220\,
            I => \N__20214\
        );

    \I__3267\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20208\
        );

    \I__3266\ : InMux
    port map (
            O => \N__20214\,
            I => \N__20203\
        );

    \I__3265\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20203\
        );

    \I__3264\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20200\
        );

    \I__3263\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20197\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__20208\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__20203\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__20200\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__20197\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__3257\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20182\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__20182\,
            I => \N__20179\
        );

    \I__3255\ : Span4Mux_s1_h
    port map (
            O => \N__20179\,
            I => \N__20176\
        );

    \I__3254\ : Span4Mux_h
    port map (
            O => \N__20176\,
            I => \N__20173\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__20173\,
            I => \POWERLED.mult1_un68_sum_i_8\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__20170\,
            I => \N__20167\
        );

    \I__3251\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20163\
        );

    \I__3250\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20160\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__20163\,
            I => \N__20155\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20155\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__20155\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__20152\,
            I => \N__20149\
        );

    \I__3245\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20146\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__20146\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__3243\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20140\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__20140\,
            I => \N__20136\
        );

    \I__3241\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20133\
        );

    \I__3240\ : Sp12to4
    port map (
            O => \N__20136\,
            I => \N__20128\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20128\
        );

    \I__3238\ : Odrv12
    port map (
            O => \N__20128\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3237\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20122\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__3235\ : Odrv12
    port map (
            O => \N__20119\,
            I => \POWERLED.un85_clk_100khz_2\
        );

    \I__3234\ : InMux
    port map (
            O => \N__20116\,
            I => \N__20112\
        );

    \I__3233\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20109\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__20112\,
            I => \N__20106\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__20109\,
            I => \N__20103\
        );

    \I__3230\ : Span12Mux_s5_h
    port map (
            O => \N__20106\,
            I => \N__20100\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__20103\,
            I => \N__20097\
        );

    \I__3228\ : Odrv12
    port map (
            O => \N__20100\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__20097\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__3225\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20086\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__20086\,
            I => \N__20083\
        );

    \I__3223\ : Span4Mux_s3_v
    port map (
            O => \N__20083\,
            I => \N__20080\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__20080\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__3221\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20074\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__20074\,
            I => \N__20070\
        );

    \I__3219\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20067\
        );

    \I__3218\ : Span4Mux_v
    port map (
            O => \N__20070\,
            I => \N__20062\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__20067\,
            I => \N__20062\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__20062\,
            I => \N__20059\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__20059\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__20056\,
            I => \N__20053\
        );

    \I__3213\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20050\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__20050\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__3211\ : InMux
    port map (
            O => \N__20047\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__3210\ : InMux
    port map (
            O => \N__20044\,
            I => \N__20041\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__20041\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__3208\ : InMux
    port map (
            O => \N__20038\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__20035\,
            I => \N__20032\
        );

    \I__3206\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20029\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__3204\ : Span4Mux_v
    port map (
            O => \N__20026\,
            I => \N__20023\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__20023\,
            I => \N__20020\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__20020\,
            I => \POWERLED.g2_1\
        );

    \I__3201\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__20011\,
            I => \POWERLED.g2_5\
        );

    \I__3198\ : InMux
    port map (
            O => \N__20008\,
            I => \N__20005\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__3196\ : Span4Mux_h
    port map (
            O => \N__20002\,
            I => \N__19999\
        );

    \I__3195\ : Span4Mux_v
    port map (
            O => \N__19999\,
            I => \N__19996\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__19996\,
            I => \POWERLED.g0_4_4\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__19993\,
            I => \POWERLED.g0_4_5_cascade_\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__19990\,
            I => \N__19986\
        );

    \I__3191\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19983\
        );

    \I__3190\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19980\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19975\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__19980\,
            I => \N__19975\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__19975\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__3185\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19966\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__19963\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__3182\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19957\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__19957\,
            I => \POWERLED.g3_1_0\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__19954\,
            I => \POWERLED.g3_1_4_cascade_\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__19951\,
            I => \POWERLED.g3_1_6_cascade_\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__3177\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19938\
        );

    \I__3176\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19938\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__19943\,
            I => \N__19935\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__19938\,
            I => \N__19932\
        );

    \I__3173\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19929\
        );

    \I__3172\ : Span4Mux_h
    port map (
            O => \N__19932\,
            I => \N__19924\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19924\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__19924\,
            I => \POWERLED.un2_count_clk_17_0_a2_5\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__19921\,
            I => \N__19918\
        );

    \I__3168\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19915\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19912\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__19912\,
            I => \POWERLED.dutycycle_RNIZ0Z_15\
        );

    \I__3165\ : InMux
    port map (
            O => \N__19909\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__3163\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19900\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19897\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__19894\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_13\
        );

    \I__3159\ : InMux
    port map (
            O => \N__19891\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__3158\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19885\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__19885\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__3156\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19879\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19875\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__19878\,
            I => \N__19872\
        );

    \I__3153\ : Span4Mux_h
    port map (
            O => \N__19875\,
            I => \N__19869\
        );

    \I__3152\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19866\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__19869\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__19866\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__3149\ : InMux
    port map (
            O => \N__19861\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__19858\,
            I => \N__19853\
        );

    \I__3147\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19843\
        );

    \I__3146\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19843\
        );

    \I__3145\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19843\
        );

    \I__3144\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19843\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__19843\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__3142\ : InMux
    port map (
            O => \N__19840\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__19837\,
            I => \N__19833\
        );

    \I__3140\ : InMux
    port map (
            O => \N__19836\,
            I => \N__19825\
        );

    \I__3139\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19825\
        );

    \I__3138\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19825\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__19825\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__3136\ : InMux
    port map (
            O => \N__19822\,
            I => \bfn_6_11_0_\
        );

    \I__3135\ : InMux
    port map (
            O => \N__19819\,
            I => \POWERLED.CO2\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__19816\,
            I => \N__19813\
        );

    \I__3133\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19807\
        );

    \I__3132\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19807\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__19807\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__19804\,
            I => \N__19801\
        );

    \I__3129\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19798\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__19798\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__3127\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19791\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19788\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19791\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__19788\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__3123\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__19777\,
            I => \N__19774\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__19774\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__3118\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19764\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19761\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__19764\,
            I => \N__19758\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__19761\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__19758\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__3113\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19750\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19747\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__19747\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__3110\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__19741\,
            I => \N__19738\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__19738\,
            I => \N__19735\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__19735\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_3\
        );

    \I__3106\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19725\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__19728\,
            I => \N__19722\
        );

    \I__3103\ : Sp12to4
    port map (
            O => \N__19725\,
            I => \N__19719\
        );

    \I__3102\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19716\
        );

    \I__3101\ : Odrv12
    port map (
            O => \N__19719\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_3\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__19716\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_3\
        );

    \I__3099\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__19708\,
            I => \N__19704\
        );

    \I__3097\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19701\
        );

    \I__3096\ : Span4Mux_s3_h
    port map (
            O => \N__19704\,
            I => \N__19696\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19696\
        );

    \I__3094\ : Span4Mux_v
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__19693\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__3092\ : InMux
    port map (
            O => \N__19690\,
            I => \POWERLED.un1_dutycycle_53_cry_3_cZ0\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__3088\ : Span4Mux_v
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__19675\,
            I => \POWERLED.dutycycle_RNIZ0Z_4\
        );

    \I__3086\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19668\
        );

    \I__3085\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19665\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__19668\,
            I => \N__19662\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19659\
        );

    \I__3082\ : Span12Mux_s5_h
    port map (
            O => \N__19662\,
            I => \N__19656\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__19659\,
            I => \N__19653\
        );

    \I__3080\ : Odrv12
    port map (
            O => \N__19656\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__19653\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__3078\ : InMux
    port map (
            O => \N__19648\,
            I => \POWERLED.un1_dutycycle_53_cry_4_cZ0\
        );

    \I__3077\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19642\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__19642\,
            I => \N__19639\
        );

    \I__3075\ : Span4Mux_h
    port map (
            O => \N__19639\,
            I => \N__19636\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__19636\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_9\
        );

    \I__3073\ : InMux
    port map (
            O => \N__19633\,
            I => \N__19629\
        );

    \I__3072\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19626\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__19629\,
            I => \N__19623\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__19626\,
            I => \N__19620\
        );

    \I__3069\ : Span12Mux_s5_h
    port map (
            O => \N__19623\,
            I => \N__19617\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__19620\,
            I => \N__19614\
        );

    \I__3067\ : Odrv12
    port map (
            O => \N__19617\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__19614\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__3065\ : InMux
    port map (
            O => \N__19609\,
            I => \POWERLED.un1_dutycycle_53_cry_5_cZ0\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__19606\,
            I => \N__19603\
        );

    \I__3063\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19600\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__19597\,
            I => \N__19594\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__19594\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_10\
        );

    \I__3059\ : InMux
    port map (
            O => \N__19591\,
            I => \POWERLED.un1_dutycycle_53_cry_6\
        );

    \I__3058\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19585\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__19582\,
            I => \N__19579\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__19579\,
            I => \POWERLED.dutycycle_RNIZ0Z_11\
        );

    \I__3054\ : InMux
    port map (
            O => \N__19576\,
            I => \bfn_6_10_0_\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__19573\,
            I => \N__19570\
        );

    \I__3052\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19567\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__19567\,
            I => \N__19564\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__19564\,
            I => \N__19561\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__19561\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_12\
        );

    \I__3048\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19555\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__19555\,
            I => \N__19551\
        );

    \I__3046\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19548\
        );

    \I__3045\ : Span4Mux_s2_v
    port map (
            O => \N__19551\,
            I => \N__19543\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__19548\,
            I => \N__19543\
        );

    \I__3043\ : Span4Mux_v
    port map (
            O => \N__19543\,
            I => \N__19540\
        );

    \I__3042\ : Odrv4
    port map (
            O => \N__19540\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__3041\ : InMux
    port map (
            O => \N__19537\,
            I => \POWERLED.un1_dutycycle_53_cry_8\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19531\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__19531\,
            I => \N__19528\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__19525\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_13\
        );

    \I__3036\ : InMux
    port map (
            O => \N__19522\,
            I => \POWERLED.un1_dutycycle_53_cry_9\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__3034\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19513\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19510\
        );

    \I__3032\ : Odrv12
    port map (
            O => \N__19510\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_14\
        );

    \I__3031\ : InMux
    port map (
            O => \N__19507\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__3029\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19495\
        );

    \I__3028\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19495\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__19495\,
            I => \N__19492\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__19492\,
            I => \POWERLED.dutycycle_en_10\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__3024\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19480\
        );

    \I__3023\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19480\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19480\,
            I => \POWERLED.dutycycleZ1Z_13\
        );

    \I__3021\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__3020\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19471\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__19468\,
            I => \N__19465\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__19465\,
            I => \POWERLED.un1_dutycycle_53_50_0\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__19462\,
            I => \POWERLED.dutycycle_RNI_12Z0Z_9_cascade_\
        );

    \I__3015\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__19456\,
            I => \POWERLED.dutycycle_RNI_15Z0Z_9\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19448\
        );

    \I__3012\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19443\
        );

    \I__3011\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19443\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__19448\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_9\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__19443\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_9\
        );

    \I__3008\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19435\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__19435\,
            I => \N__19432\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__19432\,
            I => \N__19429\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__19426\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_0\
        );

    \I__3003\ : InMux
    port map (
            O => \N__19423\,
            I => \POWERLED.un1_dutycycle_53_cry_0_cZ0\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__19420\,
            I => \N__19417\
        );

    \I__3001\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19414\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__19411\,
            I => \N__19408\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__19408\,
            I => \POWERLED.dutycycle_RNIZ0Z_2\
        );

    \I__2997\ : InMux
    port map (
            O => \N__19405\,
            I => \POWERLED.un1_dutycycle_53_cry_1_cZ0\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19396\
        );

    \I__2994\ : Span4Mux_h
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__19393\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_2\
        );

    \I__2992\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19386\
        );

    \I__2991\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19383\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__19386\,
            I => \N__19380\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19377\
        );

    \I__2988\ : Span4Mux_v
    port map (
            O => \N__19380\,
            I => \N__19374\
        );

    \I__2987\ : Span12Mux_s5_h
    port map (
            O => \N__19377\,
            I => \N__19371\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__19374\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__2985\ : Odrv12
    port map (
            O => \N__19371\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19366\,
            I => \POWERLED.un1_dutycycle_53_cry_2_cZ0\
        );

    \I__2983\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19360\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__19360\,
            I => \POWERLED.un1_clk_100khz_39_and_i_0_0\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__19357\,
            I => \POWERLED.un1_clk_100khz_30_and_i_0_0_cascade_\
        );

    \I__2980\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19351\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__19351\,
            I => \POWERLED.dutycycle_RNI4J2O7Z0Z_9\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__19348\,
            I => \N__19345\
        );

    \I__2977\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19339\
        );

    \I__2976\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19339\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__19339\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__19336\,
            I => \POWERLED.dutycycle_RNI4J2O7Z0Z_9_cascade_\
        );

    \I__2973\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19327\
        );

    \I__2972\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19327\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__19327\,
            I => \POWERLED.dutycycleZ1Z_11\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__2969\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19318\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__19318\,
            I => \POWERLED.dutycycle_en_7\
        );

    \I__2967\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19310\
        );

    \I__2966\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19307\
        );

    \I__2965\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19304\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__19310\,
            I => \N__19301\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__19307\,
            I => \N__19298\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__19304\,
            I => \N__19294\
        );

    \I__2961\ : Span4Mux_v
    port map (
            O => \N__19301\,
            I => \N__19289\
        );

    \I__2960\ : Span4Mux_s3_h
    port map (
            O => \N__19298\,
            I => \N__19289\
        );

    \I__2959\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19286\
        );

    \I__2958\ : Span4Mux_h
    port map (
            O => \N__19294\,
            I => \N__19283\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__19289\,
            I => \POWERLED.un1_dutycycle_53_20_1\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__19286\,
            I => \POWERLED.un1_dutycycle_53_20_1\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__19283\,
            I => \POWERLED.un1_dutycycle_53_20_1\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__19276\,
            I => \POWERLED.un1_dutycycle_53_3_2_1_cascade_\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__19273\,
            I => \POWERLED.un1_dutycycle_53_3_2_cascade_\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__19270\,
            I => \N__19267\
        );

    \I__2951\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19261\
        );

    \I__2950\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19261\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__19261\,
            I => \POWERLED.dutycycleZ1Z_14\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__19258\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__2947\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19252\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__19252\,
            I => \POWERLED.dutycycle_RNI_13Z0Z_9\
        );

    \I__2945\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19246\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__19246\,
            I => \POWERLED.un1_dutycycle_53_2_0\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__19243\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__19240\,
            I => \POWERLED.un1_dutycycle_53_axb_11_cascade_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19233\
        );

    \I__2940\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19230\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19227\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__19230\,
            I => \N__19222\
        );

    \I__2937\ : Span4Mux_v
    port map (
            O => \N__19227\,
            I => \N__19222\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__19222\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_4\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__19219\,
            I => \POWERLED.dutycycle_en_7_cascade_\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__19216\,
            I => \N__19212\
        );

    \I__2933\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19209\
        );

    \I__2932\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19206\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__19209\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__19206\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__2929\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19195\
        );

    \I__2928\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19195\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__19195\,
            I => \POWERLED.count_off_1_10\
        );

    \I__2926\ : InMux
    port map (
            O => \N__19192\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__2925\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19185\
        );

    \I__2924\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19182\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__19185\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__19182\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__2921\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19171\
        );

    \I__2920\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19171\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__19171\,
            I => \POWERLED.count_off_1_11\
        );

    \I__2918\ : InMux
    port map (
            O => \N__19168\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__2917\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19161\
        );

    \I__2916\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19158\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__19161\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__19158\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__2913\ : InMux
    port map (
            O => \N__19153\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__2912\ : InMux
    port map (
            O => \N__19150\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__2911\ : InMux
    port map (
            O => \N__19147\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__2910\ : InMux
    port map (
            O => \N__19144\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__2909\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19137\
        );

    \I__2908\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19134\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__19137\,
            I => \POWERLED.count_off_1_12\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__19134\,
            I => \POWERLED.count_off_1_12\
        );

    \I__2905\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19126\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__19126\,
            I => \POWERLED.count_off_0_12\
        );

    \I__2903\ : InMux
    port map (
            O => \N__19123\,
            I => \POWERLED.un3_count_off_1_cry_1\
        );

    \I__2902\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19116\
        );

    \I__2901\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19113\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19110\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__19113\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__19110\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2897\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19099\
        );

    \I__2896\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19099\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__19096\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__19096\,
            I => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\
        );

    \I__2893\ : InMux
    port map (
            O => \N__19093\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__2892\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19086\
        );

    \I__2891\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19083\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__19086\,
            I => \N__19078\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__19083\,
            I => \N__19078\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__19078\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2887\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19069\
        );

    \I__2886\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19069\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__19069\,
            I => \N__19066\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__19066\,
            I => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\
        );

    \I__2883\ : InMux
    port map (
            O => \N__19063\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__2882\ : InMux
    port map (
            O => \N__19060\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__2881\ : InMux
    port map (
            O => \N__19057\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__2880\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19050\
        );

    \I__2879\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19047\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__19050\,
            I => \N__19044\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__19047\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2876\ : Odrv12
    port map (
            O => \N__19044\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2875\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19033\
        );

    \I__2874\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19033\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__19033\,
            I => \N__19030\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__19030\,
            I => \POWERLED.count_off_1_7\
        );

    \I__2871\ : InMux
    port map (
            O => \N__19027\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__2870\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19021\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__19021\,
            I => \N__19018\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__19018\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__2867\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19012\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__19012\,
            I => \N__19008\
        );

    \I__2865\ : InMux
    port map (
            O => \N__19011\,
            I => \N__19005\
        );

    \I__2864\ : Span4Mux_s3_h
    port map (
            O => \N__19008\,
            I => \N__19000\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__19005\,
            I => \N__19000\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__19000\,
            I => \POWERLED.count_off_1_8\
        );

    \I__2861\ : InMux
    port map (
            O => \N__18997\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__2860\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18991\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__18991\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__2858\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18982\
        );

    \I__2857\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18982\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__18982\,
            I => \POWERLED.count_off_1_9\
        );

    \I__2855\ : InMux
    port map (
            O => \N__18979\,
            I => \bfn_6_5_0_\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__18970\,
            I => \N__18967\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__18967\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__2850\ : InMux
    port map (
            O => \N__18964\,
            I => \bfn_6_3_0_\
        );

    \I__2849\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18957\
        );

    \I__2848\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18954\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__18957\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__18954\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__2845\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18945\
        );

    \I__2844\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18942\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__18945\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__18942\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18933\
        );

    \I__2840\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18930\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18927\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__18930\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__18927\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__2836\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18918\
        );

    \I__2835\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18915\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__18918\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__18915\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__18910\,
            I => \N__18907\
        );

    \I__2831\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18904\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__18904\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__2829\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18897\
        );

    \I__2828\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18894\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__18897\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__18894\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2825\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18885\
        );

    \I__2824\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18882\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__18885\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__18882\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__18877\,
            I => \N__18873\
        );

    \I__2820\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18870\
        );

    \I__2819\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18867\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__18870\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__18867\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2816\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18858\
        );

    \I__2815\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18855\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__18858\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__18855\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__18850\,
            I => \N__18847\
        );

    \I__2811\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__18844\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__2809\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18837\
        );

    \I__2808\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18834\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__18837\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__18834\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__2805\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18825\
        );

    \I__2804\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18822\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__18825\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__18822\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__18817\,
            I => \N__18813\
        );

    \I__2800\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18810\
        );

    \I__2799\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18807\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__18810\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__18807\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__2796\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18798\
        );

    \I__2795\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18795\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__18798\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__18795\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__18784\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__2789\ : IoInMux
    port map (
            O => \N__18781\,
            I => \N__18778\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__2787\ : Span4Mux_s1_h
    port map (
            O => \N__18775\,
            I => \N__18772\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__18772\,
            I => \N__18768\
        );

    \I__2785\ : IoInMux
    port map (
            O => \N__18771\,
            I => \N__18765\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__18768\,
            I => \N__18761\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__18765\,
            I => \N__18758\
        );

    \I__2782\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18754\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__18761\,
            I => \N__18750\
        );

    \I__2780\ : IoSpan4Mux
    port map (
            O => \N__18758\,
            I => \N__18747\
        );

    \I__2779\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18744\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__18754\,
            I => \N__18741\
        );

    \I__2777\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18738\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__18750\,
            I => \N__18731\
        );

    \I__2775\ : Span4Mux_s2_v
    port map (
            O => \N__18747\,
            I => \N__18731\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__18744\,
            I => \N__18731\
        );

    \I__2773\ : Span4Mux_s2_v
    port map (
            O => \N__18741\,
            I => \N__18726\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__18738\,
            I => \N__18726\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__18731\,
            I => pch_pwrok
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__18726\,
            I => pch_pwrok
        );

    \I__2769\ : IoInMux
    port map (
            O => \N__18721\,
            I => \N__18718\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__18718\,
            I => \N__18715\
        );

    \I__2767\ : Odrv12
    port map (
            O => \N__18715\,
            I => vccst_pwrgd
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__18712\,
            I => \POWERLED.mult1_un138_sum_s_8_cascade_\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__2763\ : Span4Mux_v
    port map (
            O => \N__18703\,
            I => \N__18700\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__18700\,
            I => \POWERLED.un85_clk_100khz_4\
        );

    \I__2761\ : InMux
    port map (
            O => \N__18697\,
            I => \N__18693\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18690\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__18693\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__18690\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18681\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18678\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__18681\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__18678\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__18673\,
            I => \N__18669\
        );

    \I__2752\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18666\
        );

    \I__2751\ : InMux
    port map (
            O => \N__18669\,
            I => \N__18663\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__18666\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__18663\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__2748\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18654\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18651\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__18654\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18651\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__2744\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18642\
        );

    \I__2743\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18639\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__18642\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__18639\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18630\
        );

    \I__2739\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18627\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__18630\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__18627\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__18622\,
            I => \N__18618\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18615\
        );

    \I__2734\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18612\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__18615\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__18612\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18603\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18606\,
            I => \N__18600\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__18603\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__18600\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__18595\,
            I => \N__18592\
        );

    \I__2726\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18589\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__18589\,
            I => \N__18586\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__18586\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__18583\,
            I => \N__18580\
        );

    \I__2722\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18577\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18574\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__18574\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__18571\,
            I => \N__18568\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18565\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18565\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__18562\,
            I => \N__18559\
        );

    \I__2715\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18556\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__18556\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__2713\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18549\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__18552\,
            I => \N__18546\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__18549\,
            I => \N__18540\
        );

    \I__2710\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18533\
        );

    \I__2709\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18533\
        );

    \I__2708\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18533\
        );

    \I__2707\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18530\
        );

    \I__2706\ : Odrv4
    port map (
            O => \N__18540\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__18533\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__18530\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__18523\,
            I => \N__18519\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18511\
        );

    \I__2701\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18511\
        );

    \I__2700\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18511\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__18511\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__2698\ : InMux
    port map (
            O => \N__18508\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__2697\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18502\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__18502\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__2695\ : InMux
    port map (
            O => \N__18499\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__18496\,
            I => \N__18493\
        );

    \I__2693\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18490\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__18490\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__2691\ : InMux
    port map (
            O => \N__18487\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__2690\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18481\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__18481\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18475\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__18475\,
            I => \N__18471\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__18474\,
            I => \N__18468\
        );

    \I__2685\ : Span4Mux_s2_v
    port map (
            O => \N__18471\,
            I => \N__18462\
        );

    \I__2684\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18457\
        );

    \I__2683\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18457\
        );

    \I__2682\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18454\
        );

    \I__2681\ : InMux
    port map (
            O => \N__18465\,
            I => \N__18451\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__18462\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__18457\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__18454\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__18451\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2676\ : InMux
    port map (
            O => \N__18442\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__18439\,
            I => \N__18435\
        );

    \I__2674\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18427\
        );

    \I__2673\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18427\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18427\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__18427\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__18424\,
            I => \N__18421\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18418\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__18418\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__2667\ : InMux
    port map (
            O => \N__18415\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18409\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__18409\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18406\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__2663\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18400\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__18400\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__2661\ : InMux
    port map (
            O => \N__18397\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__18394\,
            I => \N__18390\
        );

    \I__2659\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18382\
        );

    \I__2658\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18382\
        );

    \I__2657\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18382\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__18382\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__18379\,
            I => \N__18376\
        );

    \I__2654\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18373\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__18373\,
            I => \N__18370\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__18370\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18367\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__2650\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18361\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18358\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__18358\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18352\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18349\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__18349\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__2644\ : InMux
    port map (
            O => \N__18346\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__18343\,
            I => \N__18340\
        );

    \I__2642\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18337\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__18337\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__18334\,
            I => \N__18331\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18328\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__18328\,
            I => \N__18325\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__18325\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__2636\ : InMux
    port map (
            O => \N__18322\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__2635\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18316\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__18316\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__18313\,
            I => \N__18310\
        );

    \I__2632\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18307\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__18307\,
            I => \N__18304\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__18304\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__2629\ : InMux
    port map (
            O => \N__18301\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__18298\,
            I => \N__18295\
        );

    \I__2627\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18292\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__18292\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18286\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__18286\,
            I => \N__18283\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__18283\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__2622\ : InMux
    port map (
            O => \N__18280\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__2621\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18274\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__18274\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__2619\ : InMux
    port map (
            O => \N__18271\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__2618\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18264\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__18267\,
            I => \N__18260\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__18264\,
            I => \N__18257\
        );

    \I__2615\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18252\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18252\
        );

    \I__2613\ : Span4Mux_s2_v
    port map (
            O => \N__18257\,
            I => \N__18247\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__18252\,
            I => \N__18244\
        );

    \I__2611\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18241\
        );

    \I__2610\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18238\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__18247\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__18244\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__18241\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__18238\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2605\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18226\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__18226\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__2603\ : InMux
    port map (
            O => \N__18223\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__18220\,
            I => \N__18215\
        );

    \I__2601\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18211\
        );

    \I__2600\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18206\
        );

    \I__2599\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18206\
        );

    \I__2598\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18203\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__18211\,
            I => \N__18200\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__18206\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__18203\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__18200\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__18193\,
            I => \N__18189\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__18192\,
            I => \N__18185\
        );

    \I__2591\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18178\
        );

    \I__2590\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18178\
        );

    \I__2589\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18178\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__18178\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__2587\ : InMux
    port map (
            O => \N__18175\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__2586\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18169\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__18169\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__2584\ : InMux
    port map (
            O => \N__18166\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__2583\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18160\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__18160\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__2581\ : InMux
    port map (
            O => \N__18157\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__2580\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18151\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__18151\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__2578\ : InMux
    port map (
            O => \N__18148\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__18145\,
            I => \N__18142\
        );

    \I__2576\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18139\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__18139\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__2574\ : InMux
    port map (
            O => \N__18136\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__2573\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18130\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__18130\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__2571\ : InMux
    port map (
            O => \N__18127\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__2569\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18118\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__18118\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__2567\ : InMux
    port map (
            O => \N__18115\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \POWERLED.mult1_un61_sum_s_8_cascade_\
        );

    \I__2565\ : InMux
    port map (
            O => \N__18109\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18103\
        );

    \I__2563\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18100\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__18100\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__2561\ : InMux
    port map (
            O => \N__18097\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__2560\ : InMux
    port map (
            O => \N__18094\,
            I => \N__18091\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__18091\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__2558\ : InMux
    port map (
            O => \N__18088\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__2557\ : InMux
    port map (
            O => \N__18085\,
            I => \N__18082\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__18082\,
            I => \N__18079\
        );

    \I__2555\ : Span4Mux_s2_v
    port map (
            O => \N__18079\,
            I => \N__18075\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__18078\,
            I => \N__18071\
        );

    \I__2553\ : Span4Mux_h
    port map (
            O => \N__18075\,
            I => \N__18067\
        );

    \I__2552\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18062\
        );

    \I__2551\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18062\
        );

    \I__2550\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18059\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__18067\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__18062\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__18059\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__18052\,
            I => \N__18049\
        );

    \I__2545\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18046\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__18046\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__2543\ : InMux
    port map (
            O => \N__18043\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__2542\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18037\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__18037\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__18034\,
            I => \N__18030\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__18033\,
            I => \N__18026\
        );

    \I__2538\ : InMux
    port map (
            O => \N__18030\,
            I => \N__18019\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18019\
        );

    \I__2536\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18019\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__18019\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__2534\ : InMux
    port map (
            O => \N__18016\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__18013\,
            I => \N__18010\
        );

    \I__2532\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__18007\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__2530\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17999\
        );

    \I__2529\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17996\
        );

    \I__2528\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17993\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__17999\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__17996\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__17993\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__17986\,
            I => \N__17983\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17980\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__17980\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__17977\,
            I => \N__17974\
        );

    \I__2520\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17971\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__17971\,
            I => \POWERLED.mult1_un47_sum_s_4_sf\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__2517\ : InMux
    port map (
            O => \N__17965\,
            I => \N__17962\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__17962\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__2515\ : InMux
    port map (
            O => \N__17959\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__17956\,
            I => \N__17953\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17950\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__17950\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__2511\ : InMux
    port map (
            O => \N__17947\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__2510\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17941\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__17941\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__2508\ : InMux
    port map (
            O => \N__17938\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__17935\,
            I => \N__17932\
        );

    \I__2506\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17929\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__17929\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__2504\ : InMux
    port map (
            O => \N__17926\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__17923\,
            I => \N__17920\
        );

    \I__2502\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17917\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__17917\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__2500\ : InMux
    port map (
            O => \N__17914\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__2499\ : InMux
    port map (
            O => \N__17911\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__2498\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17904\
        );

    \I__2497\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17901\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__17904\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__17901\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__17896\,
            I => \N__17893\
        );

    \I__2493\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17890\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__17890\,
            I => \POWERLED.un1_dutycycle_53_4_3\
        );

    \I__2491\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17884\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__17884\,
            I => \N__17879\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__17883\,
            I => \N__17876\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__17882\,
            I => \N__17873\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__17879\,
            I => \N__17869\
        );

    \I__2486\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17862\
        );

    \I__2485\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17862\
        );

    \I__2484\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17862\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__17869\,
            I => \N__17857\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N__17857\
        );

    \I__2481\ : Span4Mux_s1_h
    port map (
            O => \N__17857\,
            I => \N__17854\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__17854\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__17851\,
            I => \N__17848\
        );

    \I__2478\ : InMux
    port map (
            O => \N__17848\,
            I => \N__17845\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__17845\,
            I => \N__17840\
        );

    \I__2476\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17836\
        );

    \I__2475\ : InMux
    port map (
            O => \N__17843\,
            I => \N__17833\
        );

    \I__2474\ : Span4Mux_h
    port map (
            O => \N__17840\,
            I => \N__17830\
        );

    \I__2473\ : InMux
    port map (
            O => \N__17839\,
            I => \N__17827\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__17836\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__17833\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__17830\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__17827\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__2468\ : InMux
    port map (
            O => \N__17818\,
            I => \N__17815\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17808\
        );

    \I__2466\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17803\
        );

    \I__2465\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17803\
        );

    \I__2464\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17798\
        );

    \I__2463\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17798\
        );

    \I__2462\ : Span4Mux_h
    port map (
            O => \N__17808\,
            I => \N__17795\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__17803\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__17798\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__17795\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__2458\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17785\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17782\
        );

    \I__2456\ : Span12Mux_s6_v
    port map (
            O => \N__17782\,
            I => \N__17779\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__17779\,
            I => \POWERLED.curr_state_1_0\
        );

    \I__2454\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17773\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__17773\,
            I => \N__17770\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__17770\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_10\
        );

    \I__2451\ : InMux
    port map (
            O => \N__17767\,
            I => \N__17764\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__17764\,
            I => \N__17761\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__17761\,
            I => \POWERLED.dutycycle_RNI_9Z0Z_9\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__17758\,
            I => \N__17755\
        );

    \I__2447\ : InMux
    port map (
            O => \N__17755\,
            I => \N__17751\
        );

    \I__2446\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17748\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__17751\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__17748\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__17743\,
            I => \POWERLED.dutycycle_en_12_cascade_\
        );

    \I__2442\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17737\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__17737\,
            I => \POWERLED.un1_clk_100khz_48_and_i_i_a3_0_0\
        );

    \I__2440\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17731\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__17731\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__17728\,
            I => \N__17724\
        );

    \I__2437\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17719\
        );

    \I__2436\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17719\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__17719\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__17716\,
            I => \POWERLED.dutycycleZ0Z_13_cascade_\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__17713\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__17710\,
            I => \POWERLED.un1_dutycycle_53_axb_12_cascade_\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__17707\,
            I => \N__17704\
        );

    \I__2430\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17697\
        );

    \I__2429\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17697\
        );

    \I__2428\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17694\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__17697\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__17694\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__2425\ : InMux
    port map (
            O => \N__17689\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__17686\,
            I => \N__17683\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17680\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__17680\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17677\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__17674\,
            I => \POWERLED.dutycycle_eena_5_cascade_\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__17671\,
            I => \POWERLED.dutycycleZ1Z_5_cascade_\
        );

    \I__2418\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17665\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__17665\,
            I => \POWERLED.dutycycle_eena_5_1\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__17662\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__17659\,
            I => \POWERLED.dutycycle_eena_6_1_cascade_\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17656\,
            I => \N__17653\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__17653\,
            I => \POWERLED.dutycycle_eena_6\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__17650\,
            I => \POWERLED.dutycycle_eena_6_cascade_\
        );

    \I__2411\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17643\
        );

    \I__2410\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17640\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__17643\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__17640\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__2407\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17632\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__17632\,
            I => \POWERLED.dutycycle_eena_5\
        );

    \I__2405\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17623\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17623\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__17623\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__17620\,
            I => \POWERLED.N_4_0_cascade_\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__17617\,
            I => \POWERLED.dutycycle_eena_8_1_cascade_\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__17614\,
            I => \POWERLED.dutycycle_eena_8_cascade_\
        );

    \I__2399\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17608\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__17608\,
            I => \POWERLED.dutycycle_eena_8\
        );

    \I__2397\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17599\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17599\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__17599\,
            I => \POWERLED.dutycycleZ1Z_3\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__17596\,
            I => \POWERLED.dutycycleZ0Z_6_cascade_\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__17593\,
            I => \POWERLED.dutycycle_eena_4_1_cascade_\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__2391\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__17584\,
            I => \POWERLED.dutycycle_eena_4\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__17581\,
            I => \POWERLED.dutycycle_eena_4_cascade_\
        );

    \I__2388\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17572\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17572\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__17572\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__2385\ : InMux
    port map (
            O => \N__17569\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__17566\,
            I => \N__17563\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__2382\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17557\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__17557\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2380\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17548\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17548\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__17548\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__17545\,
            I => \N__17541\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__17544\,
            I => \N__17538\
        );

    \I__2375\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17533\
        );

    \I__2374\ : InMux
    port map (
            O => \N__17538\,
            I => \N__17533\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__17533\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__17530\,
            I => \N__17527\
        );

    \I__2371\ : InMux
    port map (
            O => \N__17527\,
            I => \N__17521\
        );

    \I__2370\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17521\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__17521\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2368\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17515\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__17515\,
            I => \POWERLED.count_off_0_9\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__17512\,
            I => \POWERLED.count_offZ0Z_9_cascade_\
        );

    \I__2365\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17506\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__17506\,
            I => \POWERLED.count_off_0_10\
        );

    \I__2363\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17500\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__17500\,
            I => \POWERLED.count_off_0_11\
        );

    \I__2361\ : InMux
    port map (
            O => \N__17497\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__2360\ : InMux
    port map (
            O => \N__17494\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__2359\ : InMux
    port map (
            O => \N__17491\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__2358\ : InMux
    port map (
            O => \N__17488\,
            I => \bfn_5_4_0_\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17485\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17482\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__2355\ : InMux
    port map (
            O => \N__17479\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__2354\ : InMux
    port map (
            O => \N__17476\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__2353\ : InMux
    port map (
            O => \N__17473\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__2352\ : InMux
    port map (
            O => \N__17470\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__2351\ : InMux
    port map (
            O => \N__17467\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__2350\ : InMux
    port map (
            O => \N__17464\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__2349\ : InMux
    port map (
            O => \N__17461\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__2348\ : InMux
    port map (
            O => \N__17458\,
            I => \bfn_5_3_0_\
        );

    \I__2347\ : InMux
    port map (
            O => \N__17455\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__2346\ : InMux
    port map (
            O => \N__17452\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__2345\ : InMux
    port map (
            O => \N__17449\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__2344\ : InMux
    port map (
            O => \N__17446\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17443\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__17440\,
            I => \N__17435\
        );

    \I__2341\ : InMux
    port map (
            O => \N__17439\,
            I => \N__17432\
        );

    \I__2340\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17429\
        );

    \I__2339\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17426\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__17432\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__17429\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__17426\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2335\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17416\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__17416\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17413\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__2332\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17405\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17400\
        );

    \I__2330\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17400\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__17405\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__17400\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__17395\,
            I => \N__17392\
        );

    \I__2326\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17389\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__17389\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__2324\ : InMux
    port map (
            O => \N__17386\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__2323\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17379\
        );

    \I__2322\ : InMux
    port map (
            O => \N__17382\,
            I => \N__17376\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__17379\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__17376\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__2319\ : InMux
    port map (
            O => \N__17371\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__2318\ : InMux
    port map (
            O => \N__17368\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__2317\ : InMux
    port map (
            O => \N__17365\,
            I => \bfn_5_2_0_\
        );

    \I__2316\ : InMux
    port map (
            O => \N__17362\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__2315\ : InMux
    port map (
            O => \N__17359\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__2314\ : InMux
    port map (
            O => \N__17356\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17353\,
            I => \N__17350\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__17350\,
            I => \N__17347\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__17347\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__2310\ : InMux
    port map (
            O => \N__17344\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__17341\,
            I => \N__17338\
        );

    \I__2308\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17335\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__17335\,
            I => \N__17332\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__17332\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__2305\ : InMux
    port map (
            O => \N__17329\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__17326\,
            I => \N__17323\
        );

    \I__2303\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17320\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__17320\,
            I => \N__17317\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__17317\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__2300\ : InMux
    port map (
            O => \N__17314\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__2299\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17306\
        );

    \I__2298\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17301\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17301\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__17306\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__17301\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17293\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__17293\,
            I => \N__17290\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__17290\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__2291\ : InMux
    port map (
            O => \N__17287\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__2290\ : InMux
    port map (
            O => \N__17284\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__2289\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17276\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__17280\,
            I => \N__17272\
        );

    \I__2287\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17269\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__17276\,
            I => \N__17266\
        );

    \I__2285\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17261\
        );

    \I__2284\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17261\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17257\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__17266\,
            I => \N__17252\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__17261\,
            I => \N__17252\
        );

    \I__2280\ : InMux
    port map (
            O => \N__17260\,
            I => \N__17249\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__17257\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__17252\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__17249\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2276\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17237\
        );

    \I__2275\ : InMux
    port map (
            O => \N__17241\,
            I => \N__17232\
        );

    \I__2274\ : InMux
    port map (
            O => \N__17240\,
            I => \N__17232\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__17237\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__17232\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__17227\,
            I => \N__17224\
        );

    \I__2270\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17220\
        );

    \I__2269\ : InMux
    port map (
            O => \N__17223\,
            I => \N__17216\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__17220\,
            I => \N__17213\
        );

    \I__2267\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17209\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__17216\,
            I => \N__17204\
        );

    \I__2265\ : Span4Mux_s0_v
    port map (
            O => \N__17213\,
            I => \N__17204\
        );

    \I__2264\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17201\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__17209\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__17204\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__17201\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2260\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17189\
        );

    \I__2259\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17184\
        );

    \I__2258\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17184\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__17189\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__17184\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2255\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17176\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__17176\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__2253\ : InMux
    port map (
            O => \N__17173\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__2252\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17165\
        );

    \I__2251\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17160\
        );

    \I__2250\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17160\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__17165\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__17160\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2247\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17152\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__17152\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__2245\ : InMux
    port map (
            O => \N__17149\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__17146\,
            I => \N__17141\
        );

    \I__2243\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17138\
        );

    \I__2242\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17135\
        );

    \I__2241\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17132\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__17138\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__17135\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__17132\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2237\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__17122\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__2235\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__17116\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__2233\ : InMux
    port map (
            O => \N__17113\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__2231\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17094\
        );

    \I__2230\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17094\
        );

    \I__2229\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17094\
        );

    \I__2228\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17087\
        );

    \I__2227\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17087\
        );

    \I__2226\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17087\
        );

    \I__2225\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17084\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__17094\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__17087\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__17084\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2221\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__17074\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__2219\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17068\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17065\
        );

    \I__2217\ : Span4Mux_s3_v
    port map (
            O => \N__17065\,
            I => \N__17062\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__17062\,
            I => vpp_ok
        );

    \I__2215\ : IoInMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__2213\ : IoSpan4Mux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__17050\,
            I => vddq_en
        );

    \I__2211\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17044\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__17044\,
            I => \N__17041\
        );

    \I__2209\ : Span4Mux_s3_h
    port map (
            O => \N__17041\,
            I => \N__17038\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__17038\,
            I => \POWERLED.mult1_un75_sum_i_8\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__17035\,
            I => \N__17032\
        );

    \I__2206\ : InMux
    port map (
            O => \N__17032\,
            I => \N__17029\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__17029\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__2204\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17023\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__17023\,
            I => \N__17020\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__17020\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__2201\ : InMux
    port map (
            O => \N__17017\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__2200\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17011\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__17011\,
            I => \N__17008\
        );

    \I__2198\ : Odrv12
    port map (
            O => \N__17008\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__2197\ : InMux
    port map (
            O => \N__17005\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__17002\,
            I => \N__16998\
        );

    \I__2195\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16990\
        );

    \I__2194\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16990\
        );

    \I__2193\ : InMux
    port map (
            O => \N__16997\,
            I => \N__16990\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__16990\,
            I => \N__16986\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16983\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__16986\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__16983\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__16978\,
            I => \N__16974\
        );

    \I__2187\ : InMux
    port map (
            O => \N__16977\,
            I => \N__16966\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16966\
        );

    \I__2185\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16966\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__16966\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__16963\,
            I => \N__16960\
        );

    \I__2182\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16957\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__16957\,
            I => \N__16954\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__16954\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__2179\ : InMux
    port map (
            O => \N__16951\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__2178\ : InMux
    port map (
            O => \N__16948\,
            I => \N__16945\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__16945\,
            I => \N__16942\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__16942\,
            I => \POWERLED.mult1_un131_sum_axb_4_l_fx\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__16939\,
            I => \N__16936\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16932\
        );

    \I__2173\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16929\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__16932\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__16929\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__2170\ : InMux
    port map (
            O => \N__16924\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__16921\,
            I => \N__16918\
        );

    \I__2168\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16915\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__16915\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16912\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__2165\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16906\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__16906\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16903\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__2162\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16897\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__16897\,
            I => \N__16894\
        );

    \I__2160\ : Odrv12
    port map (
            O => \N__16894\,
            I => \POWERLED.mult1_un131_sum_axb_7_l_fx\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__16891\,
            I => \N__16888\
        );

    \I__2158\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16884\
        );

    \I__2157\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16881\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__16884\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__16881\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__2154\ : InMux
    port map (
            O => \N__16876\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__2153\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16870\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__16870\,
            I => \N__16867\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__16867\,
            I => \N__16864\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__16864\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__16861\,
            I => \N__16858\
        );

    \I__2148\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16855\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__16855\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__2146\ : InMux
    port map (
            O => \N__16852\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__2145\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16846\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__16846\,
            I => \N__16843\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__16843\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__2142\ : InMux
    port map (
            O => \N__16840\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16834\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__16834\,
            I => \N__16831\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__16831\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__2138\ : InMux
    port map (
            O => \N__16828\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__16825\,
            I => \N__16822\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16819\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__16819\,
            I => \N__16816\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__16816\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__2133\ : InMux
    port map (
            O => \N__16813\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__16810\,
            I => \N__16807\
        );

    \I__2131\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16804\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__16804\,
            I => \N__16801\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__16801\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__2128\ : InMux
    port map (
            O => \N__16798\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__2127\ : IoInMux
    port map (
            O => \N__16795\,
            I => \N__16792\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__16792\,
            I => \N__16788\
        );

    \I__2125\ : IoInMux
    port map (
            O => \N__16791\,
            I => \N__16785\
        );

    \I__2124\ : Span4Mux_s3_h
    port map (
            O => \N__16788\,
            I => \N__16782\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__16785\,
            I => \N__16779\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__16782\,
            I => v5s_enn
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__16779\,
            I => v5s_enn
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__16774\,
            I => \N__16771\
        );

    \I__2119\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16768\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__16768\,
            I => \POWERLED.mult1_un47_sum_i\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16762\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16759\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__16759\,
            I => \N__16756\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__16756\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__2113\ : IoInMux
    port map (
            O => \N__16753\,
            I => \N__16750\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__16750\,
            I => \N__16747\
        );

    \I__2111\ : Span4Mux_s3_h
    port map (
            O => \N__16747\,
            I => \N__16744\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__16744\,
            I => v33a_enn
        );

    \I__2109\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16738\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16735\
        );

    \I__2107\ : Span4Mux_s3_h
    port map (
            O => \N__16735\,
            I => \N__16732\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__16732\,
            I => \POWERLED.un85_clk_100khz_6\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__16729\,
            I => \POWERLED.un2_count_clk_17_0_a2_1_cascade_\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__16726\,
            I => \POWERLED.un2_count_clk_17_0_a2_5_cascade_\
        );

    \I__2103\ : InMux
    port map (
            O => \N__16723\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__2102\ : InMux
    port map (
            O => \N__16720\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__2101\ : InMux
    port map (
            O => \N__16717\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__2100\ : InMux
    port map (
            O => \N__16714\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__2099\ : InMux
    port map (
            O => \N__16711\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__2098\ : InMux
    port map (
            O => \N__16708\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__2097\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16702\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__16702\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__16699\,
            I => \POWERLED.dutycycle_eena_3_1_cascade_\
        );

    \I__2094\ : InMux
    port map (
            O => \N__16696\,
            I => \N__16693\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__16693\,
            I => \POWERLED.dutycycle_eena_3\
        );

    \I__2092\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16684\
        );

    \I__2091\ : InMux
    port map (
            O => \N__16689\,
            I => \N__16684\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__16681\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__16678\,
            I => \POWERLED.dutycycle_eena_3_cascade_\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__16675\,
            I => \POWERLED.dutycycleZ0Z_2_cascade_\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__16672\,
            I => \POWERLED.un1_dutycycle_53_4_0_cascade_\
        );

    \I__2085\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16666\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__16666\,
            I => \POWERLED.un1_dutycycle_53_4_3_1\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__16663\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_12_cascade_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16657\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__16657\,
            I => \POWERLED.un1_dutycycle_53_8_3\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__16654\,
            I => \N__16650\
        );

    \I__2079\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16647\
        );

    \I__2078\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16644\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__16647\,
            I => \N__16641\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__16644\,
            I => \N__16636\
        );

    \I__2075\ : Span4Mux_h
    port map (
            O => \N__16641\,
            I => \N__16633\
        );

    \I__2074\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16628\
        );

    \I__2073\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16628\
        );

    \I__2072\ : Span12Mux_s3_h
    port map (
            O => \N__16636\,
            I => \N__16625\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__16633\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__16628\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__16625\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3\
        );

    \I__2068\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16615\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__16615\,
            I => \POWERLED.un1_dutycycle_53_56_a0_1\
        );

    \I__2066\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16609\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__16609\,
            I => \POWERLED.un1_dutycycle_53_56_a1_1\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__16606\,
            I => \POWERLED.un1_clk_100khz_45_and_i_i_a3_0_0_cascade_\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__16603\,
            I => \POWERLED.N_4_cascade_\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__16600\,
            I => \POWERLED.un1_dutycycle_53_axb_7_cascade_\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__16597\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16591\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__16591\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_10\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__16588\,
            I => \POWERLED.un1_dutycycle_53_axb_4_1_cascade_\
        );

    \I__2057\ : InMux
    port map (
            O => \N__16585\,
            I => \N__16582\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__16582\,
            I => \POWERLED.un1_dutycycle_53_8_2_0\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__16579\,
            I => \POWERLED.un1_dutycycle_53_8_2_cascade_\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__16576\,
            I => \POWERLED.un1_dutycycle_53_8_5_cascade_\
        );

    \I__2053\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16570\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__16570\,
            I => \POWERLED.count_off_0_7\
        );

    \I__2051\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16563\
        );

    \I__2050\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16560\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16563\,
            I => \N__16557\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__16560\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__16557\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__2046\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16548\
        );

    \I__2045\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16545\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16542\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__16545\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__2042\ : Odrv12
    port map (
            O => \N__16542\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__16537\,
            I => \N__16534\
        );

    \I__2040\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16531\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__16531\,
            I => \N__16527\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16524\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__16527\,
            I => \N__16521\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__16524\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__16521\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__2034\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16512\
        );

    \I__2033\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16509\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__16512\,
            I => \N__16506\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__16509\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__16506\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__2029\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16498\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__16495\,
            I => \DSW_PWRGD.un4_count_8\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__16492\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_3_cascade_\
        );

    \I__2025\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16486\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16483\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__16483\,
            I => \N__16479\
        );

    \I__2022\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16476\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__16479\,
            I => \POWERLED.un1_dutycycle_53_20_0_0\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__16476\,
            I => \POWERLED.un1_dutycycle_53_20_0_0\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__16471\,
            I => \POWERLED.o2_cascade_\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__16468\,
            I => \N__16465\
        );

    \I__2017\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16462\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16462\,
            I => \POWERLED.un1_dutycycle_53_axb_7_1\
        );

    \I__2015\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16456\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__16456\,
            I => \POWERLED.count_off_0_4\
        );

    \I__2013\ : InMux
    port map (
            O => \N__16453\,
            I => \N__16450\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__16450\,
            I => \N__16447\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__16447\,
            I => \POWERLED.count_off_0_8\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__16444\,
            I => \POWERLED.count_offZ0Z_8_cascade_\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__16441\,
            I => \N__16438\
        );

    \I__2008\ : InMux
    port map (
            O => \N__16438\,
            I => \N__16435\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__16435\,
            I => \POWERLED.count_off_0_3\
        );

    \I__2006\ : InMux
    port map (
            O => \N__16432\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__16429\,
            I => \N__16425\
        );

    \I__2004\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16420\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16415\
        );

    \I__2002\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16415\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16412\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__16420\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__16415\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__16412\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__16405\,
            I => \POWERLED.mult1_un96_sum_s_8_cascade_\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \N__16398\
        );

    \I__1995\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16390\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16390\
        );

    \I__1993\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16390\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__16390\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__1991\ : InMux
    port map (
            O => \N__16387\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__16384\,
            I => \N__16380\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__16383\,
            I => \N__16377\
        );

    \I__1988\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16372\
        );

    \I__1987\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16369\
        );

    \I__1986\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16366\
        );

    \I__1985\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16363\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__16372\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__16369\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__16366\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__16363\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__16354\,
            I => \POWERLED.mult1_un103_sum_s_8_cascade_\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__16351\,
            I => \N__16347\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__16350\,
            I => \N__16343\
        );

    \I__1977\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16336\
        );

    \I__1976\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16336\
        );

    \I__1975\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16336\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__16336\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16333\,
            I => \N__16330\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__16330\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__1971\ : InMux
    port map (
            O => \N__16327\,
            I => \POWERLED.mult1_un96_sum_cry_2_c\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__16324\,
            I => \N__16321\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16318\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__16318\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__1967\ : InMux
    port map (
            O => \N__16315\,
            I => \POWERLED.mult1_un96_sum_cry_3_c\
        );

    \I__1966\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16309\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__16309\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16306\,
            I => \POWERLED.mult1_un96_sum_cry_4_c\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__16303\,
            I => \N__16300\
        );

    \I__1962\ : InMux
    port map (
            O => \N__16300\,
            I => \N__16297\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__16297\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__1960\ : InMux
    port map (
            O => \N__16294\,
            I => \POWERLED.mult1_un96_sum_cry_5_c\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__16291\,
            I => \N__16288\
        );

    \I__1958\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16279\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16279\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16279\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__16279\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__1954\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16273\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__16273\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__1952\ : InMux
    port map (
            O => \N__16270\,
            I => \POWERLED.mult1_un96_sum_cry_6_c\
        );

    \I__1951\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16264\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__16264\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__1949\ : InMux
    port map (
            O => \N__16261\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__1948\ : InMux
    port map (
            O => \N__16258\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__1947\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16250\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__16254\,
            I => \N__16247\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__16253\,
            I => \N__16244\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__16250\,
            I => \N__16239\
        );

    \I__1943\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16236\
        );

    \I__1942\ : InMux
    port map (
            O => \N__16244\,
            I => \N__16233\
        );

    \I__1941\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16230\
        );

    \I__1940\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16227\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__16239\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__16236\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__16233\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__16230\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__16227\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__16216\,
            I => \N__16211\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__16215\,
            I => \N__16208\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__16214\,
            I => \N__16205\
        );

    \I__1931\ : InMux
    port map (
            O => \N__16211\,
            I => \N__16202\
        );

    \I__1930\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16197\
        );

    \I__1929\ : InMux
    port map (
            O => \N__16205\,
            I => \N__16197\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__16202\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__16197\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__16192\,
            I => \N__16189\
        );

    \I__1925\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16186\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__16186\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__1923\ : InMux
    port map (
            O => \N__16183\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__1922\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16177\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__16177\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__1920\ : InMux
    port map (
            O => \N__16174\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__1919\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16168\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__16168\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__1917\ : InMux
    port map (
            O => \N__16165\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__1916\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16159\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__16159\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__1914\ : InMux
    port map (
            O => \N__16156\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__1913\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16150\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__16150\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__1911\ : InMux
    port map (
            O => \N__16147\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__1910\ : InMux
    port map (
            O => \N__16144\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__1909\ : InMux
    port map (
            O => \N__16141\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__1908\ : InMux
    port map (
            O => \N__16138\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__16135\,
            I => \POWERLED.mult1_un117_sum_s_8_cascade_\
        );

    \I__1906\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16129\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__16129\,
            I => \POWERLED.un85_clk_100khz_7\
        );

    \I__1904\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16123\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__16123\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__1902\ : InMux
    port map (
            O => \N__16120\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__1901\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16114\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__16114\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__1899\ : InMux
    port map (
            O => \N__16111\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__1898\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16105\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__16105\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__1896\ : InMux
    port map (
            O => \N__16102\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__1895\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16096\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__16096\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__1893\ : InMux
    port map (
            O => \N__16093\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \N__16087\
        );

    \I__1891\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16081\
        );

    \I__1890\ : InMux
    port map (
            O => \N__16086\,
            I => \N__16081\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__16081\,
            I => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\
        );

    \I__1888\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16075\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__16075\,
            I => \POWERLED.count_0_15\
        );

    \I__1886\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16068\
        );

    \I__1885\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16064\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__16068\,
            I => \N__16061\
        );

    \I__1883\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16058\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__16064\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__16061\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__16058\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__16051\,
            I => \N__16048\
        );

    \I__1878\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16042\
        );

    \I__1877\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16042\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__16042\,
            I => \N__16039\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__16039\,
            I => \POWERLED.count_1_7\
        );

    \I__1874\ : InMux
    port map (
            O => \N__16036\,
            I => \N__16033\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__16033\,
            I => \POWERLED.count_0_7\
        );

    \I__1872\ : InMux
    port map (
            O => \N__16030\,
            I => \N__16027\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__16027\,
            I => \N__16023\
        );

    \I__1870\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16020\
        );

    \I__1869\ : Span4Mux_s3_v
    port map (
            O => \N__16023\,
            I => \N__16014\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__16020\,
            I => \N__16014\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16019\,
            I => \N__16011\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__16014\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__16011\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__16006\,
            I => \N__16002\
        );

    \I__1863\ : InMux
    port map (
            O => \N__16005\,
            I => \N__15997\
        );

    \I__1862\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15997\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__15997\,
            I => \N__15994\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__15994\,
            I => \POWERLED.count_1_8\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15988\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__15988\,
            I => \POWERLED.count_0_8\
        );

    \I__1857\ : InMux
    port map (
            O => \N__15985\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__1856\ : InMux
    port map (
            O => \N__15982\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__1855\ : InMux
    port map (
            O => \N__15979\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__1854\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15971\
        );

    \I__1853\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15968\
        );

    \I__1852\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15965\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15960\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15968\,
            I => \N__15960\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__15965\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1848\ : Odrv12
    port map (
            O => \N__15960\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1847\ : InMux
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__1846\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15949\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__15949\,
            I => \POWERLED.count_1_12\
        );

    \I__1844\ : InMux
    port map (
            O => \N__15946\,
            I => \POWERLED.un1_count_cry_11_cZ0\
        );

    \I__1843\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15938\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__15942\,
            I => \N__15935\
        );

    \I__1841\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15932\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__15938\,
            I => \N__15929\
        );

    \I__1839\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15926\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__15932\,
            I => \N__15923\
        );

    \I__1837\ : Sp12to4
    port map (
            O => \N__15929\,
            I => \N__15918\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15926\,
            I => \N__15918\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__15923\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1834\ : Odrv12
    port map (
            O => \N__15918\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__1832\ : InMux
    port map (
            O => \N__15912\,
            I => \N__15907\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__15907\,
            I => \N__15904\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__15904\,
            I => \POWERLED.count_1_13\
        );

    \I__1829\ : InMux
    port map (
            O => \N__15901\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__1828\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15894\
        );

    \I__1827\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15890\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__15894\,
            I => \N__15887\
        );

    \I__1825\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15884\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15881\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__15887\,
            I => \N__15876\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15876\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__15881\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__15876\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1819\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15865\
        );

    \I__1818\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15865\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__15865\,
            I => \N__15862\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__15862\,
            I => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\
        );

    \I__1815\ : InMux
    port map (
            O => \N__15859\,
            I => \POWERLED.un1_count_cry_13_cZ0\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__15856\,
            I => \N__15852\
        );

    \I__1813\ : InMux
    port map (
            O => \N__15855\,
            I => \N__15830\
        );

    \I__1812\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15830\
        );

    \I__1811\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15830\
        );

    \I__1810\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15821\
        );

    \I__1809\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15821\
        );

    \I__1808\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15821\
        );

    \I__1807\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15821\
        );

    \I__1806\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15814\
        );

    \I__1805\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15814\
        );

    \I__1804\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15814\
        );

    \I__1803\ : InMux
    port map (
            O => \N__15843\,
            I => \N__15807\
        );

    \I__1802\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15807\
        );

    \I__1801\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15807\
        );

    \I__1800\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15798\
        );

    \I__1799\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15798\
        );

    \I__1798\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15798\
        );

    \I__1797\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15798\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__15830\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__15821\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__15814\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__15807\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__15798\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__1791\ : InMux
    port map (
            O => \N__15787\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15781\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15781\,
            I => \N__15778\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__15778\,
            I => \N__15775\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__15775\,
            I => \POWERLED.count_0_9\
        );

    \I__1786\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15769\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__15769\,
            I => \N__15765\
        );

    \I__1784\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15762\
        );

    \I__1783\ : Odrv4
    port map (
            O => \N__15765\,
            I => \POWERLED.count_1_9\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__15762\,
            I => \POWERLED.count_1_9\
        );

    \I__1781\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15754\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15749\
        );

    \I__1779\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15746\
        );

    \I__1778\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15743\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__15749\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__15746\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__15743\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15732\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15728\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__15732\,
            I => \N__15725\
        );

    \I__1771\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15722\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__15728\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__15725\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__15722\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15712\
        );

    \I__1766\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15706\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15706\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__15706\,
            I => \N__15703\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__15703\,
            I => \POWERLED.count_1_6\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15700\,
            I => \N__15697\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15697\,
            I => \POWERLED.count_0_6\
        );

    \I__1760\ : InMux
    port map (
            O => \N__15694\,
            I => \N__15691\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__15691\,
            I => \N__15688\
        );

    \I__1758\ : Span12Mux_s1_h
    port map (
            O => \N__15688\,
            I => \N__15683\
        );

    \I__1757\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15680\
        );

    \I__1756\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15677\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__15683\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__15680\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__15677\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1752\ : InMux
    port map (
            O => \N__15670\,
            I => \N__15665\
        );

    \I__1751\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15662\
        );

    \I__1750\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15659\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__15665\,
            I => \N__15654\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15654\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__15659\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__15654\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \N__15646\
        );

    \I__1744\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15640\
        );

    \I__1743\ : InMux
    port map (
            O => \N__15645\,
            I => \N__15640\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__15640\,
            I => \POWERLED.count_1_4\
        );

    \I__1741\ : InMux
    port map (
            O => \N__15637\,
            I => \POWERLED.un1_count_cry_3\
        );

    \I__1740\ : InMux
    port map (
            O => \N__15634\,
            I => \N__15631\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__15631\,
            I => \N__15626\
        );

    \I__1738\ : InMux
    port map (
            O => \N__15630\,
            I => \N__15623\
        );

    \I__1737\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15620\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__15626\,
            I => \N__15615\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__15623\,
            I => \N__15615\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__15620\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__15615\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__15610\,
            I => \N__15607\
        );

    \I__1731\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15601\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15601\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__15601\,
            I => \POWERLED.count_1_5\
        );

    \I__1728\ : InMux
    port map (
            O => \N__15598\,
            I => \POWERLED.un1_count_cry_4\
        );

    \I__1727\ : InMux
    port map (
            O => \N__15595\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__1726\ : InMux
    port map (
            O => \N__15592\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15589\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__1724\ : InMux
    port map (
            O => \N__15586\,
            I => \bfn_2_11_0_\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15580\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__15580\,
            I => \N__15575\
        );

    \I__1721\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15572\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15569\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__15575\,
            I => \N__15562\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__15572\,
            I => \N__15562\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__15569\,
            I => \N__15562\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__15562\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15553\
        );

    \I__1714\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15553\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__15553\,
            I => \N__15550\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__15550\,
            I => \POWERLED.count_1_10\
        );

    \I__1711\ : InMux
    port map (
            O => \N__15547\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15540\
        );

    \I__1709\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15537\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__15540\,
            I => \N__15533\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15537\,
            I => \N__15530\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15536\,
            I => \N__15527\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__15533\,
            I => \N__15520\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__15530\,
            I => \N__15520\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__15527\,
            I => \N__15520\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__15520\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1701\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15511\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15511\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__15511\,
            I => \N__15508\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__15508\,
            I => \POWERLED.count_1_11\
        );

    \I__1697\ : InMux
    port map (
            O => \N__15505\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15499\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__15499\,
            I => \POWERLED.count_0_10\
        );

    \I__1694\ : InMux
    port map (
            O => \N__15496\,
            I => \N__15493\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__15493\,
            I => \POWERLED.count_0_2\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15487\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__15487\,
            I => \POWERLED.count_0_11\
        );

    \I__1690\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15481\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__15481\,
            I => \N__15476\
        );

    \I__1688\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15473\
        );

    \I__1687\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15470\
        );

    \I__1686\ : Odrv12
    port map (
            O => \N__15476\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__15473\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__15470\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1683\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15459\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__15462\,
            I => \N__15452\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__15459\,
            I => \N__15449\
        );

    \I__1680\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15446\
        );

    \I__1679\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15439\
        );

    \I__1678\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15439\
        );

    \I__1677\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15439\
        );

    \I__1676\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15436\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__15449\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__15446\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__15439\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__15436\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15427\,
            I => \N__15424\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__15424\,
            I => \N__15419\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15416\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15413\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__15419\,
            I => \N__15408\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__15416\,
            I => \N__15408\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__15413\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__15408\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__15403\,
            I => \N__15399\
        );

    \I__1662\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15394\
        );

    \I__1661\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15394\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__15394\,
            I => \POWERLED.count_1_2\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15391\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__15388\,
            I => \N__15384\
        );

    \I__1657\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15380\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15377\
        );

    \I__1655\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15374\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__15380\,
            I => \N__15369\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__15377\,
            I => \N__15369\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__15374\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__15369\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__15364\,
            I => \N__15361\
        );

    \I__1649\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15355\
        );

    \I__1648\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15355\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__15355\,
            I => \POWERLED.count_1_3\
        );

    \I__1646\ : InMux
    port map (
            O => \N__15352\,
            I => \POWERLED.un1_count_cry_2\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__15349\,
            I => \POWERLED.dutycycle_RNIZ0Z_1_cascade_\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__15346\,
            I => \N__15343\
        );

    \I__1643\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__15340\,
            I => \POWERLED.un1_dutycycle_53_axb_3_1\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__15337\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__15334\,
            I => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \I__1639\ : SRMux
    port map (
            O => \N__15331\,
            I => \N__15327\
        );

    \I__1638\ : SRMux
    port map (
            O => \N__15330\,
            I => \N__15323\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__15327\,
            I => \N__15320\
        );

    \I__1636\ : SRMux
    port map (
            O => \N__15326\,
            I => \N__15317\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__15323\,
            I => \N__15314\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__15320\,
            I => \N__15311\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15317\,
            I => \N__15308\
        );

    \I__1632\ : Span4Mux_s2_h
    port map (
            O => \N__15314\,
            I => \N__15305\
        );

    \I__1631\ : Span4Mux_s1_h
    port map (
            O => \N__15311\,
            I => \N__15300\
        );

    \I__1630\ : Span4Mux_s1_h
    port map (
            O => \N__15308\,
            I => \N__15300\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__15305\,
            I => \G_27\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__15300\,
            I => \G_27\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__15295\,
            I => \G_27_cascade_\
        );

    \I__1626\ : CEMux
    port map (
            O => \N__15292\,
            I => \N__15289\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15286\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__15286\,
            I => \DSW_PWRGD.N_29_1\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__15283\,
            I => \POWERLED.d_i1_mux_cascade_\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__15280\,
            I => \POWERLED.dutycycle_RNI_16Z0Z_9_cascade_\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__15277\,
            I => \POWERLED.d_i3_mux_cascade_\
        );

    \I__1620\ : InMux
    port map (
            O => \N__15274\,
            I => \N__15268\
        );

    \I__1619\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15268\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__15268\,
            I => \POWERLED.un1_i3_mux\
        );

    \I__1617\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15261\
        );

    \I__1616\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__15261\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__15258\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__1613\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15249\
        );

    \I__1612\ : InMux
    port map (
            O => \N__15252\,
            I => \N__15246\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__15249\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__15246\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__15241\,
            I => \N__15237\
        );

    \I__1608\ : InMux
    port map (
            O => \N__15240\,
            I => \N__15234\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15231\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__15234\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__15231\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__1604\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15222\
        );

    \I__1603\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15219\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__15222\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__15219\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__1600\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15211\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__15211\,
            I => \DSW_PWRGD.un4_count_10\
        );

    \I__1598\ : InMux
    port map (
            O => \N__15208\,
            I => \N__15204\
        );

    \I__1597\ : InMux
    port map (
            O => \N__15207\,
            I => \N__15201\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__15204\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__15201\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__1594\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15192\
        );

    \I__1593\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15189\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__15192\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__15189\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__15184\,
            I => \N__15180\
        );

    \I__1589\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15177\
        );

    \I__1588\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15174\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__15177\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__15174\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__1585\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15165\
        );

    \I__1584\ : InMux
    port map (
            O => \N__15168\,
            I => \N__15162\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__15165\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__15162\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__1581\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15154\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__15154\,
            I => \DSW_PWRGD.un4_count_11\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__15151\,
            I => \N__15147\
        );

    \I__1578\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15144\
        );

    \I__1577\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15141\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__15144\,
            I => \DSW_PWRGD.un1_curr_state10_0\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__15141\,
            I => \DSW_PWRGD.un1_curr_state10_0\
        );

    \I__1574\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15121\
        );

    \I__1573\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15121\
        );

    \I__1572\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15121\
        );

    \I__1571\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15121\
        );

    \I__1570\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15121\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__15121\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__15118\,
            I => \N__15113\
        );

    \I__1567\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15100\
        );

    \I__1566\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15100\
        );

    \I__1565\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15100\
        );

    \I__1564\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15100\
        );

    \I__1563\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15100\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__15100\,
            I => \N__15097\
        );

    \I__1561\ : Span4Mux_v
    port map (
            O => \N__15097\,
            I => \N__15094\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__15094\,
            I => \N__15091\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__15091\,
            I => v33dsw_ok
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__15088\,
            I => \N__15082\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__15087\,
            I => \N__15079\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__15086\,
            I => \N__15076\
        );

    \I__1555\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15072\
        );

    \I__1554\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15063\
        );

    \I__1553\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15063\
        );

    \I__1552\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15063\
        );

    \I__1551\ : InMux
    port map (
            O => \N__15075\,
            I => \N__15063\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__15072\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__15063\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__1548\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15055\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__15055\,
            I => \N__15050\
        );

    \I__1546\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15045\
        );

    \I__1545\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15045\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__15050\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__15045\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__1542\ : InMux
    port map (
            O => \N__15040\,
            I => \N__15037\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__1540\ : Span12Mux_s8_h
    port map (
            O => \N__15034\,
            I => \N__15031\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__15031\,
            I => gpio_fpga_soc_1
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__15028\,
            I => \N__15024\
        );

    \I__1537\ : InMux
    port map (
            O => \N__15027\,
            I => \N__15007\
        );

    \I__1536\ : InMux
    port map (
            O => \N__15024\,
            I => \N__15007\
        );

    \I__1535\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15007\
        );

    \I__1534\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15003\
        );

    \I__1533\ : InMux
    port map (
            O => \N__15021\,
            I => \N__14992\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15020\,
            I => \N__14992\
        );

    \I__1531\ : InMux
    port map (
            O => \N__15019\,
            I => \N__14992\
        );

    \I__1530\ : InMux
    port map (
            O => \N__15018\,
            I => \N__14992\
        );

    \I__1529\ : InMux
    port map (
            O => \N__15017\,
            I => \N__14992\
        );

    \I__1528\ : InMux
    port map (
            O => \N__15016\,
            I => \N__14989\
        );

    \I__1527\ : InMux
    port map (
            O => \N__15015\,
            I => \N__14986\
        );

    \I__1526\ : InMux
    port map (
            O => \N__15014\,
            I => \N__14983\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__15007\,
            I => \N__14980\
        );

    \I__1524\ : InMux
    port map (
            O => \N__15006\,
            I => \N__14977\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15003\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__14992\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14989\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__14986\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__14983\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__14980\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__14977\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__14962\,
            I => \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_\
        );

    \I__1515\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14956\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__14956\,
            I => \HDA_STRAP.curr_state_RNO_0Z0Z_0\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__14953\,
            I => \N__14945\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__14952\,
            I => \N__14942\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__14951\,
            I => \N__14938\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__14950\,
            I => \N__14933\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__14949\,
            I => \N__14930\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__14948\,
            I => \N__14925\
        );

    \I__1507\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14918\
        );

    \I__1506\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14918\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14915\
        );

    \I__1504\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14908\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14908\
        );

    \I__1502\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14908\
        );

    \I__1501\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14900\
        );

    \I__1500\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14900\
        );

    \I__1499\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14900\
        );

    \I__1498\ : InMux
    port map (
            O => \N__14928\,
            I => \N__14891\
        );

    \I__1497\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14891\
        );

    \I__1496\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14891\
        );

    \I__1495\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14891\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__14918\,
            I => \N__14884\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__14915\,
            I => \N__14884\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__14908\,
            I => \N__14884\
        );

    \I__1491\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14881\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__14900\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__14891\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__14884\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__14881\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1486\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14869\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__14869\,
            I => \HDA_STRAP.N_5_0\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14862\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14865\,
            I => \N__14859\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__14862\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14859\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__1480\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14850\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14853\,
            I => \N__14847\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14850\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__14847\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__14842\,
            I => \N__14839\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14835\
        );

    \I__1474\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14832\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__14835\,
            I => \N__14829\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__14832\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__14829\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__1470\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14820\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14817\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__14820\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__14817\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__14812\,
            I => \DSW_PWRGD.un4_count_9_cascade_\
        );

    \I__1465\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14805\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14802\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__14805\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__14802\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__14797\,
            I => \N__14793\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14790\
        );

    \I__1459\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14787\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__14790\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__14787\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__1456\ : InMux
    port map (
            O => \N__14782\,
            I => \N__14779\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__14779\,
            I => \N__14776\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__14776\,
            I => \HDA_STRAP.un4_count_12\
        );

    \I__1453\ : InMux
    port map (
            O => \N__14773\,
            I => \N__14770\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__14770\,
            I => \HDA_STRAP.count_RNO_0Z0Z_6\
        );

    \I__1451\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14763\
        );

    \I__1450\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14760\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__14763\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__14760\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__1447\ : InMux
    port map (
            O => \N__14755\,
            I => \N__14752\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__14752\,
            I => \HDA_STRAP.count_RNO_0Z0Z_8\
        );

    \I__1445\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14745\
        );

    \I__1444\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14742\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__14745\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__14742\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__1441\ : InMux
    port map (
            O => \N__14737\,
            I => \N__14734\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__14734\,
            I => \HDA_STRAP.count_RNO_0Z0Z_11\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14727\
        );

    \I__1438\ : InMux
    port map (
            O => \N__14730\,
            I => \N__14724\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__14727\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14724\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__14719\,
            I => \HDA_STRAP.N_14_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14705\
        );

    \I__1433\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14694\
        );

    \I__1432\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14694\
        );

    \I__1431\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14694\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14712\,
            I => \N__14694\
        );

    \I__1429\ : InMux
    port map (
            O => \N__14711\,
            I => \N__14694\
        );

    \I__1428\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14687\
        );

    \I__1427\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14687\
        );

    \I__1426\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14687\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__14705\,
            I => \N__14684\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__14694\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__14687\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__14684\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1421\ : InMux
    port map (
            O => \N__14677\,
            I => \N__14673\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14676\,
            I => \N__14670\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__14673\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__14670\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1417\ : IoInMux
    port map (
            O => \N__14665\,
            I => \N__14662\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14659\
        );

    \I__1415\ : IoSpan4Mux
    port map (
            O => \N__14659\,
            I => \N__14656\
        );

    \I__1414\ : Span4Mux_s1_h
    port map (
            O => \N__14656\,
            I => \N__14653\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__14653\,
            I => hda_sdo_atp
        );

    \I__1412\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14647\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__14647\,
            I => \HDA_STRAP.count_RNO_0Z0Z_0\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__14644\,
            I => \HDA_STRAP.un4_count_cascade_\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14637\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14634\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__14637\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__14634\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14629\,
            I => \N__14625\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14622\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__14625\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__14622\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__14617\,
            I => \N__14614\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14610\
        );

    \I__1399\ : InMux
    port map (
            O => \N__14613\,
            I => \N__14607\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__14610\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__14607\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14598\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14601\,
            I => \N__14595\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__14598\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__14595\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__14587\,
            I => \HDA_STRAP.un4_count_10\
        );

    \I__1390\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14581\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__14581\,
            I => \N__14578\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__14578\,
            I => \HDA_STRAP.count_RNO_0Z0Z_17\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14571\
        );

    \I__1386\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14568\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__14571\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__14568\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__14563\,
            I => \N__14560\
        );

    \I__1382\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14557\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__1380\ : Span4Mux_s2_h
    port map (
            O => \N__14554\,
            I => \N__14550\
        );

    \I__1379\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14547\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__14550\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__14547\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1376\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14535\
        );

    \I__1374\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14532\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__14535\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__14532\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__14527\,
            I => \HDA_STRAP.un4_count_9_cascade_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__14521\,
            I => \HDA_STRAP.un4_count_13\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__1367\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__14512\,
            I => \N__14509\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__14509\,
            I => \HDA_STRAP.count_RNO_0Z0Z_16\
        );

    \I__1364\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__14503\,
            I => \N__14499\
        );

    \I__1362\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14496\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__14499\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__14496\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__1359\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14488\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__14488\,
            I => \HDA_STRAP.count_RNO_0Z0Z_10\
        );

    \I__1357\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14481\
        );

    \I__1356\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14478\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__14481\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__14478\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1353\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14469\
        );

    \I__1352\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14466\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__14469\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__14466\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14457\
        );

    \I__1348\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14454\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__14457\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__14454\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__14449\,
            I => \N__14445\
        );

    \I__1344\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14442\
        );

    \I__1343\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14439\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__14442\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__14439\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14430\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14427\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14430\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__14427\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__14422\,
            I => \N__14419\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14416\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__14416\,
            I => \HDA_STRAP.un4_count_11\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14410\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__14410\,
            I => \N__14407\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__14407\,
            I => \POWERLED.un85_clk_100khz_5\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__14404\,
            I => \N__14401\
        );

    \I__1329\ : InMux
    port map (
            O => \N__14401\,
            I => \N__14398\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__14398\,
            I => \POWERLED.un85_clk_100khz_9\
        );

    \I__1327\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__14392\,
            I => \N__14389\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__14389\,
            I => \POWERLED.un85_clk_100khz_8\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__14386\,
            I => \N__14383\
        );

    \I__1323\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14380\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__14380\,
            I => \N__14377\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__14377\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__14374\,
            I => \N__14371\
        );

    \I__1319\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14368\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__14368\,
            I => \N__14365\
        );

    \I__1317\ : Odrv4
    port map (
            O => \N__14365\,
            I => \POWERLED.un85_clk_100khz_10\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__14362\,
            I => \N__14359\
        );

    \I__1315\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14356\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14353\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__14353\,
            I => \POWERLED.mult1_un89_sum_i_8\
        );

    \I__1312\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__14347\,
            I => \N__14344\
        );

    \I__1310\ : Odrv12
    port map (
            O => \N__14344\,
            I => \POWERLED.un85_clk_100khz_3\
        );

    \I__1309\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14338\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__14338\,
            I => \POWERLED.N_5118_i\
        );

    \I__1307\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14332\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__14332\,
            I => \POWERLED.N_5119_i\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14329\,
            I => \N__14326\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__14326\,
            I => \POWERLED.N_5120_i\
        );

    \I__1303\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14320\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__14320\,
            I => \POWERLED.N_5121_i\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__14317\,
            I => \N__14314\
        );

    \I__1300\ : InMux
    port map (
            O => \N__14314\,
            I => \N__14311\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__14308\,
            I => \POWERLED.N_5122_i\
        );

    \I__1297\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14302\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__14302\,
            I => \POWERLED.N_5123_i\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14296\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__14296\,
            I => \POWERLED.N_5124_i\
        );

    \I__1293\ : InMux
    port map (
            O => \N__14293\,
            I => \bfn_1_15_0_\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__14290\,
            I => \N__14287\
        );

    \I__1291\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14284\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14281\
        );

    \I__1289\ : Odrv12
    port map (
            O => \N__14281\,
            I => \POWERLED.mult1_un82_sum_i_8\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__1287\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14272\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__14272\,
            I => \POWERLED.N_5110_i\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__1284\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14263\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14260\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__14260\,
            I => \POWERLED.N_5111_i\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__14257\,
            I => \N__14254\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14251\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14248\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__14248\,
            I => \POWERLED.N_5112_i\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__14245\,
            I => \N__14242\
        );

    \I__1276\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14239\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__14239\,
            I => \POWERLED.N_5113_i\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__14236\,
            I => \N__14233\
        );

    \I__1273\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__14230\,
            I => \POWERLED.N_5114_i\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__14227\,
            I => \N__14224\
        );

    \I__1270\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14221\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__14221\,
            I => \POWERLED.N_5115_i\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \N__14215\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14212\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__14212\,
            I => \N__14209\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__14209\,
            I => \POWERLED.N_5116_i\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__14206\,
            I => \N__14203\
        );

    \I__1263\ : InMux
    port map (
            O => \N__14203\,
            I => \N__14200\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__14200\,
            I => \POWERLED.N_5117_i\
        );

    \I__1261\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14191\
        );

    \I__1260\ : InMux
    port map (
            O => \N__14196\,
            I => \N__14191\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__14191\,
            I => \POWERLED.g0_i_o3_0\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__14188\,
            I => \POWERLED.un79_clk_100khzlt6_cascade_\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__14185\,
            I => \POWERLED.un79_clk_100khzlto15_5_cascade_\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__14182\,
            I => \POWERLED.un79_clk_100khzlto15_7_cascade_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14176\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__14176\,
            I => \POWERLED.un79_clk_100khzlto15_3\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__14173\,
            I => \POWERLED.count_RNIZ0Z_8_cascade_\
        );

    \I__1252\ : SRMux
    port map (
            O => \N__14170\,
            I => \N__14167\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__14167\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__1250\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__1249\ : InMux
    port map (
            O => \N__14163\,
            I => \N__14158\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__14158\,
            I => \POWERLED.N_8\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__14155\,
            I => \N__14152\
        );

    \I__1246\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14149\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__14149\,
            I => \POWERLED.un1_count_cry_0_i\
        );

    \I__1244\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14143\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__14143\,
            I => \POWERLED.count_0_12\
        );

    \I__1242\ : IoInMux
    port map (
            O => \N__14140\,
            I => \N__14137\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__14137\,
            I => \N__14134\
        );

    \I__1240\ : Span4Mux_s0_v
    port map (
            O => \N__14134\,
            I => \N__14131\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__14131\,
            I => \N__14128\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__14128\,
            I => pwrbtn_led
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__14125\,
            I => \POWERLED.curr_state_3_0_cascade_\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__14122\,
            I => \POWERLED.curr_stateZ0Z_0_cascade_\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__14119\,
            I => \POWERLED.count_0_sqmuxa_i_cascade_\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__14116\,
            I => \POWERLED.count_1_0_cascade_\
        );

    \I__1233\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14110\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__14110\,
            I => \POWERLED.count_0_0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14101\
        );

    \I__1230\ : InMux
    port map (
            O => \N__14106\,
            I => \N__14101\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__14101\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__1228\ : InMux
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__14095\,
            I => \POWERLED.count_0_5\
        );

    \I__1226\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14089\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__14089\,
            I => \POWERLED.count_0_14\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__14086\,
            I => \POWERLED.count_1_1_cascade_\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__14083\,
            I => \POWERLED.countZ0Z_1_cascade_\
        );

    \I__1222\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14077\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__14077\,
            I => \POWERLED.count_0_1\
        );

    \I__1220\ : InMux
    port map (
            O => \N__14074\,
            I => \N__14071\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__14071\,
            I => \POWERLED.count_0_3\
        );

    \I__1218\ : InMux
    port map (
            O => \N__14068\,
            I => \DSW_PWRGD.un1_count_1_cry_11\
        );

    \I__1217\ : InMux
    port map (
            O => \N__14065\,
            I => \DSW_PWRGD.un1_count_1_cry_12\
        );

    \I__1216\ : InMux
    port map (
            O => \N__14062\,
            I => \DSW_PWRGD.un1_count_1_cry_13\
        );

    \I__1215\ : InMux
    port map (
            O => \N__14059\,
            I => \bfn_1_7_0_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__14053\,
            I => \POWERLED.count_0_4\
        );

    \I__1212\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__14047\,
            I => \POWERLED.count_0_13\
        );

    \I__1210\ : InMux
    port map (
            O => \N__14044\,
            I => \DSW_PWRGD.un1_count_1_cry_2\
        );

    \I__1209\ : InMux
    port map (
            O => \N__14041\,
            I => \DSW_PWRGD.un1_count_1_cry_3\
        );

    \I__1208\ : InMux
    port map (
            O => \N__14038\,
            I => \DSW_PWRGD.un1_count_1_cry_4\
        );

    \I__1207\ : InMux
    port map (
            O => \N__14035\,
            I => \DSW_PWRGD.un1_count_1_cry_5\
        );

    \I__1206\ : InMux
    port map (
            O => \N__14032\,
            I => \DSW_PWRGD.un1_count_1_cry_6\
        );

    \I__1205\ : InMux
    port map (
            O => \N__14029\,
            I => \bfn_1_6_0_\
        );

    \I__1204\ : InMux
    port map (
            O => \N__14026\,
            I => \DSW_PWRGD.un1_count_1_cry_8\
        );

    \I__1203\ : InMux
    port map (
            O => \N__14023\,
            I => \DSW_PWRGD.un1_count_1_cry_9\
        );

    \I__1202\ : InMux
    port map (
            O => \N__14020\,
            I => \DSW_PWRGD.un1_count_1_cry_10\
        );

    \I__1201\ : InMux
    port map (
            O => \N__14017\,
            I => \HDA_STRAP.un1_count_1_cry_12\
        );

    \I__1200\ : InMux
    port map (
            O => \N__14014\,
            I => \HDA_STRAP.un1_count_1_cry_13\
        );

    \I__1199\ : InMux
    port map (
            O => \N__14011\,
            I => \HDA_STRAP.un1_count_1_cry_14\
        );

    \I__1198\ : InMux
    port map (
            O => \N__14008\,
            I => \bfn_1_3_0_\
        );

    \I__1197\ : InMux
    port map (
            O => \N__14005\,
            I => \HDA_STRAP.un1_count_1_cry_16\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__14002\,
            I => \N__13998\
        );

    \I__1195\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13987\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__13992\,
            I => \N__13987\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__13987\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_1\
        );

    \I__1190\ : InMux
    port map (
            O => \N__13984\,
            I => \DSW_PWRGD.un1_count_1_cry_0\
        );

    \I__1189\ : InMux
    port map (
            O => \N__13981\,
            I => \DSW_PWRGD.un1_count_1_cry_1\
        );

    \I__1188\ : InMux
    port map (
            O => \N__13978\,
            I => \HDA_STRAP.un1_count_1_cry_3\
        );

    \I__1187\ : InMux
    port map (
            O => \N__13975\,
            I => \HDA_STRAP.un1_count_1_cry_4\
        );

    \I__1186\ : InMux
    port map (
            O => \N__13972\,
            I => \HDA_STRAP.un1_count_1_cry_5\
        );

    \I__1185\ : InMux
    port map (
            O => \N__13969\,
            I => \HDA_STRAP.un1_count_1_cry_6\
        );

    \I__1184\ : InMux
    port map (
            O => \N__13966\,
            I => \bfn_1_2_0_\
        );

    \I__1183\ : InMux
    port map (
            O => \N__13963\,
            I => \HDA_STRAP.un1_count_1_cry_8\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13960\,
            I => \HDA_STRAP.un1_count_1_cry_9\
        );

    \I__1181\ : InMux
    port map (
            O => \N__13957\,
            I => \HDA_STRAP.un1_count_1_cry_10\
        );

    \I__1180\ : InMux
    port map (
            O => \N__13954\,
            I => \HDA_STRAP.un1_count_1_cry_11\
        );

    \I__1179\ : InMux
    port map (
            O => \N__13951\,
            I => \HDA_STRAP.un1_count_1_cry_0\
        );

    \I__1178\ : InMux
    port map (
            O => \N__13948\,
            I => \HDA_STRAP.un1_count_1_cry_1\
        );

    \I__1177\ : InMux
    port map (
            O => \N__13945\,
            I => \HDA_STRAP.un1_count_1_cry_2\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_5_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_1_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7\,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_1_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_1_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_7\,
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_15\,
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_1_7_0_\
        );

    \N_29_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22537\,
            GLOBALBUFFEROUTPUT => \N_29_g\
        );

    \N_570_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29826\,
            GLOBALBUFFEROUTPUT => \N_570_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_0_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14553\,
            in2 => \N__14002\,
            in3 => \N__14001\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_1_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14574\,
            in2 => \_gnd_net_\,
            in3 => \N__13951\,
            lcout => \HDA_STRAP.countZ0Z_1\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_0\,
            carryout => \HDA_STRAP.un1_count_1_cry_1\,
            clk => \N__34372\,
            ce => \N__34689\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14641\,
            in2 => \_gnd_net_\,
            in3 => \N__13948\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_1\,
            carryout => \HDA_STRAP.un1_count_1_cry_2\,
            clk => \N__34372\,
            ce => \N__34689\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14613\,
            in2 => \_gnd_net_\,
            in3 => \N__13945\,
            lcout => \HDA_STRAP.countZ0Z_3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_2\,
            carryout => \HDA_STRAP.un1_count_1_cry_3\,
            clk => \N__34372\,
            ce => \N__34689\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14629\,
            in2 => \_gnd_net_\,
            in3 => \N__13978\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_3\,
            carryout => \HDA_STRAP.un1_count_1_cry_4\,
            clk => \N__34372\,
            ce => \N__34689\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14602\,
            in2 => \_gnd_net_\,
            in3 => \N__13975\,
            lcout => \HDA_STRAP.countZ0Z_5\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_4\,
            carryout => \HDA_STRAP.un1_count_1_cry_5\,
            clk => \N__34372\,
            ce => \N__34689\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_6_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14767\,
            in2 => \_gnd_net_\,
            in3 => \N__13972\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_5\,
            carryout => \HDA_STRAP.un1_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14434\,
            in2 => \_gnd_net_\,
            in3 => \N__13969\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_6\,
            carryout => \HDA_STRAP.un1_count_1_cry_7\,
            clk => \N__34372\,
            ce => \N__34689\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_8_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14749\,
            in2 => \_gnd_net_\,
            in3 => \N__13966\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14461\,
            in2 => \_gnd_net_\,
            in3 => \N__13963\,
            lcout => \HDA_STRAP.countZ0Z_9\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_8\,
            carryout => \HDA_STRAP.un1_count_1_cry_9\,
            clk => \N__34389\,
            ce => \N__34711\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_10_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14485\,
            in2 => \_gnd_net_\,
            in3 => \N__13960\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_9\,
            carryout => \HDA_STRAP.un1_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_11_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14731\,
            in2 => \_gnd_net_\,
            in3 => \N__13957\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_10\,
            carryout => \HDA_STRAP.un1_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14473\,
            in2 => \_gnd_net_\,
            in3 => \N__13954\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_11\,
            carryout => \HDA_STRAP.un1_count_1_cry_12\,
            clk => \N__34389\,
            ce => \N__34711\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14448\,
            in2 => \_gnd_net_\,
            in3 => \N__14017\,
            lcout => \HDA_STRAP.countZ0Z_13\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_12\,
            carryout => \HDA_STRAP.un1_count_1_cry_13\,
            clk => \N__34389\,
            ce => \N__34711\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14796\,
            in2 => \_gnd_net_\,
            in3 => \N__14014\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_13\,
            carryout => \HDA_STRAP.un1_count_1_cry_14\,
            clk => \N__34389\,
            ce => \N__34711\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14809\,
            in2 => \_gnd_net_\,
            in3 => \N__14011\,
            lcout => \HDA_STRAP.countZ0Z_15\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_14\,
            carryout => \HDA_STRAP.un1_count_1_cry_15\,
            clk => \N__34389\,
            ce => \N__34711\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_16_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14506\,
            in2 => \_gnd_net_\,
            in3 => \N__14008\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_17_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14542\,
            in2 => \_gnd_net_\,
            in3 => \N__14005\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_1_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15006\,
            lcout => \HDA_STRAP.curr_state_RNIH91AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34866\,
            in1 => \N__15169\,
            in2 => \N__15151\,
            in3 => \N__15150\,
            lcout => \DSW_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_0\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_1_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34862\,
            in1 => \N__16566\,
            in2 => \_gnd_net_\,
            in3 => \N__13984\,
            lcout => \DSW_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_0\,
            carryout => \DSW_PWRGD.un1_count_1_cry_1\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_2_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34867\,
            in1 => \N__15265\,
            in2 => \_gnd_net_\,
            in3 => \N__13981\,
            lcout => \DSW_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_1\,
            carryout => \DSW_PWRGD.un1_count_1_cry_2\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_3_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34863\,
            in1 => \N__15226\,
            in2 => \_gnd_net_\,
            in3 => \N__14044\,
            lcout => \DSW_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_2\,
            carryout => \DSW_PWRGD.un1_count_1_cry_3\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_4_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34868\,
            in1 => \N__16515\,
            in2 => \_gnd_net_\,
            in3 => \N__14041\,
            lcout => \DSW_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_3\,
            carryout => \DSW_PWRGD.un1_count_1_cry_4\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_5_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34864\,
            in1 => \N__15253\,
            in2 => \_gnd_net_\,
            in3 => \N__14038\,
            lcout => \DSW_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_4\,
            carryout => \DSW_PWRGD.un1_count_1_cry_5\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_6_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34869\,
            in1 => \N__16551\,
            in2 => \_gnd_net_\,
            in3 => \N__14035\,
            lcout => \DSW_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_5\,
            carryout => \DSW_PWRGD.un1_count_1_cry_6\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_7_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34865\,
            in1 => \N__15240\,
            in2 => \_gnd_net_\,
            in3 => \N__14032\,
            lcout => \DSW_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_6\,
            carryout => \DSW_PWRGD.un1_count_1_cry_7\,
            clk => \N__34373\,
            ce => 'H',
            sr => \N__15326\
        );

    \DSW_PWRGD.count_8_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34891\,
            in1 => \N__15183\,
            in2 => \_gnd_net_\,
            in3 => \N__14029\,
            lcout => \DSW_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_8\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.count_9_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34879\,
            in1 => \N__16530\,
            in2 => \_gnd_net_\,
            in3 => \N__14026\,
            lcout => \DSW_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_8\,
            carryout => \DSW_PWRGD.un1_count_1_cry_9\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.count_10_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34888\,
            in1 => \N__15196\,
            in2 => \_gnd_net_\,
            in3 => \N__14023\,
            lcout => \DSW_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_9\,
            carryout => \DSW_PWRGD.un1_count_1_cry_10\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.count_11_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34877\,
            in1 => \N__15208\,
            in2 => \_gnd_net_\,
            in3 => \N__14020\,
            lcout => \DSW_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_10\,
            carryout => \DSW_PWRGD.un1_count_1_cry_11\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.count_12_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34889\,
            in1 => \N__14824\,
            in2 => \_gnd_net_\,
            in3 => \N__14068\,
            lcout => \DSW_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_11\,
            carryout => \DSW_PWRGD.un1_count_1_cry_12\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.count_13_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34878\,
            in1 => \N__14854\,
            in2 => \_gnd_net_\,
            in3 => \N__14065\,
            lcout => \DSW_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_12\,
            carryout => \DSW_PWRGD.un1_count_1_cry_13\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.count_14_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34890\,
            in1 => \N__14866\,
            in2 => \_gnd_net_\,
            in3 => \N__14062\,
            lcout => \DSW_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_13\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14\,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__15331\
        );

    \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34500\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_14\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_15_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14838\,
            in2 => \_gnd_net_\,
            in3 => \N__14059\,
            lcout => \DSW_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34444\,
            ce => \N__15292\,
            sr => \N__15330\
        );

    \POWERLED.count_RNI0LHN_4_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14056\,
            in1 => \N__30613\,
            in2 => \_gnd_net_\,
            in3 => \N__15645\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_4_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15649\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34432\,
            ce => \N__30781\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI0M6O_13_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15913\,
            in1 => \N__14050\,
            in2 => \_gnd_net_\,
            in3 => \N__30615\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_13_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15912\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34432\,
            ce => \N__30781\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI2OIN_5_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14098\,
            in1 => \N__30614\,
            in2 => \_gnd_net_\,
            in3 => \N__15606\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15610\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34432\,
            ce => \N__30781\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI2P7O_14_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15871\,
            in1 => \N__14092\,
            in2 => \_gnd_net_\,
            in3 => \N__30616\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15870\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34432\,
            ce => \N__30781\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_1_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__15479\,
            in1 => \N__15455\,
            in2 => \_gnd_net_\,
            in3 => \N__15851\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGBFE_1_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30620\,
            in2 => \N__14086\,
            in3 => \N__14080\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => \POWERLED.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15457\,
            in2 => \N__14083\,
            in3 => \N__15855\,
            lcout => \POWERLED.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => \N__30784\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__15456\,
            in1 => \_gnd_net_\,
            in2 => \N__15856\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => \N__30784\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUHGN_3_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14074\,
            in1 => \_gnd_net_\,
            in2 => \N__30631\,
            in3 => \N__15360\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15364\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => \N__30784\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUI5O_12_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__15955\,
            in1 => \N__14146\,
            in2 => \N__30632\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15954\,
            lcout => \POWERLED.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => \N__30784\,
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNIB7P12_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__14107\,
            in1 => \N__14197\,
            in2 => \N__17883\,
            in3 => \N__14164\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__17844\,
            in1 => \N__17812\,
            in2 => \_gnd_net_\,
            in3 => \N__17872\,
            lcout => OPEN,
            ltout => \POWERLED.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI2P6L_0_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17788\,
            in1 => \_gnd_net_\,
            in2 => \N__14125\,
            in3 => \N__30577\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => \POWERLED.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIE5D5_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__30578\,
            in1 => \_gnd_net_\,
            in2 => \N__14122\,
            in3 => \N__17839\,
            lcout => \POWERLED.count_0_sqmuxa_i\,
            ltout => \POWERLED.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14119\,
            in3 => \N__15458\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIFAFE_0_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30579\,
            in1 => \_gnd_net_\,
            in2 => \N__14116\,
            in3 => \N__14113\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__14106\,
            in1 => \N__14196\,
            in2 => \N__17882\,
            in3 => \N__14163\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34460\,
            ce => 'H',
            sr => \N__14170\
        );

    \POWERLED.curr_state_RNI1KAM_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30809\,
            in2 => \_gnd_net_\,
            in3 => \N__17811\,
            lcout => \POWERLED.g0_i_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_2_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__15423\,
            in1 => \_gnd_net_\,
            in2 => \N__15388\,
            in3 => \N__15669\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_5_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__15630\,
            in1 => \N__16067\,
            in2 => \N__14188\,
            in3 => \N__15731\,
            lcout => \POWERLED.un79_clk_100khzlto15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15579\,
            in1 => \N__15543\,
            in2 => \N__15942\,
            in3 => \N__15975\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_15_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__15893\,
            in1 => \_gnd_net_\,
            in2 => \N__14185\,
            in3 => \N__15686\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_8_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16019\,
            in1 => \N__15752\,
            in2 => \N__14182\,
            in3 => \N__14179\,
            lcout => \POWERLED.count_RNIZ0Z_8\,
            ltout => \POWERLED.count_RNIZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__17814\,
            in1 => \_gnd_net_\,
            in2 => \N__14173\,
            in3 => \N__30630\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIFPNR_0_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30810\,
            in1 => \N__17813\,
            in2 => \N__30636\,
            in3 => \N__17843\,
            lcout => \POWERLED.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22552\,
            in2 => \N__14155\,
            in3 => \N__15463\,
            lcout => \POWERLED.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15484\,
            in1 => \N__22399\,
            in2 => \N__14278\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5110_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20125\,
            in2 => \N__14269\,
            in3 => \N__15427\,
            lcout => \POWERLED.N_5111_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14350\,
            in2 => \N__14257\,
            in3 => \N__15387\,
            lcout => \POWERLED.N_5112_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15670\,
            in1 => \N__18709\,
            in2 => \N__14245\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5113_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15634\,
            in1 => \N__14413\,
            in2 => \N__14236\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5114_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16741\,
            in2 => \N__14227\,
            in3 => \N__15735\,
            lcout => \POWERLED.N_5115_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16071\,
            in1 => \N__16132\,
            in2 => \N__14218\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5116_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16030\,
            in1 => \N__14395\,
            in2 => \N__14206\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5117_i\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15757\,
            in1 => \N__14341\,
            in2 => \N__14404\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5118_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15583\,
            in1 => \N__14335\,
            in2 => \N__14374\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5119_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15544\,
            in1 => \N__14329\,
            in2 => \N__14362\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5120_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14323\,
            in2 => \N__14290\,
            in3 => \N__15976\,
            lcout => \POWERLED.N_5121_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15943\,
            in1 => \N__17047\,
            in2 => \N__14317\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5122_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14305\,
            in2 => \N__20188\,
            in3 => \N__15898\,
            lcout => \POWERLED.N_5123_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15694\,
            in1 => \N__14299\,
            in2 => \N__14386\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_5124_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14293\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18478\,
            lcout => \POWERLED.un85_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16255\,
            lcout => \POWERLED.un85_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18085\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16428\,
            lcout => \POWERLED.un85_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22231\,
            lcout => \POWERLED.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB5IA5_2_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14782\,
            in1 => \N__14590\,
            in2 => \N__14422\,
            in3 => \N__14524\,
            lcout => \HDA_STRAP.un4_count\,
            ltout => \HDA_STRAP.un4_count_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010101010"
        )
    port map (
            in0 => \N__14650\,
            in1 => \N__15014\,
            in2 => \N__14644\,
            in3 => \N__14941\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34195\,
            ce => \N__34688\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI2L821_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14640\,
            in1 => \N__14628\,
            in2 => \N__14617\,
            in3 => \N__14601\,
            lcout => \HDA_STRAP.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011001100"
        )
    port map (
            in0 => \N__15023\,
            in1 => \N__14584\,
            in2 => \N__14951\,
            in3 => \N__14710\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34195\,
            ce => \N__34688\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI4CB61_17_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__14502\,
            in1 => \N__14575\,
            in2 => \N__14563\,
            in3 => \N__14538\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIH7IR1_10_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14730\,
            in2 => \N__14527\,
            in3 => \N__14484\,
            lcout => \HDA_STRAP.un4_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__14708\,
            in1 => \N__14937\,
            in2 => \N__14518\,
            in3 => \N__15027\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34195\,
            ce => \N__34688\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__14936\,
            in1 => \N__14491\,
            in2 => \N__15028\,
            in3 => \N__14709\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34195\,
            ce => \N__34688\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIBJB61_7_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14472\,
            in1 => \N__14460\,
            in2 => \N__14449\,
            in3 => \N__14433\,
            lcout => \HDA_STRAP.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDLB61_6_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__14808\,
            in1 => \N__14748\,
            in2 => \N__14797\,
            in3 => \N__14766\,
            lcout => \HDA_STRAP.un4_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011001100"
        )
    port map (
            in0 => \N__15019\,
            in1 => \N__14773\,
            in2 => \N__14953\,
            in3 => \N__14715\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34388\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__14713\,
            in1 => \N__14755\,
            in2 => \N__14950\,
            in3 => \N__15021\,
            lcout => \HDA_STRAP.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34388\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011001100"
        )
    port map (
            in0 => \N__15018\,
            in1 => \N__14737\,
            in2 => \N__14952\,
            in3 => \N__14714\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34388\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__14712\,
            in1 => \N__15020\,
            in2 => \N__14949\,
            in3 => \N__18764\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34388\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_1_2_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15017\,
            in1 => \N__14929\,
            in2 => \_gnd_net_\,
            in3 => \N__14711\,
            lcout => OPEN,
            ltout => \HDA_STRAP.N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000001100"
        )
    port map (
            in0 => \N__15022\,
            in1 => \N__14676\,
            in2 => \N__14719\,
            in3 => \N__14872\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34388\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_0_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000111111"
        )
    port map (
            in0 => \N__14716\,
            in1 => \N__20436\,
            in2 => \N__31177\,
            in3 => \N__14923\,
            lcout => \HDA_STRAP.curr_state_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__15016\,
            in1 => \N__14677\,
            in2 => \_gnd_net_\,
            in3 => \N__14928\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34322\,
            ce => \N__34706\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_1_0_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101110000"
        )
    port map (
            in0 => \N__20437\,
            in1 => \N__31176\,
            in2 => \N__14948\,
            in3 => \N__15040\,
            lcout => OPEN,
            ltout => \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15015\,
            in2 => \N__14962\,
            in3 => \N__14959\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34322\,
            ce => \N__34706\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_2_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14924\,
            in2 => \_gnd_net_\,
            in3 => \N__18753\,
            lcout => \HDA_STRAP.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25620\,
            lcout => \POWERLED.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34390\,
            ce => \N__25596\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25755\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34390\,
            ce => \N__25596\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25689\,
            lcout => \POWERLED.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34390\,
            ce => \N__25596\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19015\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34390\,
            ce => \N__25596\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14865\,
            in1 => \N__14853\,
            in2 => \N__14842\,
            in3 => \N__14823\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIB8TE4_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15157\,
            in1 => \N__15214\,
            in2 => \N__14812\,
            in3 => \N__16501\,
            lcout => \DSW_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21300\,
            in2 => \_gnd_net_\,
            in3 => \N__21805\,
            lcout => \POWERLED.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIH71P_2_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15264\,
            in1 => \N__15252\,
            in2 => \N__15241\,
            in3 => \N__15225\,
            lcout => \DSW_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIBCB91_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15207\,
            in1 => \N__15195\,
            in2 => \N__15184\,
            in3 => \N__15168\,
            lcout => \DSW_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.DSW_PWROK_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__15134\,
            in1 => \N__15111\,
            in2 => \N__15088\,
            in3 => \_gnd_net_\,
            lcout => dsw_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => \N__34713\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNIADII_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__15116\,
            in1 => \N__15075\,
            in2 => \_gnd_net_\,
            in3 => \N__15132\,
            lcout => \DSW_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_0_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101001000000"
        )
    port map (
            in0 => \N__15135\,
            in1 => \N__15112\,
            in2 => \N__15087\,
            in3 => \N__15054\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => \N__34713\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_1_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__15085\,
            in1 => \N__15058\,
            in2 => \N__15118\,
            in3 => \N__15136\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => \N__34713\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111011"
        )
    port map (
            in0 => \N__15133\,
            in1 => \N__15117\,
            in2 => \N__15086\,
            in3 => \N__15053\,
            lcout => OPEN,
            ltout => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_27_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15334\,
            in3 => \N__34841\,
            lcout => \G_27\,
            ltout => \G_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNO_0_15_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__34842\,
            in1 => \_gnd_net_\,
            in2 => \N__15295\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.N_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_9_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__21125\,
            in1 => \N__20968\,
            in2 => \_gnd_net_\,
            in3 => \N__20809\,
            lcout => OPEN,
            ltout => \POWERLED.d_i1_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_16_9_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001111"
        )
    port map (
            in0 => \N__19314\,
            in1 => \N__16489\,
            in2 => \N__15283\,
            in3 => \N__15273\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_16Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__21568\,
            in1 => \N__20811\,
            in2 => \N__15280\,
            in3 => \N__21949\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_9_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000001000"
        )
    port map (
            in0 => \N__20808\,
            in1 => \N__21124\,
            in2 => \N__20971\,
            in3 => \N__27160\,
            lcout => \POWERLED.un1_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_9_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010011010011"
        )
    port map (
            in0 => \N__27161\,
            in1 => \N__20969\,
            in2 => \N__21137\,
            in3 => \N__20810\,
            lcout => OPEN,
            ltout => \POWERLED.d_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \N__23278\,
            in1 => \N__16653\,
            in2 => \N__15277\,
            in3 => \N__15274\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__22140\,
            in1 => \N__21777\,
            in2 => \N__23797\,
            in3 => \N__26599\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_0_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__22139\,
            in2 => \_gnd_net_\,
            in3 => \N__22383\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110000111"
        )
    port map (
            in0 => \N__21802\,
            in1 => \N__22141\,
            in2 => \N__15346\,
            in3 => \N__26604\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_2_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__23792\,
            in1 => \_gnd_net_\,
            in2 => \N__15349\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_2_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__21296\,
            in1 => \N__23791\,
            in2 => \_gnd_net_\,
            in3 => \N__27117\,
            lcout => \POWERLED.un1_dutycycle_53_axb_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_9_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101000"
        )
    port map (
            in0 => \N__27118\,
            in1 => \N__20815\,
            in2 => \N__16654\,
            in3 => \N__21129\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__21130\,
            in1 => \N__20937\,
            in2 => \N__15337\,
            in3 => \N__21451\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21298\,
            in2 => \_gnd_net_\,
            in3 => \N__22382\,
            lcout => \POWERLED.mult1_un145_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_10_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__20938\,
            in1 => \N__21955\,
            in2 => \_gnd_net_\,
            in3 => \N__27119\,
            lcout => \POWERLED.g0_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_3_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21131\,
            in1 => \N__21803\,
            in2 => \_gnd_net_\,
            in3 => \N__21297\,
            lcout => \POWERLED.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15772\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34445\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIJKSP_10_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__15502\,
            in2 => \_gnd_net_\,
            in3 => \N__30604\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15558\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34445\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNISEFN_2_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15496\,
            in2 => \N__15403\,
            in3 => \N__30603\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15402\,
            lcout => \POWERLED.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34445\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNISF4O_11_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15517\,
            in1 => \N__15490\,
            in2 => \_gnd_net_\,
            in3 => \N__30605\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15516\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34445\,
            ce => \N__30783\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15480\,
            in2 => \N__15462\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIB209_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15838\,
            in1 => \N__15422\,
            in2 => \_gnd_net_\,
            in3 => \N__15391\,
            lcout => \POWERLED.count_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIC419_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15841\,
            in1 => \N__15383\,
            in2 => \_gnd_net_\,
            in3 => \N__15352\,
            lcout => \POWERLED.count_1_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2\,
            carryout => \POWERLED.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNID629_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15837\,
            in1 => \N__15668\,
            in2 => \_gnd_net_\,
            in3 => \N__15637\,
            lcout => \POWERLED.count_1_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3\,
            carryout => \POWERLED.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNIE839_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15842\,
            in1 => \N__15629\,
            in2 => \_gnd_net_\,
            in3 => \N__15598\,
            lcout => \POWERLED.count_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNIFA49_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15839\,
            in1 => \N__15736\,
            in2 => \_gnd_net_\,
            in3 => \N__15595\,
            lcout => \POWERLED.count_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIGC59_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15843\,
            in1 => \N__16072\,
            in2 => \_gnd_net_\,
            in3 => \N__15592\,
            lcout => \POWERLED.count_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIHE69_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15840\,
            in1 => \N__16026\,
            in2 => \_gnd_net_\,
            in3 => \N__15589\,
            lcout => \POWERLED.count_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNIIG79_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15844\,
            in1 => \N__15753\,
            in2 => \_gnd_net_\,
            in3 => \N__15586\,
            lcout => \POWERLED.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNIJI89_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15849\,
            in1 => \N__15578\,
            in2 => \_gnd_net_\,
            in3 => \N__15547\,
            lcout => \POWERLED.count_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15846\,
            in1 => \N__15536\,
            in2 => \_gnd_net_\,
            in3 => \N__15505\,
            lcout => \POWERLED.count_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNISEH7_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15848\,
            in1 => \N__15974\,
            in2 => \_gnd_net_\,
            in3 => \N__15946\,
            lcout => \POWERLED.count_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11_cZ0\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNITGI7_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15845\,
            in1 => \N__15941\,
            in2 => \_gnd_net_\,
            in3 => \N__15901\,
            lcout => \POWERLED.count_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15847\,
            in1 => \N__15897\,
            in2 => \_gnd_net_\,
            in3 => \N__15859\,
            lcout => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13_cZ0\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__15687\,
            in1 => \N__15850\,
            in2 => \_gnd_net_\,
            in3 => \N__15787\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIA4NN_9_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30606\,
            in1 => \N__15784\,
            in2 => \_gnd_net_\,
            in3 => \N__15768\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI4RJN_6_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15700\,
            in1 => \N__30600\,
            in2 => \_gnd_net_\,
            in3 => \N__15711\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15715\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34459\,
            ce => \N__30785\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI4S8O_15_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16078\,
            in1 => \N__30599\,
            in2 => \_gnd_net_\,
            in3 => \N__16086\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16090\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34459\,
            ce => \N__30785\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI6UKN_7_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16036\,
            in1 => \N__30601\,
            in2 => \_gnd_net_\,
            in3 => \N__16047\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16051\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34459\,
            ce => \N__30785\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI81MN_8_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__15991\,
            in1 => \N__30602\,
            in2 => \N__16006\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16005\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34459\,
            ce => \N__30785\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19711\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16873\,
            in2 => \N__16214\,
            in3 => \N__15985\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16126\,
            in2 => \N__16216\,
            in3 => \N__15982\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16117\,
            in2 => \N__16253\,
            in3 => \N__15979\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16108\,
            in2 => \N__16254\,
            in3 => \N__16144\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16989\,
            in1 => \N__16099\,
            in2 => \N__16215\,
            in3 => \N__16141\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16138\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => \POWERLED.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16135\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19672\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16765\,
            in2 => \N__16350\,
            in3 => \N__16120\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16346\,
            in2 => \N__16192\,
            in3 => \N__16111\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16180\,
            in2 => \N__16383\,
            in3 => \N__16102\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16171\,
            in2 => \N__16384\,
            in3 => \N__16093\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16243\,
            in1 => \N__16162\,
            in2 => \N__16351\,
            in3 => \N__16261\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16153\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16258\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16242\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19633\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16397\,
            in2 => \N__20092\,
            in3 => \N__16183\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16333\,
            in2 => \N__16402\,
            in3 => \N__16174\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16424\,
            in2 => \N__16324\,
            in3 => \N__16165\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16312\,
            in2 => \N__16429\,
            in3 => \N__16156\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16375\,
            in1 => \N__16401\,
            in2 => \N__16303\,
            in3 => \N__16147\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16276\,
            in2 => \_gnd_net_\,
            in3 => \N__16387\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => \POWERLED.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16354\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20116\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16287\,
            in2 => \N__20236\,
            in3 => \N__16327\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2_c\,
            carryout => \POWERLED.mult1_un96_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17026\,
            in2 => \N__16291\,
            in3 => \N__16315\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3_c\,
            carryout => \POWERLED.mult1_un96_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17353\,
            in2 => \N__17280\,
            in3 => \N__16306\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4_c\,
            carryout => \POWERLED.mult1_un96_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17275\,
            in2 => \N__17341\,
            in3 => \N__16294\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5_c\,
            carryout => \POWERLED.mult1_un96_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16423\,
            in1 => \N__16286\,
            in2 => \N__17326\,
            in3 => \N__16270\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6_c\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16432\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => \POWERLED.mult1_un96_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16405\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17212\,
            in1 => \N__17192\,
            in2 => \N__17146\,
            in3 => \N__17168\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17169\,
            in1 => \N__25096\,
            in2 => \_gnd_net_\,
            in3 => \N__17155\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000110"
        )
    port map (
            in0 => \N__17223\,
            in1 => \N__17241\,
            in2 => \N__25119\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000010010"
        )
    port map (
            in0 => \N__17409\,
            in1 => \N__25099\,
            in2 => \N__17395\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__17179\,
            in1 => \_gnd_net_\,
            in2 => \N__25120\,
            in3 => \N__17193\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__25097\,
            in2 => \_gnd_net_\,
            in3 => \N__17125\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17382\,
            in1 => \N__17408\,
            in2 => \N__17440\,
            in3 => \N__17240\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17439\,
            in1 => \N__25098\,
            in2 => \_gnd_net_\,
            in3 => \N__17419\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI94A94_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20430\,
            in2 => \_gnd_net_\,
            in3 => \N__31166\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25106\,
            in2 => \_gnd_net_\,
            in3 => \N__17219\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIV3O1A_4_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__26918\,
            in1 => \N__16459\,
            in2 => \N__25591\,
            in3 => \N__19074\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26920\,
            lcout => \POWERLED.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34271\,
            ce => \N__25597\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19075\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34271\,
            ce => \N__25597\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI7GS1A_8_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16453\,
            in1 => \N__19011\,
            in2 => \_gnd_net_\,
            in3 => \N__25579\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => \POWERLED.count_offZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_3_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19119\,
            in1 => \N__19053\,
            in2 => \N__16444\,
            in3 => \N__19090\,
            lcout => \POWERLED.un34_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIT0N1A_3_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__19104\,
            in1 => \N__25574\,
            in2 => \N__16441\,
            in3 => \N__26917\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34271\,
            ce => \N__25597\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI5DR1A_7_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16573\,
            in1 => \N__19038\,
            in2 => \_gnd_net_\,
            in3 => \N__25578\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIKA1P_1_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16567\,
            in1 => \N__16552\,
            in2 => \N__16537\,
            in3 => \N__16516\,
            lcout => \DSW_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__21105\,
            in1 => \_gnd_net_\,
            in2 => \N__21278\,
            in3 => \N__21766\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__20942\,
            in1 => \N__21796\,
            in2 => \N__16492\,
            in3 => \N__26603\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__21241\,
            in1 => \N__21762\,
            in2 => \_gnd_net_\,
            in3 => \N__20940\,
            lcout => \POWERLED.un1_dutycycle_53_20_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100011111"
        )
    port map (
            in0 => \N__20941\,
            in1 => \N__21242\,
            in2 => \N__21801\,
            in3 => \N__21104\,
            lcout => OPEN,
            ltout => \POWERLED.o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_9_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001111"
        )
    port map (
            in0 => \N__19297\,
            in1 => \N__16482\,
            in2 => \N__16471\,
            in3 => \N__20805\,
            lcout => \POWERLED.un1_dutycycle_53_axb_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__20939\,
            in1 => \N__21240\,
            in2 => \N__21800\,
            in3 => \N__21103\,
            lcout => \POWERLED.un1_dutycycle_53_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_9_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100110100110"
        )
    port map (
            in0 => \N__16594\,
            in1 => \N__20806\,
            in2 => \N__16468\,
            in3 => \N__27152\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_10_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__21900\,
            in1 => \_gnd_net_\,
            in2 => \N__16600\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001000"
        )
    port map (
            in0 => \N__21062\,
            in1 => \N__21728\,
            in2 => \N__21279\,
            in3 => \N__20949\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_3\,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_9_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__20807\,
            in1 => \N__27151\,
            in2 => \N__16597\,
            in3 => \N__26602\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_10_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21896\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_1_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011111"
        )
    port map (
            in0 => \N__21729\,
            in1 => \_gnd_net_\,
            in2 => \N__22145\,
            in3 => \N__26601\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__21249\,
            in1 => \N__19732\,
            in2 => \N__16588\,
            in3 => \N__27153\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__20950\,
            in1 => \_gnd_net_\,
            in2 => \N__21926\,
            in3 => \N__21064\,
            lcout => \POWERLED.un1_dutycycle_53_8_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_11_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000110011"
        )
    port map (
            in0 => \N__16585\,
            in1 => \N__21385\,
            in2 => \N__21450\,
            in3 => \N__23265\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_11_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16639\,
            in1 => \N__16612\,
            in2 => \N__16579\,
            in3 => \N__16660\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_8_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \N__21566\,
            in1 => \N__16618\,
            in2 => \N__16576\,
            in3 => \N__27142\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21102\,
            in1 => \N__21892\,
            in2 => \N__23273\,
            in3 => \N__20920\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_3Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001110"
        )
    port map (
            in0 => \N__21894\,
            in1 => \N__20776\,
            in2 => \N__16663\,
            in3 => \N__23261\,
            lcout => \POWERLED.un1_dutycycle_53_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16640\,
            in1 => \N__20924\,
            in2 => \N__23274\,
            in3 => \N__21895\,
            lcout => \POWERLED.un1_dutycycle_53_56_a0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21893\,
            in1 => \N__27141\,
            in2 => \N__20951\,
            in3 => \N__23260\,
            lcout => \POWERLED.un1_dutycycle_53_56_a1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_9_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__20775\,
            in1 => \N__20919\,
            in2 => \N__21388\,
            in3 => \N__21891\,
            lcout => \POWERLED.un1_dutycycle_53_50_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16696\,
            in1 => \N__20830\,
            in2 => \N__29811\,
            in3 => \N__16690\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34368\,
            ce => 'H',
            sr => \N__23685\
        );

    \POWERLED.dutycycle_RNI2O4A1_13_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__26049\,
            in1 => \N__21555\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_45_and_i_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5MDM4_13_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23372\,
            in1 => \N__25861\,
            in2 => \N__16606\,
            in3 => \N__23464\,
            lcout => OPEN,
            ltout => \POWERLED.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRBF58_13_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__26767\,
            in1 => \N__29774\,
            in2 => \N__16603\,
            in3 => \N__23073\,
            lcout => \POWERLED.dutycycle_en_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3U8C3_8_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__23371\,
            in1 => \N__26048\,
            in2 => \N__25872\,
            in3 => \N__20913\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQN4F7_8_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__23463\,
            in1 => \N__26765\,
            in2 => \N__16699\,
            in3 => \N__23072\,
            lcout => \POWERLED.dutycycle_eena_3\,
            ltout => \POWERLED.dutycycle_eena_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITTBN9_8_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__29773\,
            in1 => \N__16689\,
            in2 => \N__16678\,
            in3 => \N__20829\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => \POWERLED.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_10_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__21925\,
            in1 => \_gnd_net_\,
            in2 => \N__16675\,
            in3 => \N__21061\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_9_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__20931\,
            in1 => \N__20812\,
            in2 => \N__21387\,
            in3 => \N__21106\,
            lcout => \POWERLED.un1_dutycycle_53_4_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21380\,
            in2 => \N__21951\,
            in3 => \N__23247\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__20932\,
            in1 => \N__19315\,
            in2 => \N__16672\,
            in3 => \N__16669\,
            lcout => \POWERLED.un1_dutycycle_53_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17754\,
            in2 => \_gnd_net_\,
            in3 => \N__17907\,
            lcout => \POWERLED.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_14_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__21381\,
            in1 => \_gnd_net_\,
            in2 => \N__23268\,
            in3 => \N__25376\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_13_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20813\,
            in1 => \N__21567\,
            in2 => \N__16729\,
            in3 => \N__25405\,
            lcout => \POWERLED.un2_count_clk_17_0_a2_5\,
            ltout => \POWERLED.un2_count_clk_17_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_3_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20933\,
            in1 => \N__21307\,
            in2 => \N__16726\,
            in3 => \N__21107\,
            lcout => \POWERLED.m18_e_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19771\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16774\,
            in3 => \N__16723\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16705\,
            in2 => \N__17707\,
            in3 => \N__16720\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34556\,
            in2 => \N__17686\,
            in3 => \N__16717\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34561\,
            in2 => \N__17923\,
            in3 => \N__16714\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18214\,
            in1 => \N__18004\,
            in2 => \N__17986\,
            in3 => \N__16711\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17908\,
            in2 => \N__17758\,
            in3 => \N__16708\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__17702\,
            in1 => \N__17703\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.slp_s3n_signal_i_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__27340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26412\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19882\,
            lcout => \POWERLED.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_SUSn_RNIN4K9_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24886\,
            lcout => v33a_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17103\,
            in1 => \N__16935\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19389\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17104\,
            in2 => \_gnd_net_\,
            in3 => \N__16887\,
            lcout => \POWERLED.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_10_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20943\,
            in1 => \N__24114\,
            in2 => \N__19943\,
            in3 => \N__21952\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19707\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19671\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19390\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16973\,
            in2 => \N__16861\,
            in3 => \N__16852\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16849\,
            in2 => \N__16978\,
            in3 => \N__16840\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16837\,
            in2 => \N__17002\,
            in3 => \N__16828\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17001\,
            in2 => \N__16825\,
            in3 => \N__16813\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17101\,
            in1 => \N__16977\,
            in2 => \N__16810\,
            in3 => \N__16798\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17005\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20290\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17077\,
            in2 => \N__16963\,
            in3 => \N__16951\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16948\,
            in2 => \N__16939\,
            in3 => \N__16924\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17106\,
            in2 => \N__16921\,
            in3 => \N__16912\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16909\,
            in2 => \N__17110\,
            in3 => \N__16903\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18465\,
            in1 => \N__16900\,
            in2 => \N__16891\,
            in3 => \N__16876\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17113\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17105\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19558\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18251\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30213\,
            in2 => \_gnd_net_\,
            in3 => \N__17071\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18553\,
            lcout => \POWERLED.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20257\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17309\,
            in2 => \N__17035\,
            in3 => \N__17017\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17311\,
            in2 => \N__18379\,
            in3 => \N__17344\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18355\,
            in2 => \N__18267\,
            in3 => \N__17329\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18263\,
            in2 => \N__18334\,
            in3 => \N__17314\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17260\,
            in1 => \N__17310\,
            in2 => \N__18313\,
            in3 => \N__17287\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18289\,
            in2 => \_gnd_net_\,
            in3 => \N__17284\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17242\,
            in2 => \N__17227\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_1_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17194\,
            in2 => \_gnd_net_\,
            in3 => \N__17173\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17170\,
            in2 => \_gnd_net_\,
            in3 => \N__17149\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17144\,
            in2 => \_gnd_net_\,
            in3 => \N__17443\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17438\,
            in2 => \_gnd_net_\,
            in3 => \N__17413\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17410\,
            in2 => \_gnd_net_\,
            in3 => \N__17386\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17383\,
            in2 => \_gnd_net_\,
            in3 => \N__17371\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__34020\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18697\,
            in2 => \_gnd_net_\,
            in3 => \N__17368\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__34020\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18672\,
            in2 => \_gnd_net_\,
            in3 => \N__17365\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18685\,
            in2 => \_gnd_net_\,
            in3 => \N__17362\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18658\,
            in2 => \_gnd_net_\,
            in3 => \N__17359\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18621\,
            in2 => \_gnd_net_\,
            in3 => \N__17356\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18634\,
            in2 => \_gnd_net_\,
            in3 => \N__17470\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18646\,
            in2 => \_gnd_net_\,
            in3 => \N__17467\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18607\,
            in2 => \_gnd_net_\,
            in3 => \N__17464\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18841\,
            in2 => \_gnd_net_\,
            in3 => \N__17461\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__34163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18802\,
            in2 => \_gnd_net_\,
            in3 => \N__17458\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18829\,
            in2 => \_gnd_net_\,
            in3 => \N__17455\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18816\,
            in2 => \_gnd_net_\,
            in3 => \N__17452\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18922\,
            in2 => \_gnd_net_\,
            in3 => \N__17449\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18936\,
            in2 => \_gnd_net_\,
            in3 => \N__17446\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18949\,
            in2 => \_gnd_net_\,
            in3 => \N__17497\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18961\,
            in2 => \_gnd_net_\,
            in3 => \N__17494\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18901\,
            in2 => \_gnd_net_\,
            in3 => \N__17491\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__34185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18862\,
            in2 => \_gnd_net_\,
            in3 => \N__17488\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18876\,
            in2 => \_gnd_net_\,
            in3 => \N__17485\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18889\,
            in2 => \_gnd_net_\,
            in3 => \N__17482\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17566\,
            in3 => \N__17479\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17530\,
            in3 => \N__17476\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17545\,
            in3 => \N__17473\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17569\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17562\,
            in1 => \N__17553\,
            in2 => \N__17544\,
            in3 => \N__17526\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18988\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34196\,
            ce => \N__25590\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI9JT1A_9_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17518\,
            in1 => \N__25550\,
            in2 => \_gnd_net_\,
            in3 => \N__18987\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => \POWERLED.count_offZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_10_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19189\,
            in1 => \N__19215\,
            in2 => \N__17512\,
            in3 => \N__19165\,
            lcout => \POWERLED.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIIT20A_10_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17509\,
            in1 => \N__25551\,
            in2 => \_gnd_net_\,
            in3 => \N__19200\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34196\,
            ce => \N__25590\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIR4GU9_11_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17503\,
            in1 => \N__25552\,
            in2 => \_gnd_net_\,
            in3 => \N__19176\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34196\,
            ce => \N__25590\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIT7HU9_12_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19129\,
            in1 => \N__25553\,
            in2 => \_gnd_net_\,
            in3 => \N__19140\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3U8C3_3_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__26047\,
            in1 => \N__25865\,
            in2 => \N__23380\,
            in3 => \N__21267\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQN4F7_3_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__23070\,
            in1 => \N__26770\,
            in2 => \N__17617\,
            in3 => \N__23459\,
            lcout => \POWERLED.dutycycle_eena_8\,
            ltout => \POWERLED.dutycycle_eena_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJE6N9_3_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__21184\,
            in1 => \N__29821\,
            in2 => \N__17614\,
            in3 => \N__17604\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__17605\,
            in1 => \N__17611\,
            in2 => \N__29830\,
            in3 => \N__21183\,
            lcout => \POWERLED.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34349\,
            ce => 'H',
            sr => \N__23698\
        );

    \POWERLED.dutycycle_RNI8U6P9_10_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__17577\,
            in1 => \N__29820\,
            in2 => \N__17590\,
            in3 => \N__20682\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => \POWERLED.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3U8C3_10_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25864\,
            in1 => \N__23376\,
            in2 => \N__17596\,
            in3 => \N__26046\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQN4F7_10_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__26769\,
            in1 => \N__23458\,
            in2 => \N__17593\,
            in3 => \N__23069\,
            lcout => \POWERLED.dutycycle_eena_4\,
            ltout => \POWERLED.dutycycle_eena_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__20683\,
            in1 => \N__29825\,
            in2 => \N__17581\,
            in3 => \N__17578\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34349\,
            ce => 'H',
            sr => \N__23698\
        );

    \POWERLED.dutycycle_RNIQN4F7_7_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26741\,
            in1 => \N__23460\,
            in2 => \N__23074\,
            in3 => \N__17668\,
            lcout => \POWERLED.dutycycle_eena_5\,
            ltout => \POWERLED.dutycycle_eena_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNII46M9_7_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__29812\,
            in1 => \N__17628\,
            in2 => \N__17674\,
            in3 => \N__20985\,
            lcout => \POWERLED.dutycycleZ1Z_5\,
            ltout => \POWERLED.dutycycleZ1Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3U8C3_7_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25862\,
            in1 => \N__23374\,
            in2 => \N__17671\,
            in3 => \N__26036\,
            lcout => \POWERLED.dutycycle_eena_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILH7N9_4_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__17646\,
            in1 => \N__17656\,
            in2 => \N__29828\,
            in3 => \N__21166\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3U8C3_4_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25863\,
            in1 => \N__23375\,
            in2 => \N__17662\,
            in3 => \N__26037\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQN4F7_4_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__23461\,
            in1 => \N__26742\,
            in2 => \N__17659\,
            in3 => \N__23068\,
            lcout => \POWERLED.dutycycle_eena_6\,
            ltout => \POWERLED.dutycycle_eena_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__17647\,
            in1 => \N__29816\,
            in2 => \N__17650\,
            in3 => \N__21162\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34323\,
            ce => 'H',
            sr => \N__23696\
        );

    \POWERLED.dutycycle_7_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__17635\,
            in1 => \N__20986\,
            in2 => \N__29829\,
            in3 => \N__17629\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34323\,
            ce => 'H',
            sr => \N__23696\
        );

    \POWERLED.dutycycle_RNI5MDM4_15_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__17740\,
            in1 => \N__23462\,
            in2 => \N__25873\,
            in3 => \N__23373\,
            lcout => OPEN,
            ltout => \POWERLED.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRBF58_15_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__26766\,
            in1 => \N__23071\,
            in2 => \N__17620\,
            in3 => \N__29778\,
            lcout => \POWERLED.dutycycle_en_12\,
            ltout => \POWERLED.dutycycle_en_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__17727\,
            in1 => \N__29987\,
            in2 => \N__17743\,
            in3 => \N__21463\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34223\,
            ce => 'H',
            sr => \N__23670\
        );

    \POWERLED.dutycycle_RNI2O4A1_15_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25406\,
            lcout => \POWERLED.un1_clk_100khz_48_and_i_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIPUS6A_15_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__17734\,
            in1 => \N__29986\,
            in2 => \N__17728\,
            in3 => \N__21462\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => \POWERLED.dutycycleZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17716\,
            in3 => \N__23267\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100111100"
        )
    port map (
            in0 => \N__17767\,
            in1 => \N__19459\,
            in2 => \N__17713\,
            in3 => \N__21434\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17710\,
            in3 => \N__25407\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19878\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17968\,
            in3 => \N__17689\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17977\,
            in3 => \N__17677\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34537\,
            in2 => \N__18013\,
            in3 => \N__17914\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17911\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__22146\,
            in1 => \N__32968\,
            in2 => \N__22384\,
            in3 => \N__21109\,
            lcout => \POWERLED.g2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111101010000"
        )
    port map (
            in0 => \N__19453\,
            in1 => \N__25378\,
            in2 => \N__17896\,
            in3 => \N__21529\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21784\,
            in1 => \N__21280\,
            in2 => \_gnd_net_\,
            in3 => \N__21108\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17887\,
            in2 => \N__17851\,
            in3 => \N__17818\,
            lcout => \POWERLED.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34357\,
            ce => \N__30782\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_9_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010000"
        )
    port map (
            in0 => \N__17776\,
            in1 => \N__19237\,
            in2 => \N__20814\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_9Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__19857\,
            in1 => \_gnd_net_\,
            in2 => \N__19816\,
            in3 => \N__19836\,
            lcout => \POWERLED.mult1_un40_sum_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19856\,
            in2 => \N__19837\,
            in3 => \N__19812\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__18002\,
            in1 => \N__18003\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19858\,
            in3 => \N__19832\,
            lcout => \POWERLED.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19852\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19794\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19753\,
            in2 => \N__18192\,
            in3 => \N__17959\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18188\,
            in2 => \N__17956\,
            in3 => \N__17947\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17944\,
            in2 => \N__18220\,
            in3 => \N__17938\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18218\,
            in2 => \N__17935\,
            in3 => \N__17926\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18070\,
            in1 => \N__18133\,
            in2 => \N__18193\,
            in3 => \N__18127\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18124\,
            in3 => \N__18115\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => \POWERLED.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18112\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19990\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19783\,
            in2 => \N__18033\,
            in3 => \N__18109\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18029\,
            in2 => \N__18106\,
            in3 => \N__18097\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18094\,
            in2 => \N__18078\,
            in3 => \N__18088\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18074\,
            in2 => \N__18052\,
            in3 => \N__18043\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20212\,
            in1 => \N__18040\,
            in2 => \N__18034\,
            in3 => \N__18016\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18229\,
            in2 => \_gnd_net_\,
            in3 => \N__18223\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18219\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20170\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18389\,
            in2 => \N__19972\,
            in3 => \N__18175\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18172\,
            in2 => \N__18394\,
            in3 => \N__18166\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18163\,
            in2 => \N__20221\,
            in3 => \N__18157\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18154\,
            in2 => \N__20220\,
            in3 => \N__18148\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18543\,
            in1 => \N__18393\,
            in2 => \N__18145\,
            in3 => \N__18136\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18397\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20213\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19554\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18518\,
            in2 => \N__20152\,
            in3 => \N__18367\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18364\,
            in2 => \N__18523\,
            in3 => \N__18346\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18545\,
            in2 => \N__18343\,
            in3 => \N__18322\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18319\,
            in2 => \N__18552\,
            in3 => \N__18301\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18250\,
            in1 => \N__18522\,
            in2 => \N__18298\,
            in3 => \N__18280\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18271\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18544\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20143\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18434\,
            in2 => \N__20266\,
            in3 => \N__18508\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18505\,
            in2 => \N__18439\,
            in3 => \N__18499\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18467\,
            in2 => \N__18496\,
            in3 => \N__18487\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18484\,
            in2 => \N__18474\,
            in3 => \N__18442\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20323\,
            in1 => \N__18438\,
            in2 => \N__18424\,
            in3 => \N__18415\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18412\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18406\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => \POWERLED.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18712\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18696\,
            in1 => \N__18684\,
            in2 => \N__18673\,
            in3 => \N__18657\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18645\,
            in1 => \N__18633\,
            in2 => \N__18622\,
            in3 => \N__18606\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18595\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18583\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18562\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18790\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18850\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18964\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18960\,
            in1 => \N__18948\,
            in2 => \N__18937\,
            in3 => \N__18921\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18900\,
            in1 => \N__18888\,
            in2 => \N__18877\,
            in3 => \N__18861\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18840\,
            in1 => \N__18828\,
            in2 => \N__18817\,
            in3 => \N__18801\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_PWRGD_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30424\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22945\,
            in2 => \N__22846\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNI22EQ2_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26907\,
            in1 => \N__25456\,
            in2 => \_gnd_net_\,
            in3 => \N__19123\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19120\,
            in2 => \_gnd_net_\,
            in3 => \N__19093\,
            lcout => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19089\,
            in2 => \_gnd_net_\,
            in3 => \N__19063\,
            lcout => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNI58HQ2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26908\,
            in1 => \N__25735\,
            in2 => \_gnd_net_\,
            in3 => \N__19060\,
            lcout => \POWERLED.count_off_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNI6AIQ2_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26905\,
            in1 => \N__25669\,
            in2 => \_gnd_net_\,
            in3 => \N__19057\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNI7CJQ2_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26909\,
            in1 => \N__19054\,
            in2 => \_gnd_net_\,
            in3 => \N__19027\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNI8EKQ2_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26906\,
            in1 => \N__19024\,
            in2 => \_gnd_net_\,
            in3 => \N__18997\,
            lcout => \POWERLED.count_off_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNI9GLQ2_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26910\,
            in1 => \N__18994\,
            in2 => \_gnd_net_\,
            in3 => \N__18979\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNIAIMQ2_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26913\,
            in1 => \_gnd_net_\,
            in2 => \N__19216\,
            in3 => \N__19192\,
            lcout => \POWERLED.count_off_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNIIO3P2_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26911\,
            in1 => \N__19188\,
            in2 => \_gnd_net_\,
            in3 => \N__19168\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNIJQ4P2_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26914\,
            in1 => \N__19164\,
            in2 => \_gnd_net_\,
            in3 => \N__19153\,
            lcout => \POWERLED.count_off_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNIKS5P2_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26912\,
            in1 => \N__20553\,
            in2 => \_gnd_net_\,
            in3 => \N__19150\,
            lcout => \POWERLED.count_off_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNILU6P2_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26915\,
            in1 => \N__20538\,
            in2 => \_gnd_net_\,
            in3 => \N__19147\,
            lcout => \POWERLED.count_off_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIM08P2_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__20560\,
            in1 => \N__26916\,
            in2 => \_gnd_net_\,
            in3 => \N__19144\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19141\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34013\,
            ce => \N__25592\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001000"
        )
    port map (
            in0 => \N__21889\,
            in1 => \N__20772\,
            in2 => \N__21122\,
            in3 => \N__20964\,
            lcout => \POWERLED.un1_dutycycle_53_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__29994\,
            in1 => \N__23115\,
            in2 => \N__19270\,
            in3 => \N__21481\,
            lcout => \POWERLED.dutycycleZ1Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34085\,
            ce => 'H',
            sr => \N__23697\
        );

    \POWERLED.dutycycle_RNI_13_9_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__27054\,
            in1 => \N__20771\,
            in2 => \N__21121\,
            in3 => \N__21775\,
            lcout => \POWERLED.dutycycle_RNI_13Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI03FP9_14_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__19266\,
            in1 => \N__29984\,
            in2 => \N__23116\,
            in3 => \N__21480\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__21890\,
            in1 => \_gnd_net_\,
            in2 => \N__19258\,
            in3 => \N__21433\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_9_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110100"
        )
    port map (
            in0 => \N__19255\,
            in1 => \N__19249\,
            in2 => \N__19243\,
            in3 => \N__19236\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19240\,
            in3 => \N__25341\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_4_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20963\,
            in1 => \N__21888\,
            in2 => \N__21804\,
            in3 => \N__27053\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI4J2O7_1_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__23143\,
            in1 => \N__19363\,
            in2 => \N__26768\,
            in3 => \N__29780\,
            lcout => \POWERLED.dutycycle_en_7\,
            ltout => \POWERLED.dutycycle_en_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__29992\,
            in1 => \N__19333\,
            in2 => \N__19219\,
            in3 => \N__21583\,
            lcout => \POWERLED.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33998\,
            ce => 'H',
            sr => \N__23668\
        );

    \POWERLED.dutycycle_9_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__19354\,
            in1 => \N__29993\,
            in2 => \N__19348\,
            in3 => \N__20695\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33998\,
            ce => 'H',
            sr => \N__23668\
        );

    \POWERLED.func_state_RNI2O4A1_0_1_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__30049\,
            in1 => \N__23173\,
            in2 => \_gnd_net_\,
            in3 => \N__21386\,
            lcout => \POWERLED.un1_clk_100khz_39_and_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_9_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__23172\,
            in1 => \N__30048\,
            in2 => \_gnd_net_\,
            in3 => \N__20773\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_30_and_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4J2O7_9_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__29779\,
            in1 => \N__26755\,
            in2 => \N__19357\,
            in3 => \N__23142\,
            lcout => \POWERLED.dutycycle_RNI4J2O7Z0Z_9\,
            ltout => \POWERLED.dutycycle_RNI4J2O7Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI880A9_9_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__19344\,
            in1 => \N__29990\,
            in2 => \N__19336\,
            in3 => \N__20694\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQPBP9_11_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__29991\,
            in1 => \N__19332\,
            in2 => \N__19324\,
            in3 => \N__21582\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILOQ6A_13_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__19485\,
            in1 => \N__29988\,
            in2 => \N__19504\,
            in3 => \N__21492\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_9_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21066\,
            in1 => \N__21359\,
            in2 => \_gnd_net_\,
            in3 => \N__20763\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_13_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__19313\,
            in1 => \N__23266\,
            in2 => \N__19276\,
            in3 => \N__21528\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_13_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__19452\,
            in1 => \N__19476\,
            in2 => \N__19273\,
            in3 => \N__21361\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__19500\,
            in1 => \N__29989\,
            in2 => \N__19489\,
            in3 => \N__21493\,
            lcout => \POWERLED.dutycycleZ1Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34086\,
            ce => 'H',
            sr => \N__23646\
        );

    \POWERLED.dutycycle_RNI_12_9_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21067\,
            in1 => \N__21360\,
            in2 => \N__21806\,
            in3 => \N__20764\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_12Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_9_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__19477\,
            in1 => \_gnd_net_\,
            in2 => \N__19462\,
            in3 => \N__19451\,
            lcout => \POWERLED.dutycycle_RNI_15Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_9_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__21065\,
            in1 => \N__20762\,
            in2 => \N__27145\,
            in3 => \N__21358\,
            lcout => \POWERLED.dutycycle_RNI_11Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22357\,
            in2 => \N__21301\,
            in3 => \N__22129\,
            lcout => \POWERLED.m18_e_0\,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19438\,
            in2 => \N__22376\,
            in3 => \N__19423\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23786\,
            in2 => \N__19420\,
            in3 => \N__19405\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19402\,
            in2 => \N__23796\,
            in3 => \N__19366\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19744\,
            in2 => \N__19728\,
            in3 => \N__19690\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26595\,
            in2 => \N__19687\,
            in3 => \N__19648\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19645\,
            in2 => \N__26605\,
            in3 => \N__19609\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21939\,
            in2 => \N__19606\,
            in3 => \N__19591\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19588\,
            in2 => \N__21449\,
            in3 => \N__19576\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23269\,
            in2 => \N__19573\,
            in3 => \N__19537\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19534\,
            in2 => \N__21562\,
            in3 => \N__19522\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25366\,
            in2 => \N__19519\,
            in3 => \N__19507\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25422\,
            in2 => \N__19921\,
            in3 => \N__19909\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21551\,
            in2 => \N__19906\,
            in3 => \N__19891\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19888\,
            in2 => \N__25377\,
            in3 => \N__19861\,
            lcout => \POWERLED.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25285\,
            in2 => \N__25431\,
            in3 => \N__19840\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25426\,
            in2 => \N__19804\,
            in3 => \N__19822\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19819\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25365\,
            in2 => \_gnd_net_\,
            in3 => \N__25305\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19795\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19767\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILP0F_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__31132\,
            in1 => \N__23908\,
            in2 => \N__20035\,
            in3 => \N__20017\,
            lcout => \POWERLED.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_9_5_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20970\,
            in2 => \_gnd_net_\,
            in3 => \N__21953\,
            lcout => \POWERLED.g3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_3_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21139\,
            in1 => \N__21314\,
            in2 => \N__19948\,
            in3 => \N__21809\,
            lcout => OPEN,
            ltout => \POWERLED.g0_4_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__22378\,
            in1 => \N__20008\,
            in2 => \N__19993\,
            in3 => \N__22143\,
            lcout => \POWERLED.N_398_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19989\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_10_5_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21808\,
            in1 => \N__22142\,
            in2 => \N__21316\,
            in3 => \N__21138\,
            lcout => OPEN,
            ltout => \POWERLED.g3_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_8_5_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19960\,
            in1 => \N__22377\,
            in2 => \N__19954\,
            in3 => \N__27154\,
            lcout => OPEN,
            ltout => \POWERLED.g3_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_7_5_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__27430\,
            in1 => \N__32944\,
            in2 => \N__19951\,
            in3 => \N__19944\,
            lcout => \POWERLED.un2_count_clk_17_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20073\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20211\,
            lcout => \POWERLED.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20139\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22460\,
            lcout => \POWERLED.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20077\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20300\,
            in2 => \N__20056\,
            in3 => \N__20047\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20044\,
            in2 => \N__20305\,
            in3 => \N__20038\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20374\,
            in2 => \N__20329\,
            in3 => \N__20368\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20328\,
            in2 => \N__20365\,
            in3 => \N__20356\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22213\,
            in1 => \N__20304\,
            in2 => \N__20353\,
            in3 => \N__20344\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20341\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20335\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => \POWERLED.mult1_un145_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20332\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20324\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20283\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20250\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22717\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33853\,
            ce => \N__27844\,
            sr => \N__28226\
        );

    \PCH_PWRGD.count_RNIS94O4_13_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20391\,
            in1 => \N__22763\,
            in2 => \_gnd_net_\,
            in3 => \N__27807\,
            lcout => \PCH_PWRGD.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22765\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33853\,
            ce => \N__27844\,
            sr => \N__28226\
        );

    \PCH_PWRGD.count_RNI0G6O4_15_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22716\,
            in1 => \N__20398\,
            in2 => \_gnd_net_\,
            in3 => \N__27808\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => \PCH_PWRGD.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIS94O4_0_13_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__27809\,
            in1 => \N__20392\,
            in2 => \N__20383\,
            in3 => \N__22764\,
            lcout => \PCH_PWRGD.count_1_i_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNIAKA42_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__27702\,
            in1 => \N__22659\,
            in2 => \N__22675\,
            in3 => \N__28225\,
            lcout => \PCH_PWRGD.count_rst_10\,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISVPK4_4_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27810\,
            in1 => \_gnd_net_\,
            in2 => \N__20380\,
            in3 => \N__24159\,
            lcout => \PCH_PWRGD.un2_count_1_axb_4\,
            ltout => \PCH_PWRGD.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__27703\,
            in1 => \N__28227\,
            in2 => \N__20377\,
            in3 => \N__22660\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33853\,
            ce => \N__27844\,
            sr => \N__28226\
        );

    \PCH_PWRGD.count_14_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22741\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28224\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33996\,
            ce => \N__27834\,
            sr => \N__28243\
        );

    \PCH_PWRGD.count_RNIOPNK4_2_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20454\,
            in1 => \N__27833\,
            in2 => \_gnd_net_\,
            in3 => \N__22523\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_2_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33996\,
            ce => \N__27834\,
            sr => \N__28243\
        );

    \PCH_PWRGD.count_RNIUC5O4_14_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__28223\,
            in1 => \N__22740\,
            in2 => \N__20464\,
            in3 => \N__27832\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => \PCH_PWRGD.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOPNK4_0_2_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__22524\,
            in1 => \N__20455\,
            in2 => \N__20446\,
            in3 => \N__27811\,
            lcout => \PCH_PWRGD.count_1_i_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_12_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33996\,
            ce => \N__27834\,
            sr => \N__28243\
        );

    \PCH_PWRGD.count_RNIQ63O4_12_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20443\,
            in1 => \N__22782\,
            in2 => \_gnd_net_\,
            in3 => \N__27831\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_0_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22692\,
            in2 => \_gnd_net_\,
            in3 => \N__22707\,
            lcout => \RSMRST_PWRGD.m4_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIKA9Q3_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__24710\,
            in1 => \N__20416\,
            in2 => \N__30811\,
            in3 => \N__20406\,
            lcout => \PCH_PWRGD_delayed_vccin_ok\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28278\,
            in2 => \N__31267\,
            in3 => \N__28300\,
            lcout => \PCH_PWRGD.N_250_0\,
            ltout => \PCH_PWRGD.N_250_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__30807\,
            in1 => \N__20407\,
            in2 => \N__20410\,
            in3 => \N__24711\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI2UUH1_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28299\,
            in1 => \N__31263\,
            in2 => \_gnd_net_\,
            in3 => \N__28384\,
            lcout => \PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI39MT5_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__20472\,
            in1 => \N__29807\,
            in2 => \N__20515\,
            in3 => \N__20524\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => \POWERLED.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNII3LM3_0_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__26715\,
            in1 => \N__31158\,
            in2 => \N__20527\,
            in3 => \N__21327\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => \POWERLED.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__20473\,
            in1 => \N__20514\,
            in2 => \N__20518\,
            in3 => \N__29809\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33997\,
            ce => 'H',
            sr => \N__23669\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101011111"
        )
    port map (
            in0 => \N__20626\,
            in1 => \N__26164\,
            in2 => \N__25027\,
            in3 => \N__29332\,
            lcout => \POWERLED.dutycycle_1_0_1\,
            ltout => \POWERLED.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__20497\,
            in1 => \N__20485\,
            in2 => \N__20500\,
            in3 => \N__29810\,
            lcout => \POWERLED.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33997\,
            ce => 'H',
            sr => \N__23669\
        );

    \POWERLED.dutycycle_RNII3LM3_1_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__26716\,
            in1 => \N__31159\,
            in2 => \N__22106\,
            in3 => \N__21328\,
            lcout => \POWERLED.dutycycle_eena_0\,
            ltout => \POWERLED.dutycycle_eena_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI7KKU5_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__20491\,
            in1 => \N__20484\,
            in2 => \N__20476\,
            in3 => \N__29808\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_0_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110101111"
        )
    port map (
            in0 => \N__22322\,
            in1 => \N__26163\,
            in2 => \N__25026\,
            in3 => \N__29331\,
            lcout => \POWERLED.dutycycle_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNISKPU6_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__24282\,
            in1 => \N__29985\,
            in2 => \N__26092\,
            in3 => \N__29772\,
            lcout => \POWERLED.func_state_RNISKPU6Z0Z_0\,
            ltout => \POWERLED.func_state_RNISKPU6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIVAIU9_13_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20608\,
            in1 => \_gnd_net_\,
            in2 => \N__20611\,
            in3 => \N__20599\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20607\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34293\,
            ce => \N__25557\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20577\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34293\,
            ce => \N__25557\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20593\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34293\,
            ce => \N__25557\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI1EJU9_14_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20592\,
            in1 => \N__20584\,
            in2 => \_gnd_net_\,
            in3 => \N__25517\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI3HKU9_15_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25558\,
            in1 => \N__20578\,
            in2 => \_gnd_net_\,
            in3 => \N__20566\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => \POWERLED.count_offZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20554\,
            in1 => \N__22839\,
            in2 => \N__20542\,
            in3 => \N__20539\,
            lcout => \POWERLED.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_3_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21299\,
            in1 => \N__21807\,
            in2 => \N__20647\,
            in3 => \N__27423\,
            lcout => \POWERLED.dutycycle_RNI_10Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__23982\,
            in1 => \N__20665\,
            in2 => \N__29806\,
            in3 => \N__22882\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34084\,
            ce => 'H',
            sr => \N__23695\
        );

    \POWERLED.dutycycle_RNIEP8SA_6_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__20664\,
            in1 => \N__29759\,
            in2 => \N__23983\,
            in3 => \N__22881\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => \POWERLED.dutycycleZ1Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22094\,
            in2 => \N__20653\,
            in3 => \N__22343\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_0\,
            ltout => \POWERLED.dutycycle_RNI_5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20650\,
            in3 => \N__26579\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32969\,
            in1 => \N__22093\,
            in2 => \_gnd_net_\,
            in3 => \N__22342\,
            lcout => \POWERLED.un1_dutycycle_96_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__32971\,
            in1 => \N__27424\,
            in2 => \N__20638\,
            in3 => \N__23881\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_3_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26239\,
            in2 => \N__20629\,
            in3 => \N__26476\,
            lcout => \POWERLED.un1_dutycycle_172_m3s4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__22086\,
            in1 => \_gnd_net_\,
            in2 => \N__22356\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23005\,
            in2 => \N__22112\,
            in3 => \N__20617\,
            lcout => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23009\,
            in2 => \N__23790\,
            in3 => \N__20614\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI765B1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29944\,
            in1 => \N__23006\,
            in2 => \N__21315\,
            in3 => \N__21169\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI765BZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI886B1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29983\,
            in1 => \N__23010\,
            in2 => \N__21813\,
            in3 => \N__21148\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI886BZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23007\,
            in2 => \N__26600\,
            in3 => \N__21145\,
            lcout => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23011\,
            in2 => \N__27078\,
            in3 => \N__21142\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4A1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29943\,
            in1 => \N__23008\,
            in2 => \N__21123\,
            in3 => \N__20974\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4AZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNICGAB1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29916\,
            in1 => \N__23002\,
            in2 => \N__20962\,
            in3 => \N__20818\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNICGABZ0Z1\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23012\,
            in2 => \N__20774\,
            in3 => \N__20686\,
            lcout => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCB1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29917\,
            in1 => \N__23003\,
            in2 => \N__21954\,
            in3 => \N__20668\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCBZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23013\,
            in2 => \N__21438\,
            in3 => \N__21574\,
            lcout => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23004\,
            in2 => \N__23229\,
            in3 => \N__21571\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23014\,
            in2 => \N__21547\,
            in3 => \N__21484\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23001\,
            in2 => \N__25370\,
            in3 => \N__21469\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__25427\,
            in1 => \_gnd_net_\,
            in2 => \N__27411\,
            in3 => \N__21466\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__24233\,
            in1 => \N__21621\,
            in2 => \N__26156\,
            in3 => \N__24246\,
            lcout => \POWERLED.N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21439\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_2_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111011101"
        )
    port map (
            in0 => \N__25019\,
            in1 => \N__32956\,
            in2 => \N__24235\,
            in3 => \N__21620\,
            lcout => \POWERLED.dutycycle_RNI2O4A1_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIA02P1_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__23346\,
            in1 => \N__26212\,
            in2 => \_gnd_net_\,
            in3 => \N__21651\,
            lcout => \POWERLED.N_115_f0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_6_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26594\,
            in1 => \N__29426\,
            in2 => \N__24082\,
            in3 => \N__27069\,
            lcout => \POWERLED.N_366\,
            ltout => \POWERLED.N_366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_6_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29914\,
            in2 => \N__21640\,
            in3 => \N__24234\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI2O4A1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI4G9K2_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27412\,
            in2 => \N__21637\,
            in3 => \N__21634\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI68EU3_1_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__29425\,
            in1 => \N__29913\,
            in2 => \N__21628\,
            in3 => \N__26470\,
            lcout => \POWERLED.func_state_RNI68EU3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_0_o2_0_6_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__29061\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21965\,
            lcout => \POWERLED.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24228\,
            in1 => \N__21625\,
            in2 => \_gnd_net_\,
            in3 => \N__26151\,
            lcout => \POWERLED.func_state_RNI_0Z0Z_0\,
            ltout => \POWERLED.func_state_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28962\,
            in2 => \N__21604\,
            in3 => \N__31116\,
            lcout => \POWERLED.func_state_RNIOGRSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__21967\,
            in1 => \_gnd_net_\,
            in2 => \N__25123\,
            in3 => \_gnd_net_\,
            lcout => \SUSWARN_N_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIT69J5_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__25860\,
            in1 => \N__31115\,
            in2 => \_gnd_net_\,
            in3 => \N__21601\,
            lcout => \POWERLED.func_state_RNIT69J5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI98TE_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__21595\,
            in1 => \N__29474\,
            in2 => \N__27348\,
            in3 => \N__29318\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_0_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI919H1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111001111"
        )
    port map (
            in0 => \N__29062\,
            in1 => \N__27335\,
            in2 => \N__21970\,
            in3 => \N__21966\,
            lcout => \POWERLED.un1_dutycycle_94_cry_4_c_RNI919HZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_4_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21950\,
            in1 => \N__21820\,
            in2 => \N__21814\,
            in3 => \N__27140\,
            lcout => \POWERLED.m18_e_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_eena_14_0_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__28901\,
            in1 => \N__26404\,
            in2 => \N__27339\,
            in3 => \N__29712\,
            lcout => \POWERLED.dutycycle_eena_14_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100111111"
        )
    port map (
            in0 => \N__29459\,
            in1 => \N__23757\,
            in2 => \N__26249\,
            in3 => \N__29995\,
            lcout => \POWERLED.un1_dutycycle_172_m1_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_rep1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23534\,
            in2 => \_gnd_net_\,
            in3 => \N__25117\,
            lcout => \SUSWARN_N_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_m2_0_a2_iso_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27315\,
            in1 => \N__23473\,
            in2 => \N__26411\,
            in3 => \N__30574\,
            lcout => \POWERLED.func_m2_0_a2_isoZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIVR902_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34565\,
            in1 => \N__21661\,
            in2 => \_gnd_net_\,
            in3 => \N__30190\,
            lcout => \POWERLED.dutycycle_1_0_5\,
            ltout => \POWERLED.dutycycle_1_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIBFCJ3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__23535\,
            in1 => \N__25118\,
            in2 => \N__21655\,
            in3 => \N__26210\,
            lcout => \POWERLED.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJ2BQ2_2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__26682\,
            in1 => \N__26209\,
            in2 => \N__21994\,
            in3 => \N__21652\,
            lcout => \POWERLED.dutycycle_eena_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_155_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23536\,
            in3 => \N__25110\,
            lcout => \G_155\,
            ltout => \G_155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJDU46_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__22021\,
            in1 => \N__22002\,
            in2 => \N__22024\,
            in3 => \N__22014\,
            lcout => \POWERLED.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIFRMD2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__21976\,
            in1 => \N__29469\,
            in2 => \N__26947\,
            in3 => \N__29316\,
            lcout => \POWERLED.N_73\,
            ltout => \POWERLED.N_73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__29711\,
            in1 => \N__22015\,
            in2 => \N__22006\,
            in3 => \N__22003\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34224\,
            ce => 'H',
            sr => \N__23615\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILP0F_2_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001000"
        )
    port map (
            in0 => \N__29317\,
            in1 => \N__31120\,
            in2 => \N__29481\,
            in3 => \N__23759\,
            lcout => \POWERLED.N_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__30238\,
            in1 => \N__21985\,
            in2 => \N__31154\,
            in3 => \N__29315\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOBHB2_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29458\,
            in2 => \N__26001\,
            in3 => \N__26942\,
            lcout => \POWERLED.func_state_1_m2_am_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__23875\,
            in1 => \N__23761\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_331\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22267\,
            in2 => \N__22179\,
            in3 => \N__22261\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22175\,
            in2 => \N__22258\,
            in3 => \N__22249\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22246\,
            in2 => \N__22223\,
            in3 => \N__22240\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22237\,
            in2 => \N__22224\,
            in3 => \N__22192\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__22189\,
            in2 => \N__22180\,
            in3 => \N__22162\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22159\,
            in2 => \_gnd_net_\,
            in3 => \N__22153\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => \POWERLED.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22150\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22144\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22433\,
            in2 => \N__22510\,
            in3 => \N__22495\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22492\,
            in2 => \N__22438\,
            in3 => \N__22486\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22461\,
            in2 => \N__22483\,
            in3 => \N__22474\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22471\,
            in2 => \N__22465\,
            in3 => \N__22441\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22600\,
            in1 => \N__22437\,
            in2 => \N__22423\,
            in3 => \N__22414\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22405\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => \POWERLED.mult1_un159_sum_s_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22402\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22366\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22580\,
            in2 => \N__22282\,
            in3 => \N__22601\,
            lcout => \G_2078\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22627\,
            in2 => \N__22585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22602\,
            in2 => \N__22621\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22612\,
            in2 => \N__22606\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22584\,
            in2 => \N__22570\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__22561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22555\,
            lcout => \POWERLED.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_9_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30612\,
            in2 => \_gnd_net_\,
            in3 => \N__25122\,
            lcout => \G_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27605\,
            in2 => \N__27628\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNI8G842_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28218\,
            in1 => \N__22531\,
            in2 => \_gnd_net_\,
            in3 => \N__22513\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24140\,
            in2 => \_gnd_net_\,
            in3 => \N__22678\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22671\,
            in2 => \_gnd_net_\,
            in3 => \N__22651\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27973\,
            in2 => \_gnd_net_\,
            in3 => \N__22648\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24484\,
            in2 => \_gnd_net_\,
            in3 => \N__22645\,
            lcout => \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28009\,
            in3 => \N__22642\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27464\,
            in3 => \N__22639\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27525\,
            in2 => \_gnd_net_\,
            in3 => \N__22636\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIG0H42_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28204\,
            in1 => \N__24352\,
            in2 => \_gnd_net_\,
            in3 => \N__22633\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27898\,
            in3 => \N__22630\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNIP94V1_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28205\,
            in1 => \N__24438\,
            in2 => \_gnd_net_\,
            in3 => \N__22774\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIQB5V1_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28222\,
            in1 => \N__22771\,
            in2 => \_gnd_net_\,
            in3 => \N__22750\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22747\,
            in2 => \_gnd_net_\,
            in3 => \N__22729\,
            lcout => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNISF7V1_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__22726\,
            in1 => \N__28206\,
            in2 => \_gnd_net_\,
            in3 => \N__22720\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIHNMD2_1_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__28203\,
            in1 => \N__28357\,
            in2 => \_gnd_net_\,
            in3 => \N__29827\,
            lcout => \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34858\,
            in1 => \N__24742\,
            in2 => \N__24805\,
            in3 => \N__24804\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34851\,
            in1 => \N__22708\,
            in2 => \_gnd_net_\,
            in3 => \N__22696\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_2_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34859\,
            in1 => \N__22693\,
            in2 => \_gnd_net_\,
            in3 => \N__22681\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34852\,
            in1 => \N__24520\,
            in2 => \_gnd_net_\,
            in3 => \N__22810\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_4_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34860\,
            in1 => \N__24631\,
            in2 => \_gnd_net_\,
            in3 => \N__22807\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_5_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34853\,
            in1 => \N__24559\,
            in2 => \_gnd_net_\,
            in3 => \N__22804\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_6_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34861\,
            in1 => \N__24547\,
            in2 => \_gnd_net_\,
            in3 => \N__22801\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_7_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34854\,
            in1 => \N__24534\,
            in2 => \_gnd_net_\,
            in3 => \N__22798\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__34144\,
            ce => 'H',
            sr => \N__25165\
        );

    \RSMRST_PWRGD.count_8_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34850\,
            in1 => \N__24643\,
            in2 => \_gnd_net_\,
            in3 => \N__22795\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.count_9_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34846\,
            in1 => \N__24655\,
            in2 => \_gnd_net_\,
            in3 => \N__22792\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.count_10_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34847\,
            in1 => \N__24781\,
            in2 => \_gnd_net_\,
            in3 => \N__22789\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.count_11_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34844\,
            in1 => \N__24616\,
            in2 => \_gnd_net_\,
            in3 => \N__22786\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.count_12_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34848\,
            in1 => \N__24577\,
            in2 => \_gnd_net_\,
            in3 => \N__22867\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.count_13_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34845\,
            in1 => \N__24769\,
            in2 => \_gnd_net_\,
            in3 => \N__22864\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.count_14_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34849\,
            in1 => \N__24604\,
            in2 => \_gnd_net_\,
            in3 => \N__22861\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__34080\,
            ce => 'H',
            sr => \N__25173\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34557\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24591\,
            in2 => \_gnd_net_\,
            in3 => \N__22858\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34324\,
            ce => \N__25135\,
            sr => \N__25180\
        );

    \POWERLED.count_off_RNIBQDB2_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22837\,
            lcout => OPEN,
            ltout => \POWERLED.count_off_RNIBQDB2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI2KLI9_0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22816\,
            in2 => \N__22855\,
            in3 => \N__25496\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => \POWERLED.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22852\,
            in3 => \N__22941\,
            lcout => \POWERLED.count_off_RNIZ0Z_1\,
            ltout => \POWERLED.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22849\,
            in3 => \N__26864\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34233\,
            ce => \N__25583\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22838\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34233\,
            ce => \N__25583\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI3LLI9_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22960\,
            in1 => \N__25495\,
            in2 => \N__22954\,
            in3 => \N__26861\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => \POWERLED.count_offZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__25734\,
            in1 => \N__25668\,
            in2 => \N__22927\,
            in3 => \N__25455\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_10_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22924\,
            in1 => \N__22918\,
            in2 => \N__22906\,
            in3 => \N__22903\,
            lcout => \POWERLED.count_off_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIRGL41_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111101"
        )
    port map (
            in0 => \N__31026\,
            in1 => \N__29382\,
            in2 => \N__23089\,
            in3 => \N__22891\,
            lcout => OPEN,
            ltout => \POWERLED.N_220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI4L823_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__30149\,
            in1 => \N__26693\,
            in2 => \N__22885\,
            in3 => \N__29305\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_0_0_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__31027\,
            in1 => \N__29383\,
            in2 => \N__29573\,
            in3 => \N__28984\,
            lcout => OPEN,
            ltout => \POWERLED.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHGMD3_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__23026\,
            in1 => \N__26694\,
            in2 => \N__22870\,
            in3 => \N__29306\,
            lcout => \POWERLED.func_state_1_ss0_i_0_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26155\,
            lcout => \POWERLED.N_2216_i\,
            ltout => \POWERLED.N_2216_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJ9IE1_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001101"
        )
    port map (
            in0 => \N__29333\,
            in1 => \N__26692\,
            in2 => \N__23095\,
            in3 => \N__23848\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m2s2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIN2PE3_1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__29307\,
            in1 => \N__25186\,
            in2 => \N__23092\,
            in3 => \N__23025\,
            lcout => \POWERLED.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIMJCH1_10_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__28983\,
            in1 => \N__23088\,
            in2 => \N__29574\,
            in3 => \N__31028\,
            lcout => \POWERLED.N_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_1_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29915\,
            in1 => \N__32952\,
            in2 => \_gnd_net_\,
            in3 => \N__30037\,
            lcout => \POWERLED.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.slp_s3n_signal_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26969\,
            lcout => slp_s3n_signal,
            ltout => \slp_s3n_signal_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__28982\,
            in1 => \_gnd_net_\,
            in2 => \N__23029\,
            in3 => \N__30465\,
            lcout => \POWERLED.N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_m1_0_a2_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27347\,
            in1 => \N__29040\,
            in2 => \_gnd_net_\,
            in3 => \N__26070\,
            lcout => \POWERLED.un1_N_3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29392\,
            in3 => \N__29301\,
            lcout => \POWERLED.func_state_RNIZ0Z_1\,
            ltout => \POWERLED.func_state_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_8_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23017\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIET094_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25817\,
            in1 => \N__26211\,
            in2 => \N__23457\,
            in3 => \N__23345\,
            lcout => \POWERLED.N_399_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIV0AS_1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__26069\,
            in2 => \N__29330\,
            in3 => \N__29371\,
            lcout => \POWERLED.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4J2O7_12_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__29744\,
            in1 => \N__26678\,
            in2 => \N__23136\,
            in3 => \N__23179\,
            lcout => \POWERLED.dutycycle_en_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__23287\,
            in1 => \N__23311\,
            in2 => \N__23302\,
            in3 => \N__29939\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34449\,
            ce => 'H',
            sr => \N__23664\
        );

    \POWERLED.func_state_RNI2O4A1_1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24991\,
            in2 => \_gnd_net_\,
            in3 => \N__29202\,
            lcout => \POWERLED.func_state_RNI2O4A1Z0Z_1\,
            ltout => \POWERLED.func_state_RNI2O4A1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_1_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23314\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.func_state_RNI2O4A1_1Z0Z_1\,
            ltout => \POWERLED.func_state_RNI2O4A1_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNISSCP9_12_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23310\,
            in1 => \N__23298\,
            in2 => \N__23290\,
            in3 => \N__23286\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => \POWERLED.dutycycleZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_12_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__30038\,
            in1 => \_gnd_net_\,
            in2 => \N__23182\,
            in3 => \N__23162\,
            lcout => \POWERLED.un1_clk_100khz_42_and_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_14_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__30050\,
            in1 => \N__25375\,
            in2 => \_gnd_net_\,
            in3 => \N__23166\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_47_and_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4J2O7_14_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__26677\,
            in1 => \N__29743\,
            in2 => \N__23146\,
            in3 => \N__23129\,
            lcout => \POWERLED.dutycycle_en_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_3_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__27420\,
            in1 => \N__23494\,
            in2 => \N__32970\,
            in3 => \N__23479\,
            lcout => \POWERLED.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__23392\,
            in1 => \N__30165\,
            in2 => \N__25903\,
            in3 => \N__23398\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_m2_0_a2_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29060\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28979\,
            lcout => \POWERLED.func_m2_0_a2Z0Z_0\,
            ltout => \POWERLED.func_m2_0_a2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_m2_0_a2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26386\,
            in1 => \N__27319\,
            in2 => \N__23467\,
            in3 => \N__23532\,
            lcout => \POWERLED.func_N_5_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2O4A1_0_10_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29896\,
            in2 => \_gnd_net_\,
            in3 => \N__32951\,
            lcout => \POWERLED.count_clk_RNI2O4A1_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI91IA4_0_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010001"
        )
    port map (
            in0 => \N__25996\,
            in1 => \N__27419\,
            in2 => \N__25963\,
            in3 => \N__29588\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNI91IA4_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI4CHA7_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25939\,
            in1 => \_gnd_net_\,
            in2 => \N__23401\,
            in3 => \N__23503\,
            lcout => \POWERLED.func_state_1_m2_0\,
            ltout => \POWERLED.func_state_1_m2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIA20K9_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23391\,
            in1 => \N__30164\,
            in2 => \N__23383\,
            in3 => \N__25896\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE1QU7_5_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101010011"
        )
    port map (
            in0 => \N__23931\,
            in1 => \N__23829\,
            in2 => \N__26308\,
            in3 => \N__26199\,
            lcout => OPEN,
            ltout => \POWERLED.g0_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILMBVD_5_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001010"
        )
    port map (
            in0 => \N__23887\,
            in1 => \N__29678\,
            in2 => \N__23713\,
            in3 => \N__26304\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_fb_15_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1DAA11_5_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23542\,
            in1 => \N__23707\,
            in2 => \N__23710\,
            in3 => \N__23566\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBQG35_5_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__23806\,
            in1 => \N__23577\,
            in2 => \N__24019\,
            in3 => \N__23828\,
            lcout => \POWERLED.dutycycle_fb_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__23576\,
            in1 => \N__26689\,
            in2 => \_gnd_net_\,
            in3 => \N__23992\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_en_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__26690\,
            in1 => \N__23826\,
            in2 => \N__23701\,
            in3 => \N__23930\,
            lcout => \POWERLED.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34458\,
            ce => 'H',
            sr => \N__23616\
        );

    \POWERLED.dutycycle_RNIN2958_5_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__23578\,
            in1 => \N__24018\,
            in2 => \N__23917\,
            in3 => \N__26691\,
            lcout => \POWERLED.dutycycle_fb_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIAP426_5_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__23557\,
            in1 => \N__23551\,
            in2 => \N__24040\,
            in3 => \N__23827\,
            lcout => \POWERLED.dutycycle_fb_15_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_0_2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23533\,
            in1 => \N__28941\,
            in2 => \N__29068\,
            in3 => \N__31163\,
            lcout => \POWERLED.N_340\,
            ltout => \POWERLED.N_340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRAVV2_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__26002\,
            in1 => \N__29589\,
            in2 => \N__23506\,
            in3 => \N__26113\,
            lcout => \POWERLED.func_state_RNIRAVV2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKLAF2_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24312\,
            in1 => \N__24052\,
            in2 => \N__31167\,
            in3 => \N__23932\,
            lcout => \POWERLED.dutycycle_fb_15_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_6_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__26545\,
            in1 => \N__23880\,
            in2 => \N__27144\,
            in3 => \N__24313\,
            lcout => \POWERLED.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILP0F_0_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__24331\,
            in1 => \N__23896\,
            in2 => \N__32967\,
            in3 => \N__31164\,
            lcout => \POWERLED.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24083\,
            in1 => \N__23879\,
            in2 => \_gnd_net_\,
            in3 => \N__27110\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_6_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24084\,
            in1 => \N__24217\,
            in2 => \N__27143\,
            in3 => \N__26516\,
            lcout => \POWERLED.func_state_1_m2s2_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8OIL_5_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24306\,
            in1 => \N__24051\,
            in2 => \N__23836\,
            in3 => \N__31147\,
            lcout => \POWERLED.dutycycle_fb_14_a4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNINH5P1_2_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001111"
        )
    port map (
            in0 => \N__23719\,
            in1 => \N__24292\,
            in2 => \N__31165\,
            in3 => \N__23758\,
            lcout => \POWERLED.dutycycle_RNINH5P1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_2_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30003\,
            in2 => \_gnd_net_\,
            in3 => \N__29460\,
            lcout => \POWERLED.count_off_1_sqmuxa\,
            ltout => \POWERLED.count_off_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4G9K2_5_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__26577\,
            in1 => \N__25018\,
            in2 => \N__24127\,
            in3 => \N__24124\,
            lcout => \POWERLED.dutycycle_RNI4G9K2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_6_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__24342\,
            in1 => \N__32963\,
            in2 => \_gnd_net_\,
            in3 => \N__26576\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_6\,
            ltout => \POWERLED.dutycycle_RNI_4Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32964\,
            in1 => \N__24118\,
            in2 => \N__24088\,
            in3 => \N__24085\,
            lcout => \POWERLED.dutycycle_RNI_8Z0Z_0\,
            ltout => \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_2_5_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__24036\,
            in1 => \N__24009\,
            in2 => \N__23998\,
            in3 => \N__31145\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNO_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_1_5_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31146\,
            in1 => \N__24305\,
            in2 => \N__23995\,
            in3 => \N__23938\,
            lcout => \POWERLED.N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_4_5_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__29479\,
            in1 => \N__29981\,
            in2 => \_gnd_net_\,
            in3 => \N__26474\,
            lcout => \POWERLED.g3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILG3T6_6_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__27001\,
            in1 => \N__26700\,
            in2 => \N__24265\,
            in3 => \N__24190\,
            lcout => \POWERLED.dutycycle_eena_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_5_5_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111000001111"
        )
    port map (
            in0 => \N__26250\,
            in1 => \N__26287\,
            in2 => \N__24184\,
            in3 => \N__23959\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_3_5_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__26475\,
            in1 => \N__23947\,
            in2 => \N__23941\,
            in3 => \N__26575\,
            lcout => \POWERLED.dutycycle_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_6_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__24346\,
            in1 => \N__24330\,
            in2 => \_gnd_net_\,
            in3 => \N__32965\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2O4A1_10_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29982\,
            in2 => \_gnd_net_\,
            in3 => \N__32966\,
            lcout => \POWERLED.count_clk_RNI2O4A1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__29313\,
            in1 => \N__29478\,
            in2 => \_gnd_net_\,
            in3 => \N__26574\,
            lcout => \POWERLED.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI88TE_0_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__24286\,
            in1 => \N__27277\,
            in2 => \_gnd_net_\,
            in3 => \N__26397\,
            lcout => \POWERLED.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMQ0F_1_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24253\,
            in1 => \N__30189\,
            in2 => \N__24229\,
            in3 => \N__29302\,
            lcout => \POWERLED.N_272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_6_5_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27264\,
            in1 => \N__28885\,
            in2 => \_gnd_net_\,
            in3 => \N__26387\,
            lcout => \POWERLED.dutycycle_N_3_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISVPK4_0_4_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__24172\,
            in1 => \N__24163\,
            in2 => \N__27858\,
            in3 => \N__24141\,
            lcout => \PCH_PWRGD.count_1_i_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNI9I942_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__27692\,
            in1 => \N__28208\,
            in2 => \N__24145\,
            in3 => \N__24387\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQSOK4_3_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27780\,
            in1 => \_gnd_net_\,
            in2 => \N__24148\,
            in3 => \N__24379\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => \PCH_PWRGD.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_3_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__27693\,
            in1 => \N__28210\,
            in2 => \N__24391\,
            in3 => \N__24388\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34055\,
            ce => \N__27845\,
            sr => \N__28228\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNIESE42_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__28207\,
            in1 => \N__27691\,
            in2 => \N__27465\,
            in3 => \N__24366\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI4CUK4_8_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24358\,
            in2 => \N__24373\,
            in3 => \N__27779\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => \PCH_PWRGD.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_8_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__28209\,
            in1 => \N__27694\,
            in2 => \N__24370\,
            in3 => \N__24367\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34055\,
            ce => \N__27845\,
            sr => \N__28228\
        );

    \PCH_PWRGD.count_9_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__27695\,
            in1 => \N__28211\,
            in2 => \N__27526\,
            in3 => \N__27501\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34055\,
            ce => \N__27845\,
            sr => \N__28228\
        );

    \PCH_PWRGD.count_10_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24465\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34197\,
            ce => \N__27838\,
            sr => \N__28217\
        );

    \PCH_PWRGD.count_6_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__24493\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28216\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34197\,
            ce => \N__27838\,
            sr => \N__28217\
        );

    \PCH_PWRGD.count_RNIFRFT4_10_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24477\,
            in1 => \N__24464\,
            in2 => \_gnd_net_\,
            in3 => \N__27802\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__24669\,
            in2 => \N__28240\,
            in3 => \N__27553\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34197\,
            ce => \N__27838\,
            sr => \N__28217\
        );

    \PCH_PWRGD.count_RNI06SK4_6_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__24502\,
            in1 => \N__24492\,
            in2 => \N__28239\,
            in3 => \N__27803\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => \PCH_PWRGD.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIFRFT4_0_10_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__27804\,
            in1 => \N__24478\,
            in2 => \N__24469\,
            in3 => \N__24466\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI3VBAE_2_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__24451\,
            in1 => \N__24442\,
            in2 => \N__24427\,
            in3 => \N__24424\,
            lcout => \PCH_PWRGD.count_1_i_a2_11_0\,
            ltout => \PCH_PWRGD.count_1_i_a2_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIM6A821_1_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__24679\,
            in1 => \N__28212\,
            in2 => \N__24412\,
            in3 => \N__27552\,
            lcout => \PCH_PWRGD.count_RNIM6A821Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNIO73V1_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__28166\,
            in1 => \N__27921\,
            in2 => \N__27905\,
            in3 => \N__27685\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIO32O4_11_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27871\,
            in2 => \N__24409\,
            in3 => \N__27805\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__30951\,
            in1 => \_gnd_net_\,
            in2 => \N__25234\,
            in3 => \N__25266\,
            lcout => OPEN,
            ltout => \N_253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_11_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__24818\,
            in1 => \N__34839\,
            in2 => \N__24406\,
            in3 => \N__25232\,
            lcout => \G_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI4EPO41_0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27806\,
            in1 => \N__24403\,
            in2 => \_gnd_net_\,
            in3 => \N__24397\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => \PCH_PWRGD.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI_0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24682\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2173_i\,
            ltout => \PCH_PWRGD.N_2173_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI63UG01_1_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24670\,
            in2 => \N__24658\,
            in3 => \N__27551\,
            lcout => \PCH_PWRGD.N_364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__25267\,
            in1 => \N__30950\,
            in2 => \N__24825\,
            in3 => \N__25233\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34069\,
            ce => \N__34687\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28376\,
            lcout => \PCH_PWRGD.N_2171_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_11_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24654\,
            in1 => \N__24642\,
            in2 => \N__25273\,
            in3 => \N__24630\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.m4_0_a2_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24565\,
            in1 => \N__24508\,
            in2 => \N__24619\,
            in3 => \N__24730\,
            lcout => \N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_10_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24615\,
            in1 => \N__24603\,
            in2 => \N__24592\,
            in3 => \N__24576\,
            lcout => \RSMRST_PWRGD.m4_0_a2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_9_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24558\,
            in1 => \N__24546\,
            in2 => \N__24535\,
            in3 => \N__24519\,
            lcout => \RSMRST_PWRGD.m4_0_a2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_12_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24780\,
            in1 => \N__24768\,
            in2 => \N__24757\,
            in3 => \N__24741\,
            lcout => \RSMRST_PWRGD.m4_0_a2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32172\,
            in1 => \N__31988\,
            in2 => \N__28557\,
            in3 => \N__31798\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24955\,
            in2 => \N__24724\,
            in3 => \N__31620\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__28333\,
            in1 => \N__28270\,
            in2 => \_gnd_net_\,
            in3 => \N__24720\,
            lcout => \PCH_PWRGD.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34294\,
            ce => \N__30778\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__24721\,
            in1 => \N__28271\,
            in2 => \_gnd_net_\,
            in3 => \N__28332\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.m4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI0EA52_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24694\,
            in2 => \N__24688\,
            in3 => \N__30531\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32166\,
            in1 => \N__31790\,
            in2 => \N__30850\,
            in3 => \N__31980\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31791\,
            in1 => \N__32167\,
            in2 => \N__28599\,
            in3 => \N__31981\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPM861_8_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24970\,
            in2 => \N__24685\,
            in3 => \N__31626\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31794\,
            in1 => \N__32171\,
            in2 => \N__28600\,
            in3 => \N__31984\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34210\,
            ce => \N__31631\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__32169\,
            in1 => \N__31795\,
            in2 => \N__31990\,
            in3 => \N__28578\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34210\,
            ce => \N__31631\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31792\,
            in1 => \N__32168\,
            in2 => \N__28579\,
            in3 => \N__31982\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIRP961_9_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24964\,
            in2 => \N__24958\,
            in3 => \N__31627\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31793\,
            in1 => \N__32170\,
            in2 => \N__28558\,
            in3 => \N__31983\,
            lcout => \VPP_VDDQ.count_2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34210\,
            ce => \N__31631\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24935\,
            in1 => \N__24901\,
            in2 => \N__24882\,
            in3 => \N__24855\,
            lcout => rsmrst_pwrgd_signal,
            ltout => \rsmrst_pwrgd_signal_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a3_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25208\,
            in2 => \N__24832\,
            in3 => \N__25269\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__25209\,
            in1 => \_gnd_net_\,
            in2 => \N__24829\,
            in3 => \N__24826\,
            lcout => \RSMRST_PWRGD_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34161\,
            ce => \N__34696\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__30941\,
            in1 => \N__25207\,
            in2 => \_gnd_net_\,
            in3 => \N__25268\,
            lcout => \RSMRST_PWRGD.N_254_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__25271\,
            in1 => \_gnd_net_\,
            in2 => \N__25221\,
            in3 => \N__30940\,
            lcout => \RSMRSTn_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34161\,
            ce => \N__34696\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30939\,
            in1 => \N__25210\,
            in2 => \_gnd_net_\,
            in3 => \N__25272\,
            lcout => \RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34161\,
            ce => \N__34696\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__25270\,
            in1 => \_gnd_net_\,
            in2 => \N__25220\,
            in3 => \N__30938\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34161\,
            ce => \N__34696\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIU2UT_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000000000"
        )
    port map (
            in0 => \N__26352\,
            in1 => \N__28960\,
            in2 => \N__31108\,
            in3 => \N__26617\,
            lcout => \POWERLED.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_en_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__28961\,
            in1 => \N__26351\,
            in2 => \N__27349\,
            in3 => \N__29758\,
            lcout => \POWERLED.func_state_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34840\,
            in2 => \_gnd_net_\,
            in3 => \N__25172\,
            lcout => \RSMRST_PWRGD.N_29_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_0_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26970\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30490\,
            in2 => \_gnd_net_\,
            in3 => \N__25121\,
            lcout => suswarn_n,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_m1_e_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27341\,
            in1 => \N__28959\,
            in2 => \_gnd_net_\,
            in3 => \N__26068\,
            lcout => \POWERLED.dutycycle_N_3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25789\,
            in2 => \N__32305\,
            in3 => \N__33318\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32304\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34332\,
            ce => \N__33332\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIVI1E_9_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25783\,
            in2 => \N__32284\,
            in3 => \N__33319\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32283\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34332\,
            ce => \N__33332\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI17P1A_5_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25777\,
            in1 => \N__25759\,
            in2 => \_gnd_net_\,
            in3 => \N__25569\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI3AQ1A_6_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25570\,
            in1 => \N__25708\,
            in2 => \_gnd_net_\,
            in3 => \N__25690\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIRTL1A_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25642\,
            in1 => \N__25624\,
            in2 => \_gnd_net_\,
            in3 => \N__25568\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_15_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__25435\,
            in1 => \N__25371\,
            in2 => \_gnd_net_\,
            in3 => \N__25306\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_1_2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28980\,
            in1 => \N__29051\,
            in2 => \_gnd_net_\,
            in3 => \N__31139\,
            lcout => \POWERLED.N_340_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__25895\,
            in1 => \N__25915\,
            in2 => \N__30188\,
            in3 => \N__25921\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_0_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__26074\,
            in1 => \N__28981\,
            in2 => \N__27334\,
            in3 => \N__30051\,
            lcout => \POWERLED.N_4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI91IA4_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__25997\,
            in1 => \N__27421\,
            in2 => \N__25962\,
            in3 => \N__29587\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNI91IA4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIKML48_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__26626\,
            in1 => \N__25938\,
            in2 => \N__25924\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.func_state_1_m2_1\,
            ltout => \POWERLED.func_state_1_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRD4EA_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25914\,
            in1 => \N__30159\,
            in2 => \N__25906\,
            in3 => \N__25894\,
            lcout => \POWERLED.func_state\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__30160\,
            in1 => \N__25848\,
            in2 => \_gnd_net_\,
            in3 => \N__29424\,
            lcout => \POWERLED.un1_func_state25_6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_7_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27422\,
            in2 => \_gnd_net_\,
            in3 => \N__32915\,
            lcout => \func_state_RNI_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_0_2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__26285\,
            in1 => \N__26295\,
            in2 => \_gnd_net_\,
            in3 => \N__26259\,
            lcout => OPEN,
            ltout => \N_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S3n_RNI75Q52_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27303\,
            in1 => \N__28909\,
            in2 => \N__25792\,
            in3 => \N__26469\,
            lcout => OPEN,
            ltout => \G_34_0_a4_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_RNIH76R4_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__26353\,
            in1 => \N__26218\,
            in2 => \N__26311\,
            in3 => \N__26422\,
            lcout => \POWERLED_un1_dutycycle_172_m3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_1_2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__26296\,
            in1 => \N__26286\,
            in2 => \N__26263\,
            in3 => \N__26468\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__26354\,
            in1 => \N__28908\,
            in2 => \_gnd_net_\,
            in3 => \N__27302\,
            lcout => \POWERLED.N_319_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26147\,
            in2 => \_gnd_net_\,
            in3 => \N__29223\,
            lcout => \POWERLED.func_state_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3VDK_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000000000"
        )
    port map (
            in0 => \N__30491\,
            in1 => \N__31133\,
            in2 => \N__26157\,
            in3 => \N__29626\,
            lcout => \POWERLED.N_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBVNS_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28755\,
            in1 => \N__32494\,
            in2 => \N__28827\,
            in3 => \N__29504\,
            lcout => \POWERLED.N_284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_2_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32496\,
            in1 => \N__28756\,
            in2 => \N__28820\,
            in3 => \N__29246\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_o_N_296_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__26107\,
            in1 => \N__26785\,
            in2 => \N__26098\,
            in3 => \N__29625\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__26815\,
            in1 => \N__27428\,
            in2 => \N__26095\,
            in3 => \N__29582\,
            lcout => \POWERLED.un1_func_state25_6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI0RLE1_8_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__26946\,
            in1 => \_gnd_net_\,
            in2 => \N__29593\,
            in3 => \N__32497\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBQDB2_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__26803\,
            in1 => \N__29115\,
            in2 => \N__26929\,
            in3 => \N__26926\,
            lcout => \POWERLED.func_state_RNIBQDB2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29116\,
            in1 => \N__26814\,
            in2 => \N__26802\,
            in3 => \N__32495\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_294_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBL3Q3_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111011"
        )
    port map (
            in0 => \N__29505\,
            in1 => \N__26779\,
            in2 => \N__26759\,
            in3 => \N__29583\,
            lcout => \POWERLED.func_state_RNIBL3Q3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_0_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__29303\,
            in1 => \N__31148\,
            in2 => \_gnd_net_\,
            in3 => \N__28957\,
            lcout => \POWERLED.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_9_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29451\,
            in2 => \_gnd_net_\,
            in3 => \N__29509\,
            lcout => \POWERLED.func_state_1_m2s2_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_5_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000101010"
        )
    port map (
            in0 => \N__26578\,
            in1 => \N__30004\,
            in2 => \N__29473\,
            in3 => \N__26456\,
            lcout => \N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__28956\,
            in1 => \N__26355\,
            in2 => \N__27333\,
            in3 => \N__29447\,
            lcout => \POWERLED.func_state_RNIBVNSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_0_1_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__27429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29066\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_a2_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8H551_6_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__28911\,
            in1 => \N__27265\,
            in2 => \N__27187\,
            in3 => \N__27163\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_a2_6_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRKB61_6_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__26981\,
            in1 => \_gnd_net_\,
            in2 => \N__27184\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_309_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPUGO_0_1_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__28912\,
            in1 => \N__26992\,
            in2 => \_gnd_net_\,
            in3 => \N__26982\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNIPUGO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI7N202_1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31149\,
            in1 => \_gnd_net_\,
            in2 => \N__27181\,
            in3 => \N__26953\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_o2_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI44JG4_6_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110111011"
        )
    port map (
            in0 => \N__27178\,
            in1 => \N__27172\,
            in2 => \N__27166\,
            in3 => \N__27162\,
            lcout => \POWERLED.N_145_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29304\,
            in2 => \_gnd_net_\,
            in3 => \N__29067\,
            lcout => \POWERLED.un1_clk_100khz_51_and_i_a2_5_0\,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPUGO_1_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__28913\,
            in1 => \N__29314\,
            in2 => \N__26986\,
            in3 => \N__26983\,
            lcout => \POWERLED.func_state_RNIPUGOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__30310\,
            in1 => \N__30260\,
            in2 => \_gnd_net_\,
            in3 => \N__30076\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34417\,
            ce => \N__34712\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_1_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28169\,
            in1 => \N__27624\,
            in2 => \_gnd_net_\,
            in3 => \N__27607\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33983\,
            ce => \N__27859\,
            sr => \N__28170\
        );

    \PCH_PWRGD.count_RNIVBR74_1_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27576\,
            in1 => \N__27850\,
            in2 => \_gnd_net_\,
            in3 => \N__27583\,
            lcout => \PCH_PWRGD.un2_count_1_axb_1\,
            ltout => \PCH_PWRGD.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIG3CN1_1_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__28168\,
            in1 => \_gnd_net_\,
            in2 => \N__27610\,
            in3 => \N__27606\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => \PCH_PWRGD.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIVBR74_0_1_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001000100"
        )
    port map (
            in0 => \N__27577\,
            in1 => \N__27909\,
            in2 => \N__27568\,
            in3 => \N__27852\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI34I6I_1_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27436\,
            in1 => \N__27565\,
            in2 => \N__27556\,
            in3 => \N__28030\,
            lcout => \PCH_PWRGD.count_1_i_a2_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI6FVK4_9_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27477\,
            in1 => \N__27484\,
            in2 => \_gnd_net_\,
            in3 => \N__27849\,
            lcout => \PCH_PWRGD.un2_count_1_axb_9\,
            ltout => \PCH_PWRGD.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNIFUF42_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__28167\,
            in1 => \N__27505\,
            in2 => \N__27487\,
            in3 => \N__27696\,
            lcout => \PCH_PWRGD.count_rst_5\,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI6FVK4_0_9_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__27478\,
            in1 => \N__27466\,
            in2 => \N__27439\,
            in3 => \N__27851\,
            lcout => \PCH_PWRGD.count_1_i_a2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI29TK4_7_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28039\,
            in1 => \N__27985\,
            in2 => \_gnd_net_\,
            in3 => \N__27820\,
            lcout => \PCH_PWRGD.un2_count_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNIDQD42_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__27701\,
            in1 => \N__28024\,
            in2 => \N__28235\,
            in3 => \N__28002\,
            lcout => \PCH_PWRGD.count_rst_7\,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI29TK4_0_7_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__27857\,
            in1 => \N__27984\,
            in2 => \N__28033\,
            in3 => \N__27965\,
            lcout => \PCH_PWRGD.count_1_i_a2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__27699\,
            in1 => \N__28023\,
            in2 => \N__28234\,
            in3 => \N__28001\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34275\,
            ce => \N__27856\,
            sr => \N__28241\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIBMB42_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__28083\,
            in1 => \N__27966\,
            in2 => \N__27952\,
            in3 => \N__27700\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIU2RK4_5_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27931\,
            in1 => \_gnd_net_\,
            in2 => \N__27976\,
            in3 => \N__27821\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => \PCH_PWRGD.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_5_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__27948\,
            in1 => \N__28193\,
            in2 => \N__27934\,
            in3 => \N__27698\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34275\,
            ce => \N__27856\,
            sr => \N__28241\
        );

    \PCH_PWRGD.count_11_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__27697\,
            in1 => \N__27925\,
            in2 => \N__27910\,
            in3 => \N__28242\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34275\,
            ce => \N__27856\,
            sr => \N__28241\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_i_a2_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28309\,
            in2 => \_gnd_net_\,
            in3 => \N__27670\,
            lcout => \G_1939\,
            ltout => \G_1939_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28387\,
            in3 => \N__28353\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34292\,
            ce => \N__30779\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_i_o3_0_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__31254\,
            in1 => \N__28290\,
            in2 => \_gnd_net_\,
            in3 => \N__28383\,
            lcout => \N_218\,
            ltout => \N_218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__28339\,
            in1 => \N__28326\,
            in2 => \N__28312\,
            in3 => \N__30575\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => \PCH_PWRGD.curr_state_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIVGBJ_0_1_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28303\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2190_i\,
            ltout => \PCH_PWRGD.N_2190_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIG3CN1_1_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__28279\,
            in1 => \N__31253\,
            in2 => \N__28246\,
            in3 => \N__30576\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__31777\,
            in1 => \N__32069\,
            in2 => \N__30411\,
            in3 => \N__31908\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34374\,
            ce => \N__30780\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__31907\,
            in1 => \N__30406\,
            in2 => \N__32111\,
            in3 => \N__31778\,
            lcout => \VPP_VDDQ.curr_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34374\,
            ce => \N__30780\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101110111"
        )
    port map (
            in0 => \N__31775\,
            in1 => \N__32068\,
            in2 => \N__30412\,
            in3 => \N__31909\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28048\,
            in2 => \N__28042\,
            in3 => \N__30547\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110011"
        )
    port map (
            in0 => \N__31774\,
            in1 => \N__30410\,
            in2 => \N__28417\,
            in3 => \N__32073\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28414\,
            in2 => \N__28408\,
            in3 => \N__30546\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31776\,
            in1 => \N__28444\,
            in2 => \N__28405\,
            in3 => \N__31906\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIF7361_3_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28486\,
            in2 => \N__28402\,
            in3 => \N__31549\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__31744\,
            in1 => \N__28473\,
            in2 => \N__31953\,
            in3 => \N__32086\,
            lcout => \VPP_VDDQ.count_2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34378\,
            ce => \N__31621\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32083\,
            in1 => \N__31901\,
            in2 => \N__28474\,
            in3 => \N__31742\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID4261_2_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31547\,
            in1 => \_gnd_net_\,
            in2 => \N__28399\,
            in3 => \N__28396\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => \VPP_VDDQ.count_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_2_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28621\,
            in1 => \N__31297\,
            in2 => \N__28390\,
            in3 => \N__28458\,
            lcout => \VPP_VDDQ.un9_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31743\,
            in1 => \N__32085\,
            in2 => \N__28510\,
            in3 => \N__31927\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34378\,
            ce => \N__31621\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__28509\,
            in2 => \N__31972\,
            in3 => \N__31745\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIL79C1_15_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31548\,
            in1 => \_gnd_net_\,
            in2 => \N__28495\,
            in3 => \N__28492\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__31902\,
            in2 => \N__31797\,
            in3 => \N__28443\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34378\,
            ce => \N__31621\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32248\,
            in2 => \N__32236\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28480\,
            in2 => \_gnd_net_\,
            in3 => \N__28462\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28459\,
            in2 => \_gnd_net_\,
            in3 => \N__28429\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30891\,
            in2 => \_gnd_net_\,
            in3 => \N__28426\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31296\,
            in2 => \_gnd_net_\,
            in3 => \N__28423\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30898\,
            in2 => \_gnd_net_\,
            in3 => \N__28420\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28666\,
            in2 => \_gnd_net_\,
            in3 => \N__28624\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28617\,
            in2 => \_gnd_net_\,
            in3 => \N__28582\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28716\,
            in2 => \_gnd_net_\,
            in3 => \N__28561\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28689\,
            in2 => \_gnd_net_\,
            in3 => \N__28528\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31480\,
            in2 => \_gnd_net_\,
            in3 => \N__28525\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31428\,
            in2 => \_gnd_net_\,
            in3 => \N__28522\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31453\,
            in2 => \_gnd_net_\,
            in3 => \N__28519\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31410\,
            in2 => \_gnd_net_\,
            in3 => \N__28516\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28513\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32164\,
            in1 => \N__31952\,
            in2 => \N__31365\,
            in3 => \N__31766\,
            lcout => \VPP_VDDQ.count_2_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31949\,
            in1 => \N__28656\,
            in2 => \N__32181\,
            in3 => \N__31784\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => \VPP_VDDQ.count_2_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_0_7_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__31606\,
            in1 => \N__28645\,
            in2 => \N__28720\,
            in3 => \N__28717\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_1_7_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__31393\,
            in1 => \N__31479\,
            in2 => \N__28693\,
            in3 => \N__28690\,
            lcout => \VPP_VDDQ.un9_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_7_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31605\,
            in1 => \N__28644\,
            in2 => \_gnd_net_\,
            in3 => \N__28672\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31950\,
            in1 => \N__28657\,
            in2 => \N__32182\,
            in3 => \N__31786\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34434\,
            ce => \N__31632\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__31783\,
            in1 => \N__32173\,
            in2 => \N__32235\,
            in3 => \N__31948\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIT1QU_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31604\,
            in2 => \N__28636\,
            in3 => \N__28630\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__31785\,
            in1 => \N__32177\,
            in2 => \N__28633\,
            in3 => \N__31951\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34434\,
            ce => \N__31632\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJ0RD_3_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28741\,
            in1 => \N__33289\,
            in2 => \N__33488\,
            in3 => \N__32349\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33475\,
            in2 => \_gnd_net_\,
            in3 => \N__32350\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33999\,
            ce => \N__33324\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33483\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33999\,
            ce => \N__33324\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINA66_14_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__28726\,
            in2 => \N__33490\,
            in3 => \N__32433\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => \POWERLED.count_clkZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_13_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28735\,
            in3 => \N__32469\,
            lcout => \POWERLED.count_clk_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIL756_13_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__28732\,
            in2 => \N__33489\,
            in3 => \N__32454\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33484\,
            lcout => \POWERLED.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33999\,
            ce => \N__33324\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33476\,
            in2 => \_gnd_net_\,
            in3 => \N__32335\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33999\,
            ce => \N__33324\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33411\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIQF8B_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28762\,
            in2 => \N__28786\,
            in3 => \N__33285\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => \POWERLED.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33019\,
            in2 => \N__28783\,
            in3 => \N__33412\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIRG8B_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32587\,
            in2 => \N__28780\,
            in3 => \N__33286\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIP9UD_6_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__33288\,
            in1 => \N__33416\,
            in2 => \N__28771\,
            in3 => \N__32316\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIL3SD_4_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28777\,
            in1 => \N__33287\,
            in2 => \N__33458\,
            in3 => \N__32334\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32317\,
            in2 => \_gnd_net_\,
            in3 => \N__33418\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34438\,
            ce => \N__33317\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__33417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32612\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34438\,
            ce => \N__33317\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__32823\,
            in1 => \N__32735\,
            in2 => \N__33024\,
            in3 => \N__32414\,
            lcout => \POWERLED.count_clk_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__32413\,
            in1 => \N__33014\,
            in2 => \N__32737\,
            in3 => \N__32822\,
            lcout => \POWERLED.count_clk_RNIZ0Z_1\,
            ltout => \POWERLED.count_clk_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__29322\,
            in1 => \_gnd_net_\,
            in2 => \N__29119\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_1_1_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__31114\,
            in1 => \N__29109\,
            in2 => \N__29095\,
            in3 => \N__28910\,
            lcout => \POWERLED.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__32540\,
            in1 => \N__33539\,
            in2 => \N__32418\,
            in3 => \N__32514\,
            lcout => \POWERLED.un2_count_clk_15_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI18EF2_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101011"
        )
    port map (
            in0 => \N__29092\,
            in1 => \N__30228\,
            in2 => \N__31153\,
            in3 => \N__29621\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIH9594_1_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__29155\,
            in1 => \N__29077\,
            in2 => \N__29071\,
            in3 => \N__32484\,
            lcout => \POWERLED.func_state_RNIH9594_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOTGO_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__29591\,
            in1 => \N__29050\,
            in2 => \N__29334\,
            in3 => \N__31110\,
            lcout => \POWERLED.N_291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29049\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29488\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_4_i_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRKB61_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011111111"
        )
    port map (
            in0 => \N__29518\,
            in1 => \N__28955\,
            in2 => \N__28831\,
            in3 => \N__31109\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIUHKR2_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__28828\,
            in1 => \N__28795\,
            in2 => \N__28789\,
            in3 => \N__29620\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1U3S4_1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__30055\,
            in1 => \N__30002\,
            in2 => \N__29833\,
            in3 => \N__29713\,
            lcout => \POWERLED.count_clk_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29329\,
            in3 => \N__29590\,
            lcout => \POWERLED.func_state_RNI_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__29592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29294\,
            lcout => \POWERLED.N_176\,
            ltout => \POWERLED.N_176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29512\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2218_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__29480\,
            in1 => \N__29344\,
            in2 => \N__29335\,
            in3 => \N__32882\,
            lcout => \POWERLED.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30218\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__30371\,
            in1 => \N__30097\,
            in2 => \N__30229\,
            in3 => \N__30288\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_64_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__29127\,
            in1 => \N__30303\,
            in2 => \N__29134\,
            in3 => \N__34855\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__34856\,
            in1 => \_gnd_net_\,
            in2 => \N__29131\,
            in3 => \N__30319\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__30273\,
            in1 => \N__30370\,
            in2 => \_gnd_net_\,
            in3 => \N__30214\,
            lcout => \VPP_VDDQ.curr_state_7_0\,
            ltout => \VPP_VDDQ.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI2OB42_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30096\,
            in2 => \N__30313\,
            in3 => \N__30274\,
            lcout => \VPP_VDDQ.N_66_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__30359\,
            in1 => \N__30095\,
            in2 => \N__30237\,
            in3 => \N__30276\,
            lcout => \N_246\,
            ltout => \N_246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_43_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__30289\,
            in1 => \N__30072\,
            in2 => \N__30292\,
            in3 => \N__34843\,
            lcout => \G_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNID2IU_0_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30094\,
            in2 => \_gnd_net_\,
            in3 => \N__30275\,
            lcout => \N_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__30358\,
            in1 => \N__30277\,
            in2 => \_gnd_net_\,
            in3 => \N__30233\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34431\,
            ce => \N__34714\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33081\,
            in1 => \N__33096\,
            in2 => \N__33115\,
            in3 => \N__33657\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30649\,
            in1 => \N__30643\,
            in2 => \N__30079\,
            in3 => \N__30061\,
            lcout => \VPP_VDDQ_un6_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33672\,
            in1 => \N__33144\,
            in2 => \N__33613\,
            in3 => \N__33129\,
            lcout => \VPP_VDDQ.un6_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33627\,
            in1 => \N__33642\,
            in2 => \N__33160\,
            in3 => \N__33594\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34587\,
            in1 => \N__34473\,
            in2 => \N__33565\,
            in3 => \N__33579\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34857\,
            in2 => \_gnd_net_\,
            in3 => \N__33703\,
            lcout => \VPP_VDDQ.N_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32107\,
            lcout => \VPP_VDDQ.N_2192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30726\,
            lcout => \VPP_VDDQ.N_361_0\,
            ltout => \VPP_VDDQ.N_361_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__30548\,
            in1 => \_gnd_net_\,
            in2 => \N__30433\,
            in3 => \N__31925\,
            lcout => \VPP_VDDQ.N_62\,
            ltout => \VPP_VDDQ.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__30400\,
            in1 => \N__31971\,
            in2 => \N__30430\,
            in3 => \N__30808\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => \VPP_VDDQ.delayed_vddq_ok_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__30328\,
            in1 => \N__30718\,
            in2 => \N__30427\,
            in3 => \N__30402\,
            lcout => \VPP_VDDQ_delayed_vddq_ok\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__30401\,
            in1 => \N__30327\,
            in2 => \N__30337\,
            in3 => \N__30717\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34222\,
            ce => 'H',
            sr => \N__30703\
        );

    \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__30817\,
            in1 => \N__30803\,
            in2 => \N__30730\,
            in3 => \N__31926\,
            lcout => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30716\,
            lcout => \VPP_VDDQ.N_62_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__32090\,
            in1 => \N__31912\,
            in2 => \N__31796\,
            in3 => \N__31342\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJ48C1_14_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31324\,
            in2 => \N__30694\,
            in3 => \N__31552\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32088\,
            in1 => \N__31910\,
            in2 => \N__30687\,
            in3 => \N__31746\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIHA461_4_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30667\,
            in2 => \N__30691\,
            in3 => \N__31550\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32091\,
            in1 => \N__31913\,
            in2 => \N__30688\,
            in3 => \N__31748\,
            lcout => \VPP_VDDQ.count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34412\,
            ce => \N__31633\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31914\,
            in1 => \N__30660\,
            in2 => \N__32150\,
            in3 => \N__31770\,
            lcout => \VPP_VDDQ.count_2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34412\,
            ce => \N__31633\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32089\,
            in1 => \N__31911\,
            in2 => \N__30661\,
            in3 => \N__31747\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJD561_5_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31306\,
            in1 => \_gnd_net_\,
            in2 => \N__31300\,
            in3 => \N__31551\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__31285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31140\,
            lcout => \PCH_PWRGD.N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__31210\,
            in2 => \N__31198\,
            in3 => \N__31189\,
            lcout => OPEN,
            ltout => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__31141\,
            in1 => \_gnd_net_\,
            in2 => \N__30961\,
            in3 => \N__30958\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI38QU_6_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30879\,
            in1 => \N__30825\,
            in2 => \_gnd_net_\,
            in3 => \N__31589\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI38QU_0_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__31590\,
            in1 => \N__30892\,
            in2 => \N__30829\,
            in3 => \N__30880\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIOUR33_1_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31315\,
            in1 => \N__30868\,
            in2 => \N__30862\,
            in3 => \N__30859\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => \VPP_VDDQ.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__30846\,
            in1 => \N__32165\,
            in2 => \N__30832\,
            in3 => \N__31943\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34350\,
            ce => \N__31594\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFU5C1_12_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31372\,
            in1 => \N__31618\,
            in2 => \_gnd_net_\,
            in3 => \N__31465\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32146\,
            in1 => \N__31941\,
            in2 => \N__31386\,
            in3 => \N__31762\,
            lcout => \VPP_VDDQ.count_2_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIH17C1_13_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31348\,
            in1 => \N__31459\,
            in2 => \_gnd_net_\,
            in3 => \N__31619\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => \VPP_VDDQ.count_2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31447\,
            in1 => \N__31429\,
            in2 => \N__31417\,
            in3 => \N__31414\,
            lcout => \VPP_VDDQ.un9_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32147\,
            in1 => \N__31942\,
            in2 => \N__31387\,
            in3 => \N__31764\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34433\,
            ce => \N__31622\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31763\,
            in1 => \N__32149\,
            in2 => \N__31366\,
            in3 => \N__31947\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34433\,
            ce => \N__31622\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32148\,
            in1 => \N__31338\,
            in2 => \N__31979\,
            in3 => \N__31765\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34433\,
            ce => \N__31622\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32151\,
            in1 => \N__31973\,
            in2 => \N__32206\,
            in3 => \N__31779\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000011"
        )
    port map (
            in0 => \N__32257\,
            in1 => \N__32227\,
            in2 => \N__32194\,
            in3 => \N__31568\,
            lcout => \VPP_VDDQ.un9_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31567\,
            in1 => \N__32190\,
            in2 => \_gnd_net_\,
            in3 => \N__32256\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => \VPP_VDDQ.un1_count_2_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32239\,
            in3 => \N__32228\,
            lcout => \VPP_VDDQ.count_2_RNIZ0Z_1\,
            ltout => \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32152\,
            in1 => \N__31974\,
            in2 => \N__32197\,
            in3 => \N__31781\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34348\,
            ce => \N__31569\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31780\,
            in1 => \N__32153\,
            in2 => \N__32002\,
            in3 => \N__31975\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34348\,
            ce => \N__31569\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32154\,
            in1 => \N__32001\,
            in2 => \N__31989\,
            in3 => \N__31782\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31642\,
            in2 => \N__31636\,
            in3 => \N__31566\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32610\,
            in2 => \N__33020\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32635\,
            in3 => \N__31468\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33060\,
            in3 => \N__32338\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33543\,
            in3 => \N__32323\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__33485\,
            in1 => \_gnd_net_\,
            in2 => \N__32419\,
            in3 => \N__32320\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32544\,
            in3 => \N__32308\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__33486\,
            in1 => \_gnd_net_\,
            in2 => \N__32728\,
            in3 => \N__32290\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__33487\,
            in1 => \N__32842\,
            in2 => \_gnd_net_\,
            in3 => \N__32287\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__33453\,
            in1 => \_gnd_net_\,
            in2 => \N__32824\,
            in3 => \N__32266\,
            lcout => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33043\,
            in3 => \N__32263\,
            lcout => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9\,
            carryout => \POWERLED.un1_count_clk_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32683\,
            in3 => \N__32260\,
            lcout => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10\,
            carryout => \POWERLED.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__33455\,
            in1 => \_gnd_net_\,
            in2 => \N__32752\,
            in3 => \N__32473\,
            lcout => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11\,
            carryout => \POWERLED.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32470\,
            in3 => \N__32446\,
            lcout => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12\,
            carryout => \POWERLED.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32443\,
            in3 => \N__32425\,
            lcout => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__32356\,
            in1 => \N__33456\,
            in2 => \_gnd_net_\,
            in3 => \N__32422\,
            lcout => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32766\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34430\,
            ce => \N__33331\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIN6TD_5_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32377\,
            in2 => \N__33292\,
            in3 => \N__32388\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32389\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__33333\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__33333\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPD76_15_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33267\,
            in1 => \N__32371\,
            in2 => \_gnd_net_\,
            in3 => \N__32364\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => \POWERLED.count_clkZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_15_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32617\,
            in3 => \N__32611\,
            lcout => \POWERLED.count_clk_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__33471\,
            in1 => \N__32614\,
            in2 => \_gnd_net_\,
            in3 => \N__33018\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__33333\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNITF0E_8_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33257\,
            in1 => \N__32569\,
            in2 => \_gnd_net_\,
            in3 => \N__32580\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__33333\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32557\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33457\,
            lcout => \POWERLED.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34421\,
            ce => \N__33316\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8SH6_10_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__32563\,
            in1 => \N__33454\,
            in2 => \N__33320\,
            in3 => \N__32556\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => \POWERLED.count_clkZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33067\,
            in1 => \N__32545\,
            in2 => \N__32521\,
            in3 => \N__32679\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_8_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__32841\,
            in1 => \N__32518\,
            in2 => \N__32500\,
            in3 => \N__33496\,
            lcout => \POWERLED.N_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_10_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33066\,
            in1 => \N__33039\,
            in2 => \N__33025\,
            in3 => \N__33507\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_15_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_10_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32782\,
            in2 => \N__32980\,
            in3 => \N__32977\,
            lcout => \POWERLED.un2_count_clk_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_8_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__32840\,
            in1 => \_gnd_net_\,
            in2 => \N__32692\,
            in3 => \N__32821\,
            lcout => \POWERLED.un2_count_clk_15_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJ446_12_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33237\,
            in1 => \N__32776\,
            in2 => \_gnd_net_\,
            in3 => \N__32767\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => \POWERLED.count_clkZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_12_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32740\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_RNIZ0Z_12\,
            ltout => \POWERLED.count_clk_RNIZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_11_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32631\,
            in1 => \N__32736\,
            in2 => \N__32695\,
            in3 => \N__32678\,
            lcout => \POWERLED.un2_count_clk_15_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIH136_11_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__33469\,
            in1 => \N__33236\,
            in2 => \N__33343\,
            in3 => \N__33354\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32658\,
            in2 => \_gnd_net_\,
            in3 => \N__33470\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34450\,
            ce => \N__33334\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIHTPD_2_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__32659\,
            in1 => \N__33459\,
            in2 => \N__32644\,
            in3 => \N__33235\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => \POWERLED.count_clkZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_2_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33547\,
            in1 => \N__33520\,
            in2 => \N__33514\,
            in3 => \N__33511\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33460\,
            in2 => \_gnd_net_\,
            in3 => \N__33355\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34450\,
            ce => \N__33334\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34880\,
            in1 => \N__33159\,
            in2 => \N__33175\,
            in3 => \N__33174\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34870\,
            in1 => \N__33145\,
            in2 => \_gnd_net_\,
            in3 => \N__33133\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34881\,
            in1 => \N__33130\,
            in2 => \_gnd_net_\,
            in3 => \N__33118\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34871\,
            in1 => \N__33114\,
            in2 => \_gnd_net_\,
            in3 => \N__33100\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_4_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34882\,
            in1 => \N__33097\,
            in2 => \_gnd_net_\,
            in3 => \N__33085\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34872\,
            in1 => \N__33082\,
            in2 => \_gnd_net_\,
            in3 => \N__33070\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_6_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34883\,
            in1 => \N__33673\,
            in2 => \_gnd_net_\,
            in3 => \N__33661\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_7_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34873\,
            in1 => \N__33658\,
            in2 => \_gnd_net_\,
            in3 => \N__33646\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__34462\,
            ce => 'H',
            sr => \N__33704\
        );

    \VPP_VDDQ.count_8_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34887\,
            in1 => \N__33643\,
            in2 => \_gnd_net_\,
            in3 => \N__33631\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.count_9_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34876\,
            in1 => \N__33628\,
            in2 => \_gnd_net_\,
            in3 => \N__33616\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.count_10_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34884\,
            in1 => \N__33612\,
            in2 => \_gnd_net_\,
            in3 => \N__33598\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.count_11_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34874\,
            in1 => \N__33595\,
            in2 => \_gnd_net_\,
            in3 => \N__33583\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.count_12_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34885\,
            in1 => \N__33580\,
            in2 => \_gnd_net_\,
            in3 => \N__33568\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.count_13_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34875\,
            in1 => \N__33564\,
            in2 => \_gnd_net_\,
            in3 => \N__33550\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.count_14_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34886\,
            in1 => \N__34588\,
            in2 => \_gnd_net_\,
            in3 => \N__34576\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__33709\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34573\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34474\,
            in2 => \_gnd_net_\,
            in3 => \N__34477\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34461\,
            ce => \N__33715\,
            sr => \N__33705\
        );
end \INTERFACE\;
