// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 14 2022 10:43:49

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    input SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    input VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    input VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__39838;
    wire N__39837;
    wire N__39836;
    wire N__39829;
    wire N__39828;
    wire N__39827;
    wire N__39820;
    wire N__39819;
    wire N__39818;
    wire N__39811;
    wire N__39810;
    wire N__39809;
    wire N__39802;
    wire N__39801;
    wire N__39800;
    wire N__39793;
    wire N__39792;
    wire N__39791;
    wire N__39784;
    wire N__39783;
    wire N__39782;
    wire N__39775;
    wire N__39774;
    wire N__39773;
    wire N__39766;
    wire N__39765;
    wire N__39764;
    wire N__39757;
    wire N__39756;
    wire N__39755;
    wire N__39748;
    wire N__39747;
    wire N__39746;
    wire N__39739;
    wire N__39738;
    wire N__39737;
    wire N__39730;
    wire N__39729;
    wire N__39728;
    wire N__39721;
    wire N__39720;
    wire N__39719;
    wire N__39712;
    wire N__39711;
    wire N__39710;
    wire N__39703;
    wire N__39702;
    wire N__39701;
    wire N__39694;
    wire N__39693;
    wire N__39692;
    wire N__39685;
    wire N__39684;
    wire N__39683;
    wire N__39676;
    wire N__39675;
    wire N__39674;
    wire N__39667;
    wire N__39666;
    wire N__39665;
    wire N__39658;
    wire N__39657;
    wire N__39656;
    wire N__39649;
    wire N__39648;
    wire N__39647;
    wire N__39640;
    wire N__39639;
    wire N__39638;
    wire N__39631;
    wire N__39630;
    wire N__39629;
    wire N__39622;
    wire N__39621;
    wire N__39620;
    wire N__39613;
    wire N__39612;
    wire N__39611;
    wire N__39604;
    wire N__39603;
    wire N__39602;
    wire N__39595;
    wire N__39594;
    wire N__39593;
    wire N__39586;
    wire N__39585;
    wire N__39584;
    wire N__39577;
    wire N__39576;
    wire N__39575;
    wire N__39568;
    wire N__39567;
    wire N__39566;
    wire N__39559;
    wire N__39558;
    wire N__39557;
    wire N__39550;
    wire N__39549;
    wire N__39548;
    wire N__39541;
    wire N__39540;
    wire N__39539;
    wire N__39532;
    wire N__39531;
    wire N__39530;
    wire N__39523;
    wire N__39522;
    wire N__39521;
    wire N__39514;
    wire N__39513;
    wire N__39512;
    wire N__39505;
    wire N__39504;
    wire N__39503;
    wire N__39496;
    wire N__39495;
    wire N__39494;
    wire N__39487;
    wire N__39486;
    wire N__39485;
    wire N__39478;
    wire N__39477;
    wire N__39476;
    wire N__39469;
    wire N__39468;
    wire N__39467;
    wire N__39460;
    wire N__39459;
    wire N__39458;
    wire N__39451;
    wire N__39450;
    wire N__39449;
    wire N__39442;
    wire N__39441;
    wire N__39440;
    wire N__39433;
    wire N__39432;
    wire N__39431;
    wire N__39424;
    wire N__39423;
    wire N__39422;
    wire N__39415;
    wire N__39414;
    wire N__39413;
    wire N__39406;
    wire N__39405;
    wire N__39404;
    wire N__39397;
    wire N__39396;
    wire N__39395;
    wire N__39388;
    wire N__39387;
    wire N__39386;
    wire N__39379;
    wire N__39378;
    wire N__39377;
    wire N__39370;
    wire N__39369;
    wire N__39368;
    wire N__39361;
    wire N__39360;
    wire N__39359;
    wire N__39352;
    wire N__39351;
    wire N__39350;
    wire N__39343;
    wire N__39342;
    wire N__39341;
    wire N__39334;
    wire N__39333;
    wire N__39332;
    wire N__39325;
    wire N__39324;
    wire N__39323;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39297;
    wire N__39296;
    wire N__39295;
    wire N__39294;
    wire N__39289;
    wire N__39288;
    wire N__39287;
    wire N__39286;
    wire N__39285;
    wire N__39284;
    wire N__39283;
    wire N__39282;
    wire N__39281;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39273;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39256;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39224;
    wire N__39219;
    wire N__39214;
    wire N__39209;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39195;
    wire N__39186;
    wire N__39185;
    wire N__39184;
    wire N__39183;
    wire N__39182;
    wire N__39181;
    wire N__39180;
    wire N__39179;
    wire N__39178;
    wire N__39177;
    wire N__39176;
    wire N__39175;
    wire N__39172;
    wire N__39171;
    wire N__39170;
    wire N__39169;
    wire N__39168;
    wire N__39167;
    wire N__39166;
    wire N__39165;
    wire N__39162;
    wire N__39161;
    wire N__39160;
    wire N__39159;
    wire N__39158;
    wire N__39155;
    wire N__39154;
    wire N__39147;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39132;
    wire N__39129;
    wire N__39128;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39117;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39095;
    wire N__39094;
    wire N__39093;
    wire N__39092;
    wire N__39091;
    wire N__39088;
    wire N__39087;
    wire N__39086;
    wire N__39085;
    wire N__39084;
    wire N__39077;
    wire N__39074;
    wire N__39061;
    wire N__39060;
    wire N__39059;
    wire N__39058;
    wire N__39057;
    wire N__39056;
    wire N__39055;
    wire N__39054;
    wire N__39053;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39012;
    wire N__39007;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38987;
    wire N__38984;
    wire N__38983;
    wire N__38982;
    wire N__38981;
    wire N__38980;
    wire N__38971;
    wire N__38968;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38945;
    wire N__38942;
    wire N__38935;
    wire N__38930;
    wire N__38925;
    wire N__38918;
    wire N__38913;
    wire N__38910;
    wire N__38905;
    wire N__38900;
    wire N__38897;
    wire N__38888;
    wire N__38877;
    wire N__38862;
    wire N__38859;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38851;
    wire N__38850;
    wire N__38849;
    wire N__38848;
    wire N__38847;
    wire N__38846;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38832;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38815;
    wire N__38814;
    wire N__38813;
    wire N__38812;
    wire N__38809;
    wire N__38804;
    wire N__38803;
    wire N__38802;
    wire N__38801;
    wire N__38798;
    wire N__38791;
    wire N__38788;
    wire N__38781;
    wire N__38778;
    wire N__38773;
    wire N__38766;
    wire N__38761;
    wire N__38758;
    wire N__38749;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38725;
    wire N__38724;
    wire N__38723;
    wire N__38722;
    wire N__38719;
    wire N__38718;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38704;
    wire N__38697;
    wire N__38694;
    wire N__38693;
    wire N__38688;
    wire N__38685;
    wire N__38680;
    wire N__38679;
    wire N__38678;
    wire N__38677;
    wire N__38676;
    wire N__38675;
    wire N__38674;
    wire N__38671;
    wire N__38666;
    wire N__38659;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38645;
    wire N__38642;
    wire N__38641;
    wire N__38632;
    wire N__38627;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38615;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38595;
    wire N__38592;
    wire N__38591;
    wire N__38590;
    wire N__38589;
    wire N__38588;
    wire N__38587;
    wire N__38584;
    wire N__38579;
    wire N__38572;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38562;
    wire N__38561;
    wire N__38560;
    wire N__38557;
    wire N__38556;
    wire N__38555;
    wire N__38554;
    wire N__38553;
    wire N__38552;
    wire N__38547;
    wire N__38544;
    wire N__38539;
    wire N__38530;
    wire N__38529;
    wire N__38528;
    wire N__38527;
    wire N__38526;
    wire N__38525;
    wire N__38524;
    wire N__38523;
    wire N__38518;
    wire N__38517;
    wire N__38516;
    wire N__38515;
    wire N__38510;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38488;
    wire N__38485;
    wire N__38484;
    wire N__38477;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38447;
    wire N__38444;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38418;
    wire N__38417;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38409;
    wire N__38408;
    wire N__38405;
    wire N__38404;
    wire N__38399;
    wire N__38392;
    wire N__38391;
    wire N__38388;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38352;
    wire N__38351;
    wire N__38348;
    wire N__38347;
    wire N__38346;
    wire N__38345;
    wire N__38344;
    wire N__38343;
    wire N__38342;
    wire N__38341;
    wire N__38340;
    wire N__38339;
    wire N__38338;
    wire N__38337;
    wire N__38336;
    wire N__38333;
    wire N__38332;
    wire N__38331;
    wire N__38330;
    wire N__38329;
    wire N__38328;
    wire N__38321;
    wire N__38316;
    wire N__38313;
    wire N__38312;
    wire N__38311;
    wire N__38310;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38296;
    wire N__38295;
    wire N__38292;
    wire N__38287;
    wire N__38280;
    wire N__38275;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38259;
    wire N__38258;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38237;
    wire N__38232;
    wire N__38229;
    wire N__38228;
    wire N__38227;
    wire N__38220;
    wire N__38215;
    wire N__38204;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38183;
    wire N__38180;
    wire N__38169;
    wire N__38168;
    wire N__38167;
    wire N__38166;
    wire N__38163;
    wire N__38162;
    wire N__38161;
    wire N__38160;
    wire N__38159;
    wire N__38158;
    wire N__38155;
    wire N__38154;
    wire N__38145;
    wire N__38140;
    wire N__38137;
    wire N__38136;
    wire N__38135;
    wire N__38132;
    wire N__38131;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38108;
    wire N__38107;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38081;
    wire N__38076;
    wire N__38071;
    wire N__38064;
    wire N__38061;
    wire N__38054;
    wire N__38037;
    wire N__38036;
    wire N__38035;
    wire N__38034;
    wire N__38033;
    wire N__38032;
    wire N__38031;
    wire N__38030;
    wire N__38029;
    wire N__38028;
    wire N__38027;
    wire N__38024;
    wire N__38023;
    wire N__38022;
    wire N__38019;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38003;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37981;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37958;
    wire N__37953;
    wire N__37942;
    wire N__37935;
    wire N__37934;
    wire N__37931;
    wire N__37930;
    wire N__37929;
    wire N__37928;
    wire N__37927;
    wire N__37924;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37916;
    wire N__37915;
    wire N__37912;
    wire N__37911;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37881;
    wire N__37878;
    wire N__37877;
    wire N__37876;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37872;
    wire N__37871;
    wire N__37870;
    wire N__37865;
    wire N__37862;
    wire N__37855;
    wire N__37850;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37832;
    wire N__37825;
    wire N__37820;
    wire N__37817;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37769;
    wire N__37768;
    wire N__37767;
    wire N__37766;
    wire N__37765;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37761;
    wire N__37758;
    wire N__37757;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37749;
    wire N__37748;
    wire N__37747;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37731;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37706;
    wire N__37705;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37682;
    wire N__37677;
    wire N__37670;
    wire N__37665;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37595;
    wire N__37594;
    wire N__37593;
    wire N__37590;
    wire N__37589;
    wire N__37588;
    wire N__37585;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37565;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37549;
    wire N__37544;
    wire N__37541;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37527;
    wire N__37524;
    wire N__37519;
    wire N__37512;
    wire N__37511;
    wire N__37510;
    wire N__37509;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37503;
    wire N__37502;
    wire N__37501;
    wire N__37500;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37454;
    wire N__37449;
    wire N__37446;
    wire N__37441;
    wire N__37434;
    wire N__37433;
    wire N__37432;
    wire N__37431;
    wire N__37430;
    wire N__37429;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37417;
    wire N__37412;
    wire N__37409;
    wire N__37408;
    wire N__37403;
    wire N__37402;
    wire N__37399;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37380;
    wire N__37375;
    wire N__37372;
    wire N__37365;
    wire N__37362;
    wire N__37361;
    wire N__37358;
    wire N__37357;
    wire N__37356;
    wire N__37351;
    wire N__37350;
    wire N__37347;
    wire N__37346;
    wire N__37345;
    wire N__37344;
    wire N__37343;
    wire N__37342;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37327;
    wire N__37324;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37316;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37293;
    wire N__37292;
    wire N__37291;
    wire N__37290;
    wire N__37289;
    wire N__37284;
    wire N__37283;
    wire N__37282;
    wire N__37279;
    wire N__37278;
    wire N__37277;
    wire N__37272;
    wire N__37265;
    wire N__37262;
    wire N__37257;
    wire N__37254;
    wire N__37249;
    wire N__37246;
    wire N__37241;
    wire N__37234;
    wire N__37229;
    wire N__37224;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37190;
    wire N__37187;
    wire N__37182;
    wire N__37179;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37154;
    wire N__37149;
    wire N__37148;
    wire N__37145;
    wire N__37144;
    wire N__37143;
    wire N__37142;
    wire N__37141;
    wire N__37140;
    wire N__37139;
    wire N__37136;
    wire N__37135;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37127;
    wire N__37126;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37109;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37101;
    wire N__37100;
    wire N__37099;
    wire N__37096;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37088;
    wire N__37087;
    wire N__37086;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37072;
    wire N__37071;
    wire N__37070;
    wire N__37069;
    wire N__37068;
    wire N__37067;
    wire N__37064;
    wire N__37063;
    wire N__37062;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37027;
    wire N__37022;
    wire N__37019;
    wire N__37018;
    wire N__37015;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37007;
    wire N__37006;
    wire N__37003;
    wire N__37002;
    wire N__37001;
    wire N__36998;
    wire N__36997;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36973;
    wire N__36970;
    wire N__36969;
    wire N__36968;
    wire N__36967;
    wire N__36966;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36955;
    wire N__36948;
    wire N__36943;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36891;
    wire N__36890;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36863;
    wire N__36862;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36840;
    wire N__36837;
    wire N__36836;
    wire N__36835;
    wire N__36834;
    wire N__36831;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36823;
    wire N__36822;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36810;
    wire N__36805;
    wire N__36802;
    wire N__36801;
    wire N__36800;
    wire N__36793;
    wire N__36788;
    wire N__36781;
    wire N__36776;
    wire N__36775;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36745;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36733;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36709;
    wire N__36704;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36673;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36655;
    wire N__36652;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36640;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36612;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36573;
    wire N__36570;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36544;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36528;
    wire N__36523;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36498;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36482;
    wire N__36473;
    wire N__36470;
    wire N__36463;
    wire N__36454;
    wire N__36447;
    wire N__36438;
    wire N__36437;
    wire N__36436;
    wire N__36433;
    wire N__36428;
    wire N__36427;
    wire N__36424;
    wire N__36421;
    wire N__36414;
    wire N__36407;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36391;
    wire N__36388;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36366;
    wire N__36363;
    wire N__36362;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36341;
    wire N__36338;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36310;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36274;
    wire N__36271;
    wire N__36266;
    wire N__36263;
    wire N__36256;
    wire N__36253;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36223;
    wire N__36222;
    wire N__36221;
    wire N__36220;
    wire N__36217;
    wire N__36216;
    wire N__36215;
    wire N__36212;
    wire N__36211;
    wire N__36210;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36205;
    wire N__36204;
    wire N__36203;
    wire N__36200;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36175;
    wire N__36174;
    wire N__36173;
    wire N__36170;
    wire N__36163;
    wire N__36158;
    wire N__36151;
    wire N__36140;
    wire N__36129;
    wire N__36126;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36096;
    wire N__36091;
    wire N__36088;
    wire N__36085;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36061;
    wire N__36060;
    wire N__36059;
    wire N__36058;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36042;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36032;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__36006;
    wire N__36005;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35985;
    wire N__35980;
    wire N__35975;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35948;
    wire N__35947;
    wire N__35946;
    wire N__35941;
    wire N__35932;
    wire N__35921;
    wire N__35920;
    wire N__35919;
    wire N__35914;
    wire N__35907;
    wire N__35902;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35888;
    wire N__35883;
    wire N__35880;
    wire N__35879;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35864;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35856;
    wire N__35853;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35845;
    wire N__35838;
    wire N__35837;
    wire N__35836;
    wire N__35835;
    wire N__35834;
    wire N__35833;
    wire N__35832;
    wire N__35831;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35817;
    wire N__35812;
    wire N__35809;
    wire N__35808;
    wire N__35805;
    wire N__35800;
    wire N__35799;
    wire N__35798;
    wire N__35793;
    wire N__35792;
    wire N__35791;
    wire N__35790;
    wire N__35789;
    wire N__35788;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35776;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35670;
    wire N__35661;
    wire N__35658;
    wire N__35653;
    wire N__35646;
    wire N__35643;
    wire N__35638;
    wire N__35633;
    wire N__35628;
    wire N__35621;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35579;
    wire N__35574;
    wire N__35571;
    wire N__35570;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35555;
    wire N__35554;
    wire N__35549;
    wire N__35546;
    wire N__35545;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35537;
    wire N__35536;
    wire N__35531;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35502;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35486;
    wire N__35481;
    wire N__35478;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35468;
    wire N__35467;
    wire N__35466;
    wire N__35465;
    wire N__35464;
    wire N__35463;
    wire N__35462;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35450;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35435;
    wire N__35434;
    wire N__35429;
    wire N__35424;
    wire N__35423;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35388;
    wire N__35385;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35223;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35210;
    wire N__35209;
    wire N__35206;
    wire N__35205;
    wire N__35204;
    wire N__35203;
    wire N__35200;
    wire N__35199;
    wire N__35196;
    wire N__35195;
    wire N__35194;
    wire N__35193;
    wire N__35190;
    wire N__35189;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35177;
    wire N__35170;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35138;
    wire N__35135;
    wire N__35120;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35108;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35088;
    wire N__35085;
    wire N__35084;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35070;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35038;
    wire N__35031;
    wire N__35028;
    wire N__35027;
    wire N__35026;
    wire N__35025;
    wire N__35020;
    wire N__35017;
    wire N__35016;
    wire N__35015;
    wire N__35012;
    wire N__35011;
    wire N__35010;
    wire N__35009;
    wire N__35008;
    wire N__35007;
    wire N__35006;
    wire N__35003;
    wire N__35002;
    wire N__34997;
    wire N__34994;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34982;
    wire N__34979;
    wire N__34978;
    wire N__34977;
    wire N__34976;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34955;
    wire N__34954;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34936;
    wire N__34933;
    wire N__34926;
    wire N__34923;
    wire N__34918;
    wire N__34915;
    wire N__34910;
    wire N__34901;
    wire N__34878;
    wire N__34875;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34838;
    wire N__34837;
    wire N__34834;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34823;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34801;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34786;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34771;
    wire N__34770;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34748;
    wire N__34741;
    wire N__34738;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34673;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34631;
    wire N__34626;
    wire N__34623;
    wire N__34622;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34607;
    wire N__34606;
    wire N__34605;
    wire N__34604;
    wire N__34601;
    wire N__34600;
    wire N__34599;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34580;
    wire N__34575;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34552;
    wire N__34549;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34528;
    wire N__34521;
    wire N__34512;
    wire N__34509;
    wire N__34508;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34455;
    wire N__34452;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34412;
    wire N__34411;
    wire N__34408;
    wire N__34403;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34388;
    wire N__34387;
    wire N__34384;
    wire N__34383;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34379;
    wire N__34378;
    wire N__34373;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34363;
    wire N__34362;
    wire N__34357;
    wire N__34356;
    wire N__34355;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34343;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34324;
    wire N__34323;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34285;
    wire N__34278;
    wire N__34275;
    wire N__34266;
    wire N__34265;
    wire N__34262;
    wire N__34261;
    wire N__34260;
    wire N__34259;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34251;
    wire N__34242;
    wire N__34241;
    wire N__34240;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34224;
    wire N__34221;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34193;
    wire N__34190;
    wire N__34189;
    wire N__34188;
    wire N__34187;
    wire N__34184;
    wire N__34183;
    wire N__34178;
    wire N__34175;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34165;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34136;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34097;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34051;
    wire N__34050;
    wire N__34049;
    wire N__34048;
    wire N__34047;
    wire N__34042;
    wire N__34037;
    wire N__34036;
    wire N__34033;
    wire N__34032;
    wire N__34031;
    wire N__34030;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34008;
    wire N__34005;
    wire N__34000;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33984;
    wire N__33981;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33942;
    wire N__33941;
    wire N__33940;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33894;
    wire N__33893;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33836;
    wire N__33835;
    wire N__33832;
    wire N__33831;
    wire N__33830;
    wire N__33827;
    wire N__33826;
    wire N__33825;
    wire N__33824;
    wire N__33823;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33812;
    wire N__33811;
    wire N__33810;
    wire N__33809;
    wire N__33808;
    wire N__33807;
    wire N__33804;
    wire N__33803;
    wire N__33802;
    wire N__33801;
    wire N__33798;
    wire N__33797;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33769;
    wire N__33768;
    wire N__33767;
    wire N__33764;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33756;
    wire N__33753;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33733;
    wire N__33732;
    wire N__33731;
    wire N__33730;
    wire N__33719;
    wire N__33716;
    wire N__33711;
    wire N__33708;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33681;
    wire N__33678;
    wire N__33671;
    wire N__33668;
    wire N__33659;
    wire N__33652;
    wire N__33639;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33631;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33612;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33591;
    wire N__33590;
    wire N__33589;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33560;
    wire N__33557;
    wire N__33552;
    wire N__33551;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33530;
    wire N__33529;
    wire N__33526;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33464;
    wire N__33463;
    wire N__33462;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33455;
    wire N__33454;
    wire N__33453;
    wire N__33452;
    wire N__33451;
    wire N__33450;
    wire N__33447;
    wire N__33446;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33438;
    wire N__33435;
    wire N__33430;
    wire N__33427;
    wire N__33422;
    wire N__33419;
    wire N__33418;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33410;
    wire N__33409;
    wire N__33408;
    wire N__33407;
    wire N__33398;
    wire N__33389;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33385;
    wire N__33384;
    wire N__33383;
    wire N__33380;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33374;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33350;
    wire N__33347;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33326;
    wire N__33319;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33297;
    wire N__33288;
    wire N__33285;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33265;
    wire N__33260;
    wire N__33251;
    wire N__33240;
    wire N__33239;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33230;
    wire N__33229;
    wire N__33224;
    wire N__33223;
    wire N__33222;
    wire N__33221;
    wire N__33220;
    wire N__33219;
    wire N__33218;
    wire N__33217;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33199;
    wire N__33198;
    wire N__33197;
    wire N__33196;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33188;
    wire N__33187;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33175;
    wire N__33164;
    wire N__33163;
    wire N__33162;
    wire N__33161;
    wire N__33160;
    wire N__33159;
    wire N__33158;
    wire N__33157;
    wire N__33156;
    wire N__33155;
    wire N__33152;
    wire N__33147;
    wire N__33144;
    wire N__33143;
    wire N__33142;
    wire N__33141;
    wire N__33140;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33126;
    wire N__33123;
    wire N__33118;
    wire N__33107;
    wire N__33102;
    wire N__33101;
    wire N__33098;
    wire N__33093;
    wire N__33090;
    wire N__33085;
    wire N__33076;
    wire N__33069;
    wire N__33066;
    wire N__33063;
    wire N__33054;
    wire N__33045;
    wire N__33042;
    wire N__33033;
    wire N__33030;
    wire N__33025;
    wire N__33022;
    wire N__33015;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32966;
    wire N__32961;
    wire N__32958;
    wire N__32957;
    wire N__32956;
    wire N__32949;
    wire N__32946;
    wire N__32945;
    wire N__32944;
    wire N__32941;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32909;
    wire N__32904;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32879;
    wire N__32874;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32856;
    wire N__32855;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32831;
    wire N__32826;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32814;
    wire N__32811;
    wire N__32810;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32738;
    wire N__32735;
    wire N__32734;
    wire N__32729;
    wire N__32726;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32701;
    wire N__32698;
    wire N__32693;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32662;
    wire N__32657;
    wire N__32652;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32627;
    wire N__32622;
    wire N__32619;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32611;
    wire N__32608;
    wire N__32603;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32582;
    wire N__32579;
    wire N__32574;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32547;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32535;
    wire N__32534;
    wire N__32529;
    wire N__32526;
    wire N__32525;
    wire N__32524;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32483;
    wire N__32478;
    wire N__32475;
    wire N__32474;
    wire N__32471;
    wire N__32470;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32408;
    wire N__32405;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32385;
    wire N__32384;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32343;
    wire N__32340;
    wire N__32339;
    wire N__32334;
    wire N__32331;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32323;
    wire N__32318;
    wire N__32315;
    wire N__32310;
    wire N__32309;
    wire N__32308;
    wire N__32307;
    wire N__32306;
    wire N__32305;
    wire N__32304;
    wire N__32303;
    wire N__32302;
    wire N__32301;
    wire N__32298;
    wire N__32297;
    wire N__32296;
    wire N__32295;
    wire N__32294;
    wire N__32293;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32285;
    wire N__32284;
    wire N__32283;
    wire N__32282;
    wire N__32279;
    wire N__32278;
    wire N__32277;
    wire N__32276;
    wire N__32275;
    wire N__32274;
    wire N__32273;
    wire N__32270;
    wire N__32269;
    wire N__32268;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32253;
    wire N__32250;
    wire N__32249;
    wire N__32248;
    wire N__32243;
    wire N__32234;
    wire N__32229;
    wire N__32226;
    wire N__32217;
    wire N__32214;
    wire N__32205;
    wire N__32204;
    wire N__32203;
    wire N__32200;
    wire N__32199;
    wire N__32198;
    wire N__32197;
    wire N__32196;
    wire N__32193;
    wire N__32186;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32167;
    wire N__32164;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32125;
    wire N__32120;
    wire N__32107;
    wire N__32104;
    wire N__32097;
    wire N__32094;
    wire N__32087;
    wire N__32082;
    wire N__32073;
    wire N__32070;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31985;
    wire N__31984;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31966;
    wire N__31965;
    wire N__31962;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31903;
    wire N__31898;
    wire N__31887;
    wire N__31884;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31778;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31598;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31583;
    wire N__31582;
    wire N__31581;
    wire N__31578;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31559;
    wire N__31558;
    wire N__31557;
    wire N__31556;
    wire N__31555;
    wire N__31554;
    wire N__31553;
    wire N__31552;
    wire N__31549;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31534;
    wire N__31533;
    wire N__31532;
    wire N__31529;
    wire N__31528;
    wire N__31527;
    wire N__31524;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31501;
    wire N__31494;
    wire N__31489;
    wire N__31484;
    wire N__31477;
    wire N__31464;
    wire N__31463;
    wire N__31462;
    wire N__31461;
    wire N__31460;
    wire N__31457;
    wire N__31456;
    wire N__31455;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31449;
    wire N__31448;
    wire N__31445;
    wire N__31444;
    wire N__31443;
    wire N__31442;
    wire N__31441;
    wire N__31440;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31425;
    wire N__31424;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31406;
    wire N__31399;
    wire N__31396;
    wire N__31395;
    wire N__31394;
    wire N__31393;
    wire N__31390;
    wire N__31385;
    wire N__31382;
    wire N__31375;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31355;
    wire N__31352;
    wire N__31341;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31300;
    wire N__31299;
    wire N__31298;
    wire N__31297;
    wire N__31296;
    wire N__31295;
    wire N__31292;
    wire N__31291;
    wire N__31290;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31258;
    wire N__31257;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31222;
    wire N__31219;
    wire N__31210;
    wire N__31207;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30947;
    wire N__30946;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30925;
    wire N__30922;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30828;
    wire N__30825;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30801;
    wire N__30800;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30792;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30771;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30762;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30754;
    wire N__30753;
    wire N__30750;
    wire N__30749;
    wire N__30748;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30732;
    wire N__30729;
    wire N__30722;
    wire N__30719;
    wire N__30714;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30698;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30683;
    wire N__30682;
    wire N__30681;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30662;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30644;
    wire N__30643;
    wire N__30638;
    wire N__30637;
    wire N__30636;
    wire N__30635;
    wire N__30634;
    wire N__30633;
    wire N__30630;
    wire N__30629;
    wire N__30628;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30605;
    wire N__30600;
    wire N__30595;
    wire N__30592;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30521;
    wire N__30520;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30498;
    wire N__30497;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30479;
    wire N__30478;
    wire N__30471;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30456;
    wire N__30455;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30431;
    wire N__30430;
    wire N__30429;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30406;
    wire N__30403;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30381;
    wire N__30378;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30338;
    wire N__30337;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30291;
    wire N__30290;
    wire N__30289;
    wire N__30288;
    wire N__30287;
    wire N__30286;
    wire N__30285;
    wire N__30284;
    wire N__30283;
    wire N__30282;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30276;
    wire N__30267;
    wire N__30266;
    wire N__30265;
    wire N__30264;
    wire N__30255;
    wire N__30254;
    wire N__30253;
    wire N__30252;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30230;
    wire N__30227;
    wire N__30220;
    wire N__30211;
    wire N__30204;
    wire N__30201;
    wire N__30200;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30179;
    wire N__30174;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30153;
    wire N__30152;
    wire N__30151;
    wire N__30150;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30129;
    wire N__30126;
    wire N__30125;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30099;
    wire N__30096;
    wire N__30095;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30084;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30070;
    wire N__30067;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30036;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29978;
    wire N__29977;
    wire N__29976;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29946;
    wire N__29945;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29916;
    wire N__29913;
    wire N__29912;
    wire N__29907;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29880;
    wire N__29877;
    wire N__29876;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29855;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29819;
    wire N__29818;
    wire N__29817;
    wire N__29816;
    wire N__29815;
    wire N__29814;
    wire N__29813;
    wire N__29810;
    wire N__29797;
    wire N__29796;
    wire N__29795;
    wire N__29794;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29783;
    wire N__29782;
    wire N__29781;
    wire N__29780;
    wire N__29779;
    wire N__29770;
    wire N__29763;
    wire N__29754;
    wire N__29751;
    wire N__29742;
    wire N__29739;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29718;
    wire N__29717;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29699;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29681;
    wire N__29678;
    wire N__29673;
    wire N__29672;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29654;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29627;
    wire N__29624;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29567;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29477;
    wire N__29476;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29442;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29425;
    wire N__29422;
    wire N__29415;
    wire N__29414;
    wire N__29413;
    wire N__29410;
    wire N__29409;
    wire N__29406;
    wire N__29399;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29363;
    wire N__29358;
    wire N__29355;
    wire N__29354;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29277;
    wire N__29276;
    wire N__29275;
    wire N__29272;
    wire N__29263;
    wire N__29258;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29243;
    wire N__29242;
    wire N__29241;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29225;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29198;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29151;
    wire N__29150;
    wire N__29149;
    wire N__29146;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29113;
    wire N__29112;
    wire N__29109;
    wire N__29108;
    wire N__29107;
    wire N__29104;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29089;
    wire N__29088;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29051;
    wire N__29048;
    wire N__29043;
    wire N__29038;
    wire N__29031;
    wire N__29028;
    wire N__29027;
    wire N__29022;
    wire N__29019;
    wire N__29018;
    wire N__29013;
    wire N__29010;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28988;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28964;
    wire N__28961;
    wire N__28960;
    wire N__28957;
    wire N__28956;
    wire N__28953;
    wire N__28946;
    wire N__28943;
    wire N__28938;
    wire N__28935;
    wire N__28934;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28913;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28901;
    wire N__28896;
    wire N__28893;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28880;
    wire N__28877;
    wire N__28872;
    wire N__28871;
    wire N__28868;
    wire N__28863;
    wire N__28862;
    wire N__28861;
    wire N__28860;
    wire N__28859;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28842;
    wire N__28839;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28814;
    wire N__28811;
    wire N__28810;
    wire N__28809;
    wire N__28808;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28796;
    wire N__28795;
    wire N__28794;
    wire N__28791;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28774;
    wire N__28771;
    wire N__28770;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28754;
    wire N__28749;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28733;
    wire N__28730;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28718;
    wire N__28715;
    wire N__28714;
    wire N__28711;
    wire N__28706;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28680;
    wire N__28679;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28671;
    wire N__28670;
    wire N__28667;
    wire N__28666;
    wire N__28663;
    wire N__28658;
    wire N__28651;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28632;
    wire N__28631;
    wire N__28630;
    wire N__28629;
    wire N__28628;
    wire N__28623;
    wire N__28618;
    wire N__28615;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28580;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28550;
    wire N__28549;
    wire N__28548;
    wire N__28547;
    wire N__28546;
    wire N__28545;
    wire N__28544;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28533;
    wire N__28532;
    wire N__28531;
    wire N__28528;
    wire N__28527;
    wire N__28526;
    wire N__28525;
    wire N__28524;
    wire N__28521;
    wire N__28512;
    wire N__28503;
    wire N__28502;
    wire N__28501;
    wire N__28500;
    wire N__28499;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28482;
    wire N__28479;
    wire N__28472;
    wire N__28469;
    wire N__28464;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28436;
    wire N__28433;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28413;
    wire N__28410;
    wire N__28409;
    wire N__28408;
    wire N__28407;
    wire N__28406;
    wire N__28405;
    wire N__28404;
    wire N__28403;
    wire N__28402;
    wire N__28401;
    wire N__28400;
    wire N__28399;
    wire N__28398;
    wire N__28397;
    wire N__28396;
    wire N__28395;
    wire N__28394;
    wire N__28393;
    wire N__28392;
    wire N__28391;
    wire N__28390;
    wire N__28389;
    wire N__28388;
    wire N__28387;
    wire N__28384;
    wire N__28383;
    wire N__28382;
    wire N__28379;
    wire N__28372;
    wire N__28365;
    wire N__28362;
    wire N__28353;
    wire N__28352;
    wire N__28351;
    wire N__28344;
    wire N__28343;
    wire N__28340;
    wire N__28331;
    wire N__28330;
    wire N__28329;
    wire N__28328;
    wire N__28327;
    wire N__28326;
    wire N__28325;
    wire N__28324;
    wire N__28321;
    wire N__28320;
    wire N__28319;
    wire N__28314;
    wire N__28311;
    wire N__28306;
    wire N__28295;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28279;
    wire N__28274;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28260;
    wire N__28259;
    wire N__28258;
    wire N__28257;
    wire N__28254;
    wire N__28249;
    wire N__28242;
    wire N__28241;
    wire N__28240;
    wire N__28235;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28192;
    wire N__28185;
    wire N__28180;
    wire N__28161;
    wire N__28158;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28146;
    wire N__28145;
    wire N__28144;
    wire N__28143;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28125;
    wire N__28116;
    wire N__28115;
    wire N__28114;
    wire N__28113;
    wire N__28112;
    wire N__28111;
    wire N__28108;
    wire N__28107;
    wire N__28104;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28086;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28078;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28028;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28004;
    wire N__28003;
    wire N__27998;
    wire N__27995;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27959;
    wire N__27958;
    wire N__27951;
    wire N__27948;
    wire N__27947;
    wire N__27946;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27908;
    wire N__27903;
    wire N__27900;
    wire N__27899;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27887;
    wire N__27884;
    wire N__27879;
    wire N__27876;
    wire N__27875;
    wire N__27874;
    wire N__27869;
    wire N__27866;
    wire N__27861;
    wire N__27860;
    wire N__27859;
    wire N__27858;
    wire N__27855;
    wire N__27848;
    wire N__27843;
    wire N__27842;
    wire N__27841;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27809;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27782;
    wire N__27779;
    wire N__27778;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27766;
    wire N__27763;
    wire N__27762;
    wire N__27761;
    wire N__27754;
    wire N__27749;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27734;
    wire N__27733;
    wire N__27732;
    wire N__27731;
    wire N__27730;
    wire N__27727;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27645;
    wire N__27642;
    wire N__27641;
    wire N__27640;
    wire N__27637;
    wire N__27632;
    wire N__27627;
    wire N__27626;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27609;
    wire N__27606;
    wire N__27605;
    wire N__27600;
    wire N__27597;
    wire N__27596;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27584;
    wire N__27579;
    wire N__27576;
    wire N__27575;
    wire N__27570;
    wire N__27567;
    wire N__27566;
    wire N__27565;
    wire N__27564;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27552;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27538;
    wire N__27537;
    wire N__27536;
    wire N__27535;
    wire N__27534;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27467;
    wire N__27466;
    wire N__27465;
    wire N__27462;
    wire N__27457;
    wire N__27452;
    wire N__27449;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27393;
    wire N__27390;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27042;
    wire N__27039;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27014;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26996;
    wire N__26995;
    wire N__26992;
    wire N__26985;
    wire N__26982;
    wire N__26981;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26939;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26915;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26861;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26819;
    wire N__26814;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26777;
    wire N__26776;
    wire N__26775;
    wire N__26774;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26762;
    wire N__26757;
    wire N__26748;
    wire N__26747;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26734;
    wire N__26733;
    wire N__26732;
    wire N__26725;
    wire N__26720;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26693;
    wire N__26692;
    wire N__26691;
    wire N__26682;
    wire N__26681;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26673;
    wire N__26672;
    wire N__26671;
    wire N__26670;
    wire N__26669;
    wire N__26666;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26654;
    wire N__26645;
    wire N__26640;
    wire N__26635;
    wire N__26628;
    wire N__26627;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26553;
    wire N__26552;
    wire N__26549;
    wire N__26548;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26534;
    wire N__26533;
    wire N__26532;
    wire N__26531;
    wire N__26530;
    wire N__26529;
    wire N__26528;
    wire N__26527;
    wire N__26526;
    wire N__26525;
    wire N__26524;
    wire N__26523;
    wire N__26522;
    wire N__26517;
    wire N__26506;
    wire N__26489;
    wire N__26474;
    wire N__26473;
    wire N__26472;
    wire N__26471;
    wire N__26468;
    wire N__26467;
    wire N__26466;
    wire N__26461;
    wire N__26460;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26452;
    wire N__26439;
    wire N__26436;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26351;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26295;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26287;
    wire N__26282;
    wire N__26279;
    wire N__26278;
    wire N__26277;
    wire N__26276;
    wire N__26271;
    wire N__26270;
    wire N__26267;
    wire N__26266;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26262;
    wire N__26259;
    wire N__26258;
    wire N__26257;
    wire N__26256;
    wire N__26255;
    wire N__26254;
    wire N__26253;
    wire N__26252;
    wire N__26251;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26233;
    wire N__26224;
    wire N__26223;
    wire N__26222;
    wire N__26221;
    wire N__26216;
    wire N__26209;
    wire N__26202;
    wire N__26193;
    wire N__26190;
    wire N__26185;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26136;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26108;
    wire N__26105;
    wire N__26104;
    wire N__26103;
    wire N__26102;
    wire N__26091;
    wire N__26090;
    wire N__26089;
    wire N__26088;
    wire N__26087;
    wire N__26086;
    wire N__26085;
    wire N__26082;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26070;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26046;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26031;
    wire N__26028;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26017;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26005;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25991;
    wire N__25990;
    wire N__25989;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25981;
    wire N__25980;
    wire N__25979;
    wire N__25978;
    wire N__25977;
    wire N__25976;
    wire N__25975;
    wire N__25974;
    wire N__25971;
    wire N__25970;
    wire N__25967;
    wire N__25966;
    wire N__25965;
    wire N__25964;
    wire N__25963;
    wire N__25962;
    wire N__25961;
    wire N__25960;
    wire N__25959;
    wire N__25958;
    wire N__25955;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25937;
    wire N__25934;
    wire N__25929;
    wire N__25926;
    wire N__25915;
    wire N__25904;
    wire N__25903;
    wire N__25902;
    wire N__25899;
    wire N__25898;
    wire N__25897;
    wire N__25896;
    wire N__25893;
    wire N__25884;
    wire N__25883;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25869;
    wire N__25858;
    wire N__25857;
    wire N__25856;
    wire N__25855;
    wire N__25854;
    wire N__25853;
    wire N__25850;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25832;
    wire N__25827;
    wire N__25816;
    wire N__25811;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25712;
    wire N__25711;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25683;
    wire N__25680;
    wire N__25679;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25635;
    wire N__25632;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25560;
    wire N__25557;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25542;
    wire N__25541;
    wire N__25538;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25508;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25490;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25463;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25355;
    wire N__25352;
    wire N__25351;
    wire N__25348;
    wire N__25347;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25333;
    wire N__25326;
    wire N__25325;
    wire N__25322;
    wire N__25321;
    wire N__25318;
    wire N__25317;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25303;
    wire N__25296;
    wire N__25295;
    wire N__25292;
    wire N__25291;
    wire N__25288;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25262;
    wire N__25261;
    wire N__25256;
    wire N__25253;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25198;
    wire N__25197;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25013;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24991;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24961;
    wire N__24958;
    wire N__24953;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24938;
    wire N__24935;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24923;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24905;
    wire N__24904;
    wire N__24901;
    wire N__24896;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24878;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24716;
    wire N__24715;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24698;
    wire N__24695;
    wire N__24694;
    wire N__24691;
    wire N__24684;
    wire N__24681;
    wire N__24680;
    wire N__24679;
    wire N__24674;
    wire N__24671;
    wire N__24666;
    wire N__24665;
    wire N__24664;
    wire N__24663;
    wire N__24662;
    wire N__24659;
    wire N__24650;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24609;
    wire N__24606;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24545;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24522;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24510;
    wire N__24507;
    wire N__24506;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24494;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24484;
    wire N__24479;
    wire N__24476;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24435;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24423;
    wire N__24420;
    wire N__24419;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24404;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24335;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24264;
    wire N__24263;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24194;
    wire N__24191;
    wire N__24190;
    wire N__24187;
    wire N__24186;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24172;
    wire N__24165;
    wire N__24164;
    wire N__24161;
    wire N__24160;
    wire N__24157;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24098;
    wire N__24095;
    wire N__24094;
    wire N__24091;
    wire N__24090;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24076;
    wire N__24069;
    wire N__24068;
    wire N__24065;
    wire N__24064;
    wire N__24061;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24020;
    wire N__24017;
    wire N__24016;
    wire N__24013;
    wire N__24012;
    wire N__24009;
    wire N__24004;
    wire N__24001;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23986;
    wire N__23983;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23945;
    wire N__23942;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23915;
    wire N__23912;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23873;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23765;
    wire N__23762;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23750;
    wire N__23749;
    wire N__23748;
    wire N__23747;
    wire N__23746;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23730;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23640;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23625;
    wire N__23622;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23607;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23472;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23457;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23427;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23415;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23400;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23372;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23310;
    wire N__23307;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23240;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23225;
    wire N__23222;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23210;
    wire N__23205;
    wire N__23202;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23159;
    wire N__23154;
    wire N__23153;
    wire N__23152;
    wire N__23151;
    wire N__23150;
    wire N__23149;
    wire N__23148;
    wire N__23147;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23072;
    wire N__23069;
    wire N__23068;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23049;
    wire N__23040;
    wire N__23037;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23022;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__22999;
    wire N__22992;
    wire N__22989;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22974;
    wire N__22971;
    wire N__22970;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22922;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22901;
    wire N__22900;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22845;
    wire N__22842;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22827;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22779;
    wire N__22778;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22766;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22751;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22739;
    wire N__22736;
    wire N__22735;
    wire N__22732;
    wire N__22727;
    wire N__22724;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22625;
    wire N__22624;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22618;
    wire N__22617;
    wire N__22616;
    wire N__22615;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22605;
    wire N__22604;
    wire N__22603;
    wire N__22602;
    wire N__22601;
    wire N__22590;
    wire N__22579;
    wire N__22574;
    wire N__22565;
    wire N__22552;
    wire N__22543;
    wire N__22542;
    wire N__22541;
    wire N__22540;
    wire N__22539;
    wire N__22538;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22472;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22446;
    wire N__22445;
    wire N__22444;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22430;
    wire N__22429;
    wire N__22426;
    wire N__22421;
    wire N__22416;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22404;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22344;
    wire N__22343;
    wire N__22342;
    wire N__22341;
    wire N__22340;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22325;
    wire N__22320;
    wire N__22315;
    wire N__22314;
    wire N__22309;
    wire N__22300;
    wire N__22297;
    wire N__22290;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22266;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22093;
    wire N__22092;
    wire N__22091;
    wire N__22088;
    wire N__22081;
    wire N__22078;
    wire N__22073;
    wire N__22068;
    wire N__22067;
    wire N__22064;
    wire N__22063;
    wire N__22060;
    wire N__22059;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22045;
    wire N__22038;
    wire N__22037;
    wire N__22034;
    wire N__22033;
    wire N__22030;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21989;
    wire N__21986;
    wire N__21985;
    wire N__21982;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21876;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21809;
    wire N__21806;
    wire N__21805;
    wire N__21802;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21753;
    wire N__21750;
    wire N__21745;
    wire N__21742;
    wire N__21735;
    wire N__21732;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21618;
    wire N__21615;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21537;
    wire N__21534;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21522;
    wire N__21519;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21504;
    wire N__21501;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21471;
    wire N__21468;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21456;
    wire N__21453;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21441;
    wire N__21438;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21395;
    wire N__21394;
    wire N__21391;
    wire N__21386;
    wire N__21381;
    wire N__21380;
    wire N__21379;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21359;
    wire N__21358;
    wire N__21351;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21339;
    wire N__21336;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21328;
    wire N__21325;
    wire N__21320;
    wire N__21315;
    wire N__21314;
    wire N__21309;
    wire N__21308;
    wire N__21307;
    wire N__21304;
    wire N__21299;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21263;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21240;
    wire N__21237;
    wire N__21236;
    wire N__21233;
    wire N__21228;
    wire N__21225;
    wire N__21224;
    wire N__21221;
    wire N__21216;
    wire N__21213;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21194;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21129;
    wire N__21126;
    wire N__21125;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21110;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21084;
    wire N__21083;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21050;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20975;
    wire N__20974;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20937;
    wire N__20934;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20864;
    wire N__20863;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20822;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20804;
    wire N__20803;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20754;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20726;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20712;
    wire N__20709;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20684;
    wire N__20683;
    wire N__20680;
    wire N__20675;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20607;
    wire N__20604;
    wire N__20603;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20580;
    wire N__20577;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20568;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20554;
    wire N__20547;
    wire N__20546;
    wire N__20543;
    wire N__20542;
    wire N__20539;
    wire N__20532;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20486;
    wire N__20485;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20477;
    wire N__20476;
    wire N__20475;
    wire N__20470;
    wire N__20465;
    wire N__20462;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20424;
    wire N__20423;
    wire N__20420;
    wire N__20419;
    wire N__20416;
    wire N__20415;
    wire N__20412;
    wire N__20407;
    wire N__20404;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20378;
    wire N__20375;
    wire N__20374;
    wire N__20371;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20188;
    wire N__20185;
    wire N__20184;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20170;
    wire N__20163;
    wire N__20162;
    wire N__20159;
    wire N__20158;
    wire N__20155;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20120;
    wire N__20117;
    wire N__20116;
    wire N__20113;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20084;
    wire N__20081;
    wire N__20074;
    wire N__20071;
    wire N__20064;
    wire N__20063;
    wire N__20062;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20055;
    wire N__20054;
    wire N__20053;
    wire N__20052;
    wire N__20051;
    wire N__20050;
    wire N__20043;
    wire N__20034;
    wire N__20031;
    wire N__20022;
    wire N__20015;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20007;
    wire N__20004;
    wire N__19999;
    wire N__19992;
    wire N__19987;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19970;
    wire N__19967;
    wire N__19966;
    wire N__19963;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19925;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19907;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19895;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19805;
    wire N__19804;
    wire N__19803;
    wire N__19802;
    wire N__19799;
    wire N__19798;
    wire N__19797;
    wire N__19786;
    wire N__19783;
    wire N__19782;
    wire N__19781;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19777;
    wire N__19776;
    wire N__19775;
    wire N__19774;
    wire N__19773;
    wire N__19772;
    wire N__19771;
    wire N__19770;
    wire N__19769;
    wire N__19768;
    wire N__19767;
    wire N__19766;
    wire N__19765;
    wire N__19764;
    wire N__19763;
    wire N__19762;
    wire N__19759;
    wire N__19754;
    wire N__19749;
    wire N__19746;
    wire N__19735;
    wire N__19726;
    wire N__19715;
    wire N__19706;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19684;
    wire N__19681;
    wire N__19676;
    wire N__19671;
    wire N__19668;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19625;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19613;
    wire N__19610;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19595;
    wire N__19594;
    wire N__19591;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19559;
    wire N__19558;
    wire N__19557;
    wire N__19550;
    wire N__19549;
    wire N__19548;
    wire N__19547;
    wire N__19544;
    wire N__19543;
    wire N__19542;
    wire N__19541;
    wire N__19538;
    wire N__19531;
    wire N__19530;
    wire N__19527;
    wire N__19526;
    wire N__19525;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19510;
    wire N__19509;
    wire N__19508;
    wire N__19507;
    wire N__19506;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19481;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19469;
    wire N__19468;
    wire N__19467;
    wire N__19464;
    wire N__19463;
    wire N__19462;
    wire N__19461;
    wire N__19460;
    wire N__19459;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19453;
    wire N__19446;
    wire N__19445;
    wire N__19444;
    wire N__19437;
    wire N__19434;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19416;
    wire N__19409;
    wire N__19402;
    wire N__19397;
    wire N__19392;
    wire N__19385;
    wire N__19382;
    wire N__19377;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19357;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19277;
    wire N__19276;
    wire N__19275;
    wire N__19274;
    wire N__19273;
    wire N__19272;
    wire N__19271;
    wire N__19266;
    wire N__19263;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19253;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19243;
    wire N__19242;
    wire N__19241;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19224;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19210;
    wire N__19207;
    wire N__19200;
    wire N__19195;
    wire N__19190;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19172;
    wire N__19159;
    wire N__19146;
    wire N__19145;
    wire N__19142;
    wire N__19141;
    wire N__19138;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19109;
    wire N__19106;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19082;
    wire N__19081;
    wire N__19080;
    wire N__19077;
    wire N__19074;
    wire N__19073;
    wire N__19072;
    wire N__19071;
    wire N__19070;
    wire N__19069;
    wire N__19068;
    wire N__19065;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19061;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19049;
    wire N__19044;
    wire N__19037;
    wire N__19026;
    wire N__19025;
    wire N__19022;
    wire N__19021;
    wire N__19020;
    wire N__19019;
    wire N__19014;
    wire N__19009;
    wire N__19004;
    wire N__18993;
    wire N__18988;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18957;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18935;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18893;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18843;
    wire N__18842;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18818;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18800;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18779;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18744;
    wire N__18743;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18725;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18698;
    wire N__18695;
    wire N__18694;
    wire N__18691;
    wire N__18684;
    wire N__18681;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18669;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18648;
    wire N__18645;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18633;
    wire N__18630;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18615;
    wire N__18612;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18600;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18585;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18567;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18552;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18537;
    wire N__18534;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18522;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18504;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18474;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18456;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18441;
    wire N__18438;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18426;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18414;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18393;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18381;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18348;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18333;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18321;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18303;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18291;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18270;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18246;
    wire N__18245;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18222;
    wire N__18221;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18170;
    wire N__18165;
    wire N__18162;
    wire N__18161;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18141;
    wire N__18138;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18111;
    wire N__18110;
    wire N__18107;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18081;
    wire N__18078;
    wire N__18077;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18054;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18032;
    wire N__18029;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18008;
    wire N__18005;
    wire N__18000;
    wire N__17999;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17976;
    wire N__17973;
    wire N__17972;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17945;
    wire N__17942;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17927;
    wire N__17924;
    wire N__17919;
    wire N__17916;
    wire N__17915;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17886;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17880;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17864;
    wire N__17861;
    wire N__17860;
    wire N__17859;
    wire N__17856;
    wire N__17855;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17839;
    wire N__17836;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17805;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17787;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17775;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17754;
    wire N__17753;
    wire N__17750;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17732;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17717;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17696;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17681;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17663;
    wire N__17662;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17610;
    wire N__17607;
    wire N__17606;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17588;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17570;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17541;
    wire N__17538;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17511;
    wire N__17510;
    wire N__17505;
    wire N__17502;
    wire N__17499;
    wire N__17498;
    wire N__17495;
    wire N__17494;
    wire N__17493;
    wire N__17492;
    wire N__17491;
    wire N__17490;
    wire N__17489;
    wire N__17488;
    wire N__17487;
    wire N__17480;
    wire N__17479;
    wire N__17478;
    wire N__17477;
    wire N__17476;
    wire N__17475;
    wire N__17464;
    wire N__17459;
    wire N__17456;
    wire N__17445;
    wire N__17440;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17420;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17397;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17346;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17327;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17271;
    wire N__17270;
    wire N__17269;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17250;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17238;
    wire N__17235;
    wire N__17234;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17217;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17172;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17136;
    wire N__17133;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17097;
    wire N__17096;
    wire N__17091;
    wire N__17088;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire N__17070;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17046;
    wire N__17045;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17012;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__17001;
    wire N__16994;
    wire N__16993;
    wire N__16992;
    wire N__16991;
    wire N__16990;
    wire N__16989;
    wire N__16988;
    wire N__16987;
    wire N__16986;
    wire N__16985;
    wire N__16984;
    wire N__16983;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16968;
    wire N__16959;
    wire N__16948;
    wire N__16947;
    wire N__16946;
    wire N__16945;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16939;
    wire N__16938;
    wire N__16937;
    wire N__16936;
    wire N__16935;
    wire N__16924;
    wire N__16917;
    wire N__16916;
    wire N__16915;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16893;
    wire N__16888;
    wire N__16881;
    wire N__16866;
    wire N__16865;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16815;
    wire N__16812;
    wire N__16811;
    wire N__16810;
    wire N__16809;
    wire N__16806;
    wire N__16801;
    wire N__16798;
    wire N__16791;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16769;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16754;
    wire N__16753;
    wire N__16748;
    wire N__16745;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16706;
    wire N__16705;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16686;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16664;
    wire N__16659;
    wire N__16656;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16644;
    wire N__16641;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16629;
    wire N__16628;
    wire N__16625;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16610;
    wire N__16607;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16592;
    wire N__16589;
    wire N__16584;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16559;
    wire N__16556;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16539;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16496;
    wire N__16495;
    wire N__16492;
    wire N__16487;
    wire N__16484;
    wire N__16479;
    wire N__16478;
    wire N__16475;
    wire N__16474;
    wire N__16469;
    wire N__16466;
    wire N__16461;
    wire N__16458;
    wire N__16457;
    wire N__16452;
    wire N__16449;
    wire N__16446;
    wire N__16445;
    wire N__16444;
    wire N__16439;
    wire N__16436;
    wire N__16431;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16403;
    wire N__16402;
    wire N__16397;
    wire N__16394;
    wire N__16389;
    wire N__16386;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16374;
    wire N__16373;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16355;
    wire N__16354;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16337;
    wire N__16336;
    wire N__16333;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16311;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16262;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16247;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16226;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16199;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16019;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15984;
    wire N__15981;
    wire N__15980;
    wire N__15977;
    wire N__15972;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15881;
    wire N__15876;
    wire N__15873;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15845;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15806;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15752;
    wire N__15747;
    wire VCCG0;
    wire GNDG0;
    wire \b2v_inst36.countZ0Z_10_cascade_ ;
    wire \b2v_inst36.count_2_10 ;
    wire \b2v_inst36.count_rst_9 ;
    wire \b2v_inst36.count_rst_9_cascade_ ;
    wire \b2v_inst36.un2_count_1_axb_5_cascade_ ;
    wire \b2v_inst36.count_2_5 ;
    wire \b2v_inst36.count_rst_7_cascade_ ;
    wire \b2v_inst36.countZ0Z_6_cascade_ ;
    wire \b2v_inst36.count_2_4 ;
    wire \b2v_inst36.countZ0Z_11_cascade_ ;
    wire \b2v_inst36.count_2_11 ;
    wire \b2v_inst36.count_2_6 ;
    wire \b2v_inst36.count_rst_6 ;
    wire \b2v_inst36.count_rst_6_cascade_ ;
    wire \b2v_inst36.un2_count_1_axb_8_cascade_ ;
    wire \b2v_inst36.count_2_8 ;
    wire \b2v_inst36.count_rst_4 ;
    wire \b2v_inst36.count_rst_3 ;
    wire \b2v_inst36.count_rst_13 ;
    wire \b2v_inst36.count_rst_13_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_1 ;
    wire \b2v_inst36.un12_clk_100khz_0_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_2 ;
    wire \b2v_inst36.un12_clk_100khz_7 ;
    wire \b2v_inst36.un12_clk_100khz_12_cascade_ ;
    wire \b2v_inst36.N_1_i_cascade_ ;
    wire \b2v_inst36.count_2_0 ;
    wire \b2v_inst36.count_rst_14 ;
    wire \b2v_inst36.countZ0Z_0_cascade_ ;
    wire \b2v_inst36.count_2_1 ;
    wire \b2v_inst16.count_rst_0_cascade_ ;
    wire \b2v_inst16.countZ0Z_11_cascade_ ;
    wire \b2v_inst16.count_4_11 ;
    wire \b2v_inst16.count_rst_9_cascade_ ;
    wire \b2v_inst16.countZ0Z_4_cascade_ ;
    wire \b2v_inst16.count_4_4 ;
    wire \b2v_inst16.countZ0Z_3_cascade_ ;
    wire \b2v_inst16.count_4_3 ;
    wire \b2v_inst16.count_4_i_a3_9_0 ;
    wire \b2v_inst16.count_4_i_a3_8_0_cascade_ ;
    wire \b2v_inst16.count_4_i_a3_10_0 ;
    wire \b2v_inst16.N_414_cascade_ ;
    wire \b2v_inst16.N_416_cascade_ ;
    wire \b2v_inst16.count_rst_8 ;
    wire \b2v_inst16.count_RNIE4RF_2Z0Z_1_cascade_ ;
    wire \b2v_inst16.count_rst_5_cascade_ ;
    wire \b2v_inst16.N_414 ;
    wire \b2v_inst16.countZ0Z_0_cascade_ ;
    wire \b2v_inst16.count_4_0 ;
    wire \b2v_inst16.countZ0Z_1 ;
    wire \b2v_inst16.count_4_i_a3_7_0 ;
    wire \b2v_inst16.count_RNIE4RF_2Z0Z_1 ;
    wire \b2v_inst16.count_4_1 ;
    wire \b2v_inst16.countZ0Z_7_cascade_ ;
    wire \b2v_inst16.count_4_7 ;
    wire \b2v_inst16.count_rst_10_cascade_ ;
    wire \b2v_inst16.countZ0Z_5_cascade_ ;
    wire \b2v_inst16.count_4_5 ;
    wire \b2v_inst16.countZ0Z_8_cascade_ ;
    wire \b2v_inst16.count_4_8 ;
    wire \b2v_inst16.count_rst_12 ;
    wire \b2v_inst16.curr_state_7_0_1_cascade_ ;
    wire vddq_ok;
    wire \b2v_inst16.N_208_0_cascade_ ;
    wire \b2v_inst16.curr_state_RNIBO6I1Z0Z_0_cascade_ ;
    wire \b2v_inst16.curr_state_2_1 ;
    wire \b2v_inst16.curr_state_2_0 ;
    wire \b2v_inst11.count_0_7 ;
    wire bfn_1_11_0_;
    wire \b2v_inst11.un1_count_cry_1_cZ0 ;
    wire \b2v_inst11.un1_count_cry_2_cZ0 ;
    wire \b2v_inst11.un1_count_cry_3 ;
    wire \b2v_inst11.un1_count_cry_4 ;
    wire \b2v_inst11.un1_count_cry_5 ;
    wire \b2v_inst11.count_1_7 ;
    wire \b2v_inst11.un1_count_cry_6 ;
    wire \b2v_inst11.un1_count_cry_7 ;
    wire \b2v_inst11.un1_count_cry_8 ;
    wire bfn_1_12_0_;
    wire \b2v_inst11.un1_count_cry_9 ;
    wire \b2v_inst11.un1_count_cry_10 ;
    wire \b2v_inst11.un1_count_cry_11 ;
    wire \b2v_inst11.un1_count_cry_12 ;
    wire \b2v_inst11.un1_count_cry_13 ;
    wire \b2v_inst11.un1_count_cry_14 ;
    wire \b2v_inst11.count_1_5 ;
    wire \b2v_inst11.count_0_5 ;
    wire \b2v_inst11.count_1_14 ;
    wire \b2v_inst11.count_0_14 ;
    wire \b2v_inst11.count_1_6 ;
    wire \b2v_inst11.count_0_6 ;
    wire \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ;
    wire \b2v_inst11.count_0_15 ;
    wire bfn_1_14_0_;
    wire \b2v_inst11.un85_clk_100khz_0_cry_0 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_1 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_2 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_3 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_4 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_5 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_6 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_7 ;
    wire bfn_1_15_0_;
    wire \b2v_inst11.un85_clk_100khz_0_cry_8 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_9 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_10 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_11 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_12 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_13 ;
    wire \b2v_inst11.un85_clk_100khz_0_cry_14 ;
    wire \b2v_inst11.un85_clk_100khz0 ;
    wire bfn_1_16_0_;
    wire \b2v_inst36.count_rst_12_cascade_ ;
    wire \b2v_inst36.count_rst_12 ;
    wire \b2v_inst36.countZ0Z_3_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_3 ;
    wire \b2v_inst36.count_rst_11 ;
    wire \b2v_inst36.count_2_2 ;
    wire \b2v_inst36.count_2_3 ;
    wire \b2v_inst36.count_2_7 ;
    wire \b2v_inst36.un2_count_1_axb_1 ;
    wire bfn_2_2_0_;
    wire \b2v_inst36.un2_count_1_axb_2 ;
    wire \b2v_inst36.un2_count_1_cry_1_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_1 ;
    wire \b2v_inst36.countZ0Z_3 ;
    wire \b2v_inst36.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_2 ;
    wire \b2v_inst36.un2_count_1_axb_4 ;
    wire \b2v_inst36.count_rst_10 ;
    wire \b2v_inst36.un2_count_1_cry_3 ;
    wire \b2v_inst36.un2_count_1_axb_5 ;
    wire \b2v_inst36.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_4 ;
    wire \b2v_inst36.un2_count_1_axb_6 ;
    wire \b2v_inst36.un2_count_1_cry_5_c_RNIE2FZ0Z8 ;
    wire \b2v_inst36.un2_count_1_cry_5 ;
    wire \b2v_inst36.countZ0Z_7 ;
    wire \b2v_inst36.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_6 ;
    wire \b2v_inst36.un2_count_1_axb_8 ;
    wire \b2v_inst36.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_7 ;
    wire \b2v_inst36.un2_count_1_cry_8 ;
    wire bfn_2_3_0_;
    wire \b2v_inst36.countZ0Z_10 ;
    wire \b2v_inst36.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_9 ;
    wire \b2v_inst36.countZ0Z_11 ;
    wire \b2v_inst36.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_10 ;
    wire \b2v_inst36.un2_count_1_cry_11 ;
    wire \b2v_inst36.un2_count_1_cry_12 ;
    wire \b2v_inst36.un2_count_1_cry_13 ;
    wire \b2v_inst36.un2_count_1_cry_14 ;
    wire \b2v_inst36.un2_count_1_axb_9 ;
    wire \b2v_inst36.count_2_12 ;
    wire \b2v_inst36.count_rst_2 ;
    wire \b2v_inst36.countZ0Z_12 ;
    wire \b2v_inst36.count_rst_5 ;
    wire \b2v_inst36.countZ0Z_12_cascade_ ;
    wire \b2v_inst36.count_2_9 ;
    wire \b2v_inst36.un12_clk_100khz_6 ;
    wire \b2v_inst36.countZ0Z_14 ;
    wire \b2v_inst36.countZ0Z_14_cascade_ ;
    wire \b2v_inst36.countZ0Z_0 ;
    wire \b2v_inst36.un12_clk_100khz_10 ;
    wire \b2v_inst36.count_2_13 ;
    wire \b2v_inst36.count_rst_1 ;
    wire \b2v_inst36.countZ0Z_13 ;
    wire \b2v_inst36.count_rst_0 ;
    wire \b2v_inst36.count_2_14 ;
    wire \b2v_inst36.curr_state_RNINSDSZ0Z_0 ;
    wire \b2v_inst36.count_rst ;
    wire \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_ ;
    wire \b2v_inst36.count_2_15 ;
    wire \b2v_inst36.countZ0Z_15 ;
    wire \b2v_inst16.count_en_cascade_ ;
    wire \b2v_inst16.un4_count_1_axb_1 ;
    wire \b2v_inst16.countZ0Z_0 ;
    wire bfn_2_6_0_;
    wire \b2v_inst16.countZ0Z_2 ;
    wire \b2v_inst16.un4_count_1_cry_1 ;
    wire \b2v_inst16.countZ0Z_3 ;
    wire \b2v_inst16.un4_count_1_cry_2_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_2 ;
    wire \b2v_inst16.countZ0Z_4 ;
    wire \b2v_inst16.un4_count_1_cry_3_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_3 ;
    wire \b2v_inst16.countZ0Z_5 ;
    wire \b2v_inst16.un4_count_1_cry_4_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_4 ;
    wire \b2v_inst16.countZ0Z_6 ;
    wire \b2v_inst16.un4_count_1_cry_5 ;
    wire \b2v_inst16.countZ0Z_7 ;
    wire \b2v_inst16.un4_count_1_cry_6_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_6 ;
    wire \b2v_inst16.un4_count_1_cry_7 ;
    wire \b2v_inst16.un4_count_1_cry_8 ;
    wire bfn_2_7_0_;
    wire \b2v_inst16.un4_count_1_cry_9 ;
    wire \b2v_inst16.countZ0Z_11 ;
    wire \b2v_inst16.un4_count_1_cry_10_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_10 ;
    wire \b2v_inst16.un4_count_1_cry_11 ;
    wire \b2v_inst16.un4_count_1_cry_12 ;
    wire \b2v_inst16.un4_count_1_cry_13 ;
    wire \b2v_inst16.un4_count_1_cry_14 ;
    wire \b2v_inst16.countZ0Z_12 ;
    wire \b2v_inst16.un4_count_1_cry_7_THRU_CO ;
    wire \b2v_inst16.countZ0Z_8 ;
    wire \b2v_inst16.count_rst_13 ;
    wire \b2v_inst16.count_rst_14_cascade_ ;
    wire \b2v_inst16.countZ0Z_9 ;
    wire \b2v_inst16.un4_count_1_cry_8_THRU_CO ;
    wire \b2v_inst16.countZ0Z_9_cascade_ ;
    wire \b2v_inst16.N_416 ;
    wire \b2v_inst16.count_4_9 ;
    wire \b2v_inst16.count_4_10 ;
    wire \b2v_inst16.count_rst ;
    wire \b2v_inst16.countZ0Z_10 ;
    wire \b2v_inst16.count_rst_1 ;
    wire \b2v_inst16.count_4_12 ;
    wire \b2v_inst11.curr_state_3_0_cascade_ ;
    wire \b2v_inst11.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJZ0Z62 ;
    wire \b2v_inst11.curr_state_4_0 ;
    wire \b2v_inst11.count_0_0 ;
    wire \b2v_inst11.countZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_1_1_cascade_ ;
    wire CONSTANT_ONE_NET_cascade_;
    wire \b2v_inst11.N_5852_i ;
    wire \b2v_inst11.countZ0Z_1 ;
    wire \b2v_inst11.count_0_1 ;
    wire \b2v_inst11.count_0_8 ;
    wire \b2v_inst11.count_1_8 ;
    wire \b2v_inst11.count_1_9 ;
    wire \b2v_inst11.count_0_9 ;
    wire \b2v_inst11.count_1_10 ;
    wire \b2v_inst11.count_0_10 ;
    wire \b2v_inst11.count_1_11 ;
    wire \b2v_inst11.count_0_11 ;
    wire \b2v_inst11.count_1_2 ;
    wire \b2v_inst11.count_0_2 ;
    wire \b2v_inst11.count_1_12 ;
    wire \b2v_inst11.count_0_12 ;
    wire \b2v_inst11.count_1_3 ;
    wire \b2v_inst11.count_0_3 ;
    wire \b2v_inst11.count_1_13 ;
    wire \b2v_inst11.count_0_13 ;
    wire \b2v_inst11.count_1_4 ;
    wire \b2v_inst11.count_0_4 ;
    wire \b2v_inst11.countZ0Z_2 ;
    wire \b2v_inst11.countZ0Z_3 ;
    wire \b2v_inst11.countZ0Z_4 ;
    wire \b2v_inst11.countZ0Z_7 ;
    wire \b2v_inst11.countZ0Z_6 ;
    wire \b2v_inst11.un79_clk_100khzlt6_cascade_ ;
    wire \b2v_inst11.countZ0Z_5 ;
    wire \b2v_inst11.countZ0Z_10 ;
    wire \b2v_inst11.countZ0Z_12 ;
    wire \b2v_inst11.countZ0Z_11 ;
    wire \b2v_inst11.countZ0Z_13 ;
    wire \b2v_inst11.countZ0Z_14 ;
    wire \b2v_inst11.un79_clk_100khzlto15_5_cascade_ ;
    wire \b2v_inst11.countZ0Z_15 ;
    wire \b2v_inst11.un79_clk_100khzlto15_3 ;
    wire \b2v_inst11.countZ0Z_8 ;
    wire \b2v_inst11.un79_clk_100khzlto15_7_cascade_ ;
    wire \b2v_inst11.countZ0Z_9 ;
    wire \b2v_inst11.count_RNIZ0Z_8 ;
    wire \b2v_inst11.curr_stateZ0Z_0 ;
    wire \b2v_inst11.count_RNIZ0Z_8_cascade_ ;
    wire \b2v_inst11.curr_state_3_i_m2_0_rep1_1 ;
    wire \b2v_inst11.N_5853_i ;
    wire \b2v_inst11.un85_clk_100khz_0 ;
    wire bfn_2_14_0_;
    wire \b2v_inst11.N_5854_i ;
    wire \b2v_inst11.un85_clk_100khz_0_0 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_1 ;
    wire \b2v_inst11.N_5855_i ;
    wire \b2v_inst11.un85_clk_100khz_0_1 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_2 ;
    wire \b2v_inst11.N_5856_i ;
    wire \b2v_inst11.un85_clk_100khz_0_2 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_3 ;
    wire \b2v_inst11.N_5857_i ;
    wire \b2v_inst11.un85_clk_100khz_0_3 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_4 ;
    wire \b2v_inst11.N_5858_i ;
    wire \b2v_inst11.un85_clk_100khz_0_4 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_5 ;
    wire \b2v_inst11.N_5859_i ;
    wire \b2v_inst11.un85_clk_100khz_0_5 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_6 ;
    wire \b2v_inst11.N_5860_i ;
    wire \b2v_inst11.un85_clk_100khz_0_6 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_7 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_8 ;
    wire \b2v_inst11.N_5861_i ;
    wire \b2v_inst11.un85_clk_100khz_0_7 ;
    wire bfn_2_15_0_;
    wire \b2v_inst11.N_5862_i ;
    wire \b2v_inst11.un85_clk_100khz_1_8 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_9 ;
    wire \b2v_inst11.N_5863_i ;
    wire \b2v_inst11.un85_clk_100khz_1_9 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_10 ;
    wire \b2v_inst11.N_5864_i ;
    wire \b2v_inst11.un85_clk_100khz_1_10 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_11 ;
    wire \b2v_inst11.N_5865_i ;
    wire \b2v_inst11.un85_clk_100khz_1_11 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_12 ;
    wire \b2v_inst11.N_5866_i ;
    wire \b2v_inst11.un85_clk_100khz_1_12 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_13 ;
    wire \b2v_inst11.N_5867_i ;
    wire \b2v_inst11.un85_clk_100khz_1_13 ;
    wire \b2v_inst11.un85_clk_100khz_1_cry_14 ;
    wire \b2v_inst11.un85_clk_100khz1 ;
    wire bfn_2_16_0_;
    wire \b2v_inst11.mult1_un103_sum_cry_2 ;
    wire \b2v_inst11.mult1_un103_sum_cry_3 ;
    wire \b2v_inst11.mult1_un103_sum_cry_4 ;
    wire \b2v_inst11.mult1_un103_sum_cry_5 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6 ;
    wire \b2v_inst11.mult1_un103_sum_cry_7 ;
    wire \b2v_inst11.mult1_un96_sum_i_0_8 ;
    wire \b2v_inst200.un25_clk_100khz_1_cascade_ ;
    wire \b2v_inst200.un2_count_1_axb_1_cascade_ ;
    wire \b2v_inst200.count_RNIZ0Z_1 ;
    wire \b2v_inst200.countZ0Z_16 ;
    wire \b2v_inst200.un25_clk_100khz_0 ;
    wire \b2v_inst200.count_3_1 ;
    wire \b2v_inst200.un25_clk_100khz_3_cascade_ ;
    wire \b2v_inst200.count_3_3 ;
    wire \b2v_inst200.un25_clk_100khz_2 ;
    wire \b2v_inst200.count_3_13 ;
    wire \b2v_inst200.un25_clk_100khz_5 ;
    wire \b2v_inst200.count_3_12 ;
    wire \b2v_inst200.count_3_9 ;
    wire \b2v_inst200.countZ0Z_12_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_4 ;
    wire \b2v_inst200.count_3_5 ;
    wire \b2v_inst16.countZ0Z_15 ;
    wire \b2v_inst16.count_rst_4 ;
    wire \b2v_inst16.count_4_15 ;
    wire \b2v_inst16.countZ0Z_13 ;
    wire \b2v_inst16.count_rst_2 ;
    wire \b2v_inst16.count_4_13 ;
    wire \b2v_inst16.countZ0Z_14 ;
    wire \b2v_inst16.count_rst_3 ;
    wire \b2v_inst16.count_4_14 ;
    wire \b2v_inst16.count_rst_7 ;
    wire \b2v_inst16.count_4_2 ;
    wire \b2v_inst16.count_rst_11 ;
    wire \b2v_inst16.count_4_6 ;
    wire \b2v_inst16.count_en ;
    wire \b2v_inst16.N_3037_i ;
    wire \b2v_inst36.curr_state_0_1 ;
    wire \b2v_inst36.curr_state_7_1_cascade_ ;
    wire \b2v_inst36.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst36.N_1_i ;
    wire \b2v_inst36.curr_state_0_0 ;
    wire \b2v_inst36.curr_state_7_0_cascade_ ;
    wire \b2v_inst36.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst36.count_0_sqmuxa ;
    wire \b2v_inst11.count_off_0_11 ;
    wire \b2v_inst11.count_off_0_10 ;
    wire \b2v_inst11.count_off_0_12 ;
    wire \b2v_inst11.count_off_0_3 ;
    wire \b2v_inst11.count_off_0_14 ;
    wire \b2v_inst11.count_offZ0Z_14_cascade_ ;
    wire \b2v_inst11.count_off_0_13 ;
    wire \b2v_inst11.g0_i_o3_0 ;
    wire \b2v_inst11.un85_clk_100khz1_THRU_CO ;
    wire \b2v_inst11.un85_clk_100khz0_THRU_CO ;
    wire \b2v_inst11.N_6_cascade_ ;
    wire \b2v_inst11.g0_0_0_rep1_1 ;
    wire \b2v_inst11.pwm_outZ0 ;
    wire \b2v_inst11.g0_i_a3_0_1 ;
    wire \b2v_inst11.N_6 ;
    wire pwrbtn_led;
    wire \b2v_inst200.count_enZ0 ;
    wire \b2v_inst16.delayed_vddq_pwrgd_en_cascade_ ;
    wire vpp_en;
    wire \b2v_inst16.curr_state_RNIBO6I1Z0Z_0 ;
    wire \b2v_inst16.N_268 ;
    wire \b2v_inst16.N_268_cascade_ ;
    wire \b2v_inst16.N_26 ;
    wire \b2v_inst11.countZ0Z_0 ;
    wire \b2v_inst11.count_0_sqmuxa_i ;
    wire \b2v_inst11.count_1_0 ;
    wire bfn_4_11_0_;
    wire \b2v_inst11.mult1_un166_sum_cry_0 ;
    wire \b2v_inst11.mult1_un166_sum_cry_1 ;
    wire \b2v_inst11.mult1_un166_sum_cry_2 ;
    wire \b2v_inst11.mult1_un166_sum_cry_3 ;
    wire G_2848;
    wire \b2v_inst11.mult1_un166_sum_cry_4 ;
    wire \b2v_inst11.mult1_un166_sum_cry_5 ;
    wire \b2v_inst11.mult1_un166_sum_s_6 ;
    wire bfn_4_12_0_;
    wire \b2v_inst11.mult1_un145_sum_cry_2 ;
    wire \b2v_inst11.mult1_un145_sum_cry_3 ;
    wire \b2v_inst11.mult1_un145_sum_cry_4 ;
    wire \b2v_inst11.mult1_un145_sum_cry_5 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6 ;
    wire \b2v_inst11.mult1_un145_sum_cry_7 ;
    wire \b2v_inst11.mult1_un138_sum_i_0_8 ;
    wire bfn_4_13_0_;
    wire \b2v_inst11.mult1_un138_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_2 ;
    wire \b2v_inst11.mult1_un138_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_3 ;
    wire \b2v_inst11.mult1_un138_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_4 ;
    wire \b2v_inst11.mult1_un138_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_5 ;
    wire \b2v_inst11.mult1_un145_sum_axb_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_6 ;
    wire \b2v_inst11.mult1_un138_sum_cry_7 ;
    wire \b2v_inst11.mult1_un138_sum_s_8 ;
    wire \b2v_inst11.mult1_un131_sum_i_0_8 ;
    wire bfn_4_14_0_;
    wire \b2v_inst11.mult1_un117_sum_cry_2 ;
    wire \b2v_inst11.mult1_un117_sum_cry_3 ;
    wire \b2v_inst11.mult1_un117_sum_cry_4 ;
    wire \b2v_inst11.mult1_un117_sum_cry_5 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6 ;
    wire \b2v_inst11.mult1_un117_sum_cry_7 ;
    wire \b2v_inst11.mult1_un117_sum_s_8_cascade_ ;
    wire bfn_4_15_0_;
    wire \b2v_inst11.mult1_un124_sum_cry_2 ;
    wire \b2v_inst11.mult1_un117_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_3 ;
    wire \b2v_inst11.mult1_un117_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_4 ;
    wire \b2v_inst11.mult1_un117_sum_s_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_5 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un117_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un124_sum_cry_6 ;
    wire \b2v_inst11.mult1_un124_sum_axb_8 ;
    wire \b2v_inst11.mult1_un124_sum_cry_7 ;
    wire \b2v_inst11.mult1_un117_sum_i ;
    wire bfn_4_16_0_;
    wire \b2v_inst11.mult1_un131_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_2 ;
    wire \b2v_inst11.mult1_un124_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_3 ;
    wire \b2v_inst11.mult1_un124_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_4 ;
    wire \b2v_inst11.mult1_un124_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_5 ;
    wire \b2v_inst11.mult1_un124_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un138_sum_axb_8 ;
    wire \b2v_inst11.mult1_un131_sum_cry_6 ;
    wire \b2v_inst11.mult1_un131_sum_axb_8 ;
    wire \b2v_inst11.mult1_un131_sum_cry_7 ;
    wire \b2v_inst11.mult1_un131_sum_s_8 ;
    wire \b2v_inst11.mult1_un124_sum_s_8 ;
    wire \b2v_inst11.mult1_un124_sum_i_0_8 ;
    wire \b2v_inst16.N_208_0 ;
    wire \b2v_inst16.delayed_vddq_pwrgd_en ;
    wire \b2v_inst16.curr_stateZ0Z_1 ;
    wire \b2v_inst16.delayed_vddq_pwrgdZ0 ;
    wire \b2v_inst200.count_1_0_cascade_ ;
    wire \b2v_inst200.un2_count_1_axb_1 ;
    wire bfn_5_2_0_;
    wire \b2v_inst200.countZ0Z_2 ;
    wire \b2v_inst200.un2_count_1_cry_1 ;
    wire \b2v_inst200.un2_count_1_axb_3 ;
    wire \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_2 ;
    wire \b2v_inst200.countZ0Z_4 ;
    wire \b2v_inst200.un2_count_1_cry_3 ;
    wire \b2v_inst200.un2_count_1_axb_5 ;
    wire \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_4 ;
    wire \b2v_inst200.un2_count_1_cry_5_cZ0 ;
    wire \b2v_inst200.countZ0Z_7 ;
    wire \b2v_inst200.un2_count_1_cry_6 ;
    wire \b2v_inst200.un2_count_1_cry_7 ;
    wire \b2v_inst200.un2_count_1_cry_8 ;
    wire \b2v_inst200.un2_count_1_axb_9 ;
    wire \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ;
    wire bfn_5_3_0_;
    wire \b2v_inst200.un2_count_1_cry_9 ;
    wire \b2v_inst200.countZ0Z_11 ;
    wire \b2v_inst200.un2_count_1_cry_10 ;
    wire \b2v_inst200.countZ0Z_12 ;
    wire \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ;
    wire \b2v_inst200.un2_count_1_cry_11 ;
    wire \b2v_inst200.un2_count_1_axb_13 ;
    wire \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ;
    wire \b2v_inst200.un2_count_1_cry_12 ;
    wire \b2v_inst200.countZ0Z_14 ;
    wire \b2v_inst200.un2_count_1_cry_13 ;
    wire \b2v_inst200.un2_count_1_cry_14 ;
    wire \b2v_inst200.un2_count_1_axb_16 ;
    wire \b2v_inst200.count_1_16 ;
    wire \b2v_inst200.un2_count_1_cry_15 ;
    wire \b2v_inst200.un2_count_1_cry_16 ;
    wire \b2v_inst200.countZ0Z_17 ;
    wire bfn_5_4_0_;
    wire \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ;
    wire \b2v_inst200.count_0_17 ;
    wire \b2v_inst200.N_56_cascade_ ;
    wire gpio_fpga_soc_1;
    wire \b2v_inst200.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst200.m6_i_0_cascade_ ;
    wire \b2v_inst200.N_58_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_0_cascade_ ;
    wire N_411;
    wire N_411_cascade_;
    wire \b2v_inst200.m6_i_0 ;
    wire \b2v_inst200.curr_state_3_0 ;
    wire bfn_5_6_0_;
    wire \b2v_inst11.un3_count_off_1_cry_1 ;
    wire \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ;
    wire \b2v_inst11.un3_count_off_1_cry_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_3 ;
    wire \b2v_inst11.un3_count_off_1_cry_4 ;
    wire \b2v_inst11.un3_count_off_1_cry_5 ;
    wire \b2v_inst11.un3_count_off_1_cry_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_7 ;
    wire \b2v_inst11.un3_count_off_1_cry_8 ;
    wire bfn_5_7_0_;
    wire \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ;
    wire \b2v_inst11.un3_count_off_1_cry_9 ;
    wire \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ;
    wire \b2v_inst11.un3_count_off_1_cry_10 ;
    wire \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ;
    wire \b2v_inst11.un3_count_off_1_cry_11 ;
    wire \b2v_inst11.count_offZ0Z_13 ;
    wire \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ;
    wire \b2v_inst11.un3_count_off_1_cry_12 ;
    wire \b2v_inst11.count_offZ0Z_14 ;
    wire \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ;
    wire \b2v_inst11.un3_count_off_1_cry_13 ;
    wire \b2v_inst11.count_offZ0Z_15 ;
    wire \b2v_inst11.un3_count_off_1_cry_14 ;
    wire \b2v_inst11.count_offZ0Z_12 ;
    wire \b2v_inst11.count_offZ0Z_11 ;
    wire \b2v_inst11.count_offZ0Z_10 ;
    wire \b2v_inst11.count_offZ0Z_9 ;
    wire \b2v_inst200.curr_state_i_2_cascade_ ;
    wire \b2v_inst200.i4_mux ;
    wire \b2v_inst200.N_2989_i ;
    wire \b2v_inst200.N_205_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_2 ;
    wire \b2v_inst200.HDA_SDO_ATP_0 ;
    wire \b2v_inst200.N_205 ;
    wire \b2v_inst200.curr_state_i_2 ;
    wire hda_sdo_atp;
    wire \b2v_inst200.N_282 ;
    wire \b2v_inst200.curr_stateZ0Z_1 ;
    wire \b2v_inst200.curr_stateZ0Z_0 ;
    wire \b2v_inst200.curr_state_3_1 ;
    wire bfn_5_9_0_;
    wire \b2v_inst20.counter_1_cry_1 ;
    wire \b2v_inst20.counter_1_cry_2 ;
    wire \b2v_inst20.counter_1_cry_3 ;
    wire \b2v_inst20.counter_1_cry_4 ;
    wire \b2v_inst20.counter_1_cry_5 ;
    wire \b2v_inst20.counter_1_cry_6 ;
    wire \b2v_inst20.counterZ0Z_8 ;
    wire \b2v_inst20.counter_1_cry_7 ;
    wire \b2v_inst20.counter_1_cry_8 ;
    wire \b2v_inst20.counterZ0Z_9 ;
    wire bfn_5_10_0_;
    wire \b2v_inst20.counterZ0Z_10 ;
    wire \b2v_inst20.counter_1_cry_9 ;
    wire \b2v_inst20.counterZ0Z_11 ;
    wire \b2v_inst20.counter_1_cry_10 ;
    wire \b2v_inst20.counter_1_cry_11 ;
    wire \b2v_inst20.counter_1_cry_12 ;
    wire \b2v_inst20.counter_1_cry_13 ;
    wire \b2v_inst20.counter_1_cry_14 ;
    wire \b2v_inst20.counter_1_cry_15 ;
    wire \b2v_inst20.counter_1_cry_16 ;
    wire bfn_5_11_0_;
    wire \b2v_inst20.counter_1_cry_17 ;
    wire \b2v_inst20.counter_1_cry_18 ;
    wire \b2v_inst20.counterZ0Z_20 ;
    wire \b2v_inst20.counter_1_cry_19 ;
    wire \b2v_inst20.counterZ0Z_21 ;
    wire \b2v_inst20.counter_1_cry_20 ;
    wire \b2v_inst20.counterZ0Z_22 ;
    wire \b2v_inst20.counter_1_cry_21 ;
    wire \b2v_inst20.counterZ0Z_23 ;
    wire \b2v_inst20.counter_1_cry_22 ;
    wire \b2v_inst20.counter_1_cry_23 ;
    wire \b2v_inst20.counter_1_cry_24 ;
    wire bfn_5_12_0_;
    wire \b2v_inst20.counter_1_cry_25 ;
    wire \b2v_inst20.counter_1_cry_26 ;
    wire \b2v_inst20.counterZ0Z_28 ;
    wire \b2v_inst20.counter_1_cry_27 ;
    wire \b2v_inst20.counterZ0Z_29 ;
    wire \b2v_inst20.counter_1_cry_28 ;
    wire \b2v_inst20.counterZ0Z_30 ;
    wire \b2v_inst20.counter_1_cry_29 ;
    wire \b2v_inst20.counter_1_cry_30 ;
    wire \b2v_inst20.counterZ0Z_31 ;
    wire \b2v_inst11.mult1_un138_sum_i ;
    wire \b2v_inst11.mult1_un124_sum_i ;
    wire \b2v_inst11.mult1_un110_sum_i ;
    wire bfn_5_14_0_;
    wire \b2v_inst11.mult1_un103_sum_i ;
    wire \b2v_inst11.mult1_un110_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_2 ;
    wire \b2v_inst11.mult1_un103_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_3 ;
    wire \b2v_inst11.mult1_un103_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_4 ;
    wire \b2v_inst11.mult1_un103_sum_s_8 ;
    wire \b2v_inst11.mult1_un103_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_5 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un103_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un117_sum_axb_8 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6 ;
    wire \b2v_inst11.mult1_un110_sum_axb_8 ;
    wire \b2v_inst11.mult1_un110_sum_cry_7 ;
    wire \b2v_inst11.mult1_un110_sum_s_8 ;
    wire \b2v_inst11.mult1_un110_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un110_sum_i_0_8 ;
    wire bfn_5_15_0_;
    wire \b2v_inst11.mult1_un89_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6 ;
    wire \b2v_inst11.mult1_un89_sum_cry_7 ;
    wire \b2v_inst11.mult1_un82_sum_i_0_8 ;
    wire bfn_5_16_0_;
    wire \b2v_inst11.mult1_un96_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un103_sum_axb_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_6 ;
    wire \b2v_inst11.mult1_un96_sum_axb_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_7 ;
    wire \b2v_inst11.mult1_un96_sum_s_8 ;
    wire \b2v_inst11.mult1_un89_sum_s_8 ;
    wire \b2v_inst11.mult1_un89_sum_i_0_8 ;
    wire \b2v_inst200.un2_count_1_axb_15 ;
    wire \b2v_inst200.un2_count_1_axb_8 ;
    wire \b2v_inst200.count_3_15 ;
    wire \b2v_inst200.countZ0Z_6 ;
    wire \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71 ;
    wire \b2v_inst200.count_1_8 ;
    wire \b2v_inst200.count_3_8 ;
    wire \b2v_inst200.countZ0Z_10 ;
    wire \b2v_inst200.un25_clk_100khz_14 ;
    wire \b2v_inst200.un25_clk_100khz_6 ;
    wire \b2v_inst200.un25_clk_100khz_7_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_13 ;
    wire \b2v_inst200.count_RNI5RUP8Z0Z_8 ;
    wire \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_ ;
    wire \b2v_inst200.countZ0Z_0 ;
    wire \b2v_inst200.count_3_0 ;
    wire \b2v_inst200.count_1_11 ;
    wire \b2v_inst200.count_3_11 ;
    wire \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ;
    wire \b2v_inst200.count_3_14 ;
    wire \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ;
    wire \b2v_inst200.count_3_2 ;
    wire \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ;
    wire \b2v_inst200.count_3_4 ;
    wire \b2v_inst200.count_1_6 ;
    wire \b2v_inst200.count_3_6 ;
    wire \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ;
    wire \b2v_inst200.count_3_7 ;
    wire \b2v_inst200.count_1_10 ;
    wire \b2v_inst200.count_3_10 ;
    wire \b2v_inst200.count_en_g ;
    wire bfn_6_3_0_;
    wire \b2v_inst5.un2_count_1_cry_0 ;
    wire \b2v_inst5.un2_count_1_cry_1 ;
    wire \b2v_inst5.un2_count_1_cry_2 ;
    wire \b2v_inst5.un2_count_1_cry_3 ;
    wire \b2v_inst5.un2_count_1_cry_4 ;
    wire \b2v_inst5.un2_count_1_cry_5 ;
    wire \b2v_inst5.un2_count_1_cry_6 ;
    wire \b2v_inst5.un2_count_1_cry_7 ;
    wire bfn_6_4_0_;
    wire \b2v_inst5.un2_count_1_cry_8 ;
    wire \b2v_inst5.un2_count_1_cry_9 ;
    wire \b2v_inst5.un2_count_1_cry_10 ;
    wire \b2v_inst5.un2_count_1_cry_11 ;
    wire \b2v_inst5.un2_count_1_cry_12 ;
    wire \b2v_inst5.un2_count_1_cry_13 ;
    wire \b2v_inst5.un2_count_1_cry_14 ;
    wire \b2v_inst5.countZ0Z_4_cascade_ ;
    wire \b2v_inst5.count_rst_6 ;
    wire \b2v_inst5.count_rst_6_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_8 ;
    wire \b2v_inst5.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst5.un2_count_1_axb_8_cascade_ ;
    wire \b2v_inst5.count_1_8 ;
    wire \b2v_inst5.count_rst_10 ;
    wire \b2v_inst5.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst5.countZ0Z_4 ;
    wire \b2v_inst5.count_1_4 ;
    wire \b2v_inst11.count_off_0_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ;
    wire \b2v_inst11.count_off_0_0 ;
    wire \b2v_inst11.count_offZ0Z_0 ;
    wire \b2v_inst11.count_offZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_off_RNIZ0Z_1 ;
    wire \b2v_inst11.count_off_0_1 ;
    wire \b2v_inst11.count_off_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_offZ0Z_1 ;
    wire \b2v_inst11.count_offZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_offZ0Z_2 ;
    wire \b2v_inst20.counterZ0Z_7 ;
    wire \b2v_inst20.counter_1_cry_4_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_5 ;
    wire \b2v_inst20.counter_1_cry_5_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_6 ;
    wire \b2v_inst11.count_offZ0Z_3 ;
    wire \b2v_inst20.counterZ0Z_1 ;
    wire v33dsw_ok;
    wire \b2v_inst36.curr_stateZ0Z_1 ;
    wire \b2v_inst36.curr_stateZ0Z_0 ;
    wire \b2v_inst11.count_offZ0Z_4 ;
    wire \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ;
    wire \b2v_inst11.count_off_0_4 ;
    wire \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ;
    wire \b2v_inst11.count_off_0_15 ;
    wire \b2v_inst11.count_off_0_5 ;
    wire \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ;
    wire \b2v_inst11.count_offZ0Z_5 ;
    wire \b2v_inst11.count_off_0_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ;
    wire \b2v_inst11.count_offZ0Z_6 ;
    wire bfn_6_9_0_;
    wire \b2v_inst20.un4_counter_1_and ;
    wire \b2v_inst20.un4_counter_0 ;
    wire \b2v_inst20.un4_counter_2_and ;
    wire \b2v_inst20.un4_counter_1 ;
    wire \b2v_inst20.un4_counter_2 ;
    wire \b2v_inst20.un4_counter_3 ;
    wire \b2v_inst20.un4_counter_5_and ;
    wire \b2v_inst20.un4_counter_4 ;
    wire \b2v_inst20.un4_counter_5 ;
    wire \b2v_inst20.un4_counter_7_and ;
    wire \b2v_inst20.un4_counter_6 ;
    wire b2v_inst20_un4_counter_7;
    wire bfn_6_10_0_;
    wire \b2v_inst20.counterZ0Z_16 ;
    wire \b2v_inst20.counterZ0Z_17 ;
    wire \b2v_inst20.counterZ0Z_18 ;
    wire \b2v_inst20.counterZ0Z_19 ;
    wire \b2v_inst20.un4_counter_4_and ;
    wire \b2v_inst20.counterZ0Z_15 ;
    wire \b2v_inst20.counterZ0Z_13 ;
    wire \b2v_inst20.counterZ0Z_14 ;
    wire \b2v_inst20.counterZ0Z_12 ;
    wire \b2v_inst20.un4_counter_3_and ;
    wire \b2v_inst20.counterZ0Z_24 ;
    wire \b2v_inst20.counterZ0Z_26 ;
    wire \b2v_inst20.counterZ0Z_25 ;
    wire \b2v_inst20.counterZ0Z_27 ;
    wire \b2v_inst20.un4_counter_6_and ;
    wire bfn_6_11_0_;
    wire \b2v_inst11.mult1_un159_sum_cry_2_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_1 ;
    wire \b2v_inst11.mult1_un159_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_2 ;
    wire \b2v_inst11.mult1_un159_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_3 ;
    wire \b2v_inst11.mult1_un159_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_4 ;
    wire \b2v_inst11.mult1_un166_sum_axb_6 ;
    wire \b2v_inst11.mult1_un159_sum_cry_5 ;
    wire \b2v_inst11.mult1_un159_sum_cry_6 ;
    wire \b2v_inst11.mult1_un159_sum_s_7 ;
    wire \b2v_inst11.mult1_un159_sum_i ;
    wire bfn_6_12_0_;
    wire \b2v_inst11.mult1_un145_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un152_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_2 ;
    wire \b2v_inst11.mult1_un145_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un152_sum_axb_4_l_fx ;
    wire \b2v_inst11.mult1_un152_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_3 ;
    wire \b2v_inst11.mult1_un145_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_4 ;
    wire \b2v_inst11.mult1_un145_sum_s_8 ;
    wire \b2v_inst11.mult1_un145_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_5 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un152_sum_axb_7_l_fx ;
    wire \b2v_inst11.mult1_un159_sum_axb_7 ;
    wire \b2v_inst11.mult1_un152_sum_cry_6 ;
    wire \b2v_inst11.mult1_un152_sum_axb_8 ;
    wire \b2v_inst11.mult1_un152_sum_cry_7 ;
    wire \b2v_inst11.mult1_un152_sum_s_8 ;
    wire \b2v_inst11.mult1_un152_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un152_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un82_sum_i ;
    wire \b2v_inst11.mult1_un96_sum_i ;
    wire pch_pwrok;
    wire bfn_6_14_0_;
    wire \b2v_inst11.mult1_un75_sum_i ;
    wire \b2v_inst11.mult1_un82_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_2 ;
    wire \b2v_inst11.mult1_un82_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_3 ;
    wire \b2v_inst11.mult1_un82_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_4 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_axb_8 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6 ;
    wire \b2v_inst11.mult1_un82_sum_cry_7 ;
    wire \b2v_inst11.mult1_un82_sum_s_8 ;
    wire \b2v_inst11.mult1_un75_sum_i_0_8 ;
    wire bfn_6_15_0_;
    wire \b2v_inst11.mult1_un68_sum_i ;
    wire \b2v_inst11.mult1_un75_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_2 ;
    wire \b2v_inst11.mult1_un75_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_3 ;
    wire \b2v_inst11.mult1_un75_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_4 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_5 ;
    wire \b2v_inst11.mult1_un82_sum_axb_8 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6 ;
    wire \b2v_inst11.mult1_un75_sum_cry_7 ;
    wire \b2v_inst11.mult1_un75_sum_s_8 ;
    wire \b2v_inst11.mult1_un68_sum_i_0_8 ;
    wire \b2v_inst5.un2_count_1_cry_4_c_RNIPKTZ0Z9 ;
    wire \b2v_inst5.count_1_5 ;
    wire \b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9 ;
    wire \b2v_inst5.count_1_6 ;
    wire \b2v_inst5.countZ0Z_13_cascade_ ;
    wire \b2v_inst5.count_1_13 ;
    wire \b2v_inst5.countZ0Z_3 ;
    wire \b2v_inst5.countZ0Z_3_cascade_ ;
    wire \b2v_inst5.countZ0Z_1 ;
    wire \b2v_inst5.un2_count_1_cry_0_c_RNILCPZ0Z9 ;
    wire \b2v_inst5.count_1_1 ;
    wire \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2 ;
    wire \b2v_inst5.count_1_12 ;
    wire \b2v_inst5.count_1_14 ;
    wire \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ;
    wire \b2v_inst5.countZ0Z_14 ;
    wire \b2v_inst5.countZ0Z_14_cascade_ ;
    wire \b2v_inst5.countZ0Z_12 ;
    wire \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_0 ;
    wire \b2v_inst5.curr_state_0_1 ;
    wire \b2v_inst5.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst5.count_1_0 ;
    wire \b2v_inst5.count_rst_14 ;
    wire \b2v_inst5.count_i_0 ;
    wire \b2v_inst5.curr_stateZ0Z_1 ;
    wire \b2v_inst5.count_1_15 ;
    wire \b2v_inst5.count_rst ;
    wire \b2v_inst5.countZ0Z_15 ;
    wire \b2v_inst5.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst5.N_51 ;
    wire \b2v_inst5.m4_0 ;
    wire curr_state_RNID8DP1_0_0_cascade_;
    wire N_413;
    wire \b2v_inst5.curr_state_0_0 ;
    wire \b2v_inst5.curr_stateZ0Z_0 ;
    wire \b2v_inst5.N_2856_i ;
    wire \b2v_inst5.curr_state_RNIZ0Z_1 ;
    wire \b2v_inst5.N_2856_i_cascade_ ;
    wire \b2v_inst11.count_off_0_7 ;
    wire \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ;
    wire \b2v_inst11.count_offZ0Z_7 ;
    wire \b2v_inst11.un34_clk_100khz_11 ;
    wire \b2v_inst11.un34_clk_100khz_9 ;
    wire \b2v_inst11.un34_clk_100khz_10 ;
    wire \b2v_inst11.un34_clk_100khz_8 ;
    wire \b2v_inst11.count_off_RNI_1Z0Z_1_cascade_ ;
    wire \b2v_inst11.func_state_1_m0_0_0_1_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ;
    wire \b2v_inst11.count_off_0_8 ;
    wire \b2v_inst11.count_offZ0Z_8 ;
    wire \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ;
    wire \b2v_inst11.count_off_0_9 ;
    wire \b2v_inst11.N_76_cascade_ ;
    wire \b2v_inst11.func_state_RNICMPB4Z0Z_0 ;
    wire \b2v_inst11.func_state_1_m2_1_cascade_ ;
    wire \b2v_inst11.func_state_cascade_ ;
    wire \b2v_inst11.N_339 ;
    wire \b2v_inst11.N_339_cascade_ ;
    wire \b2v_inst11.func_state_RNI6IFF4Z0Z_1 ;
    wire \b2v_inst36.DSW_PWROK_0 ;
    wire \b2v_inst36.curr_state_RNI3E27Z0Z_0 ;
    wire dsw_pwrok;
    wire \b2v_inst11.func_state_1_m2_1 ;
    wire \b2v_inst11.func_stateZ0Z_1 ;
    wire \b2v_inst11.un1_clk_100khz_51_and_i_a3_0_1_cascade_ ;
    wire vpp_ok;
    wire VCCST_EN_i_0_o3_0_cascade_;
    wire vddq_en;
    wire \b2v_inst11.count_clk_en_0_xZ0Z1_cascade_ ;
    wire \b2v_inst11.N_335 ;
    wire v5s_enn_cascade_;
    wire \b2v_inst20.counterZ0Z_0 ;
    wire \b2v_inst20.un4_counter_0_and ;
    wire \b2v_inst20.counter_1_cry_1_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_2 ;
    wire \b2v_inst20.counter_1_cry_2_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_3 ;
    wire \b2v_inst20.counter_1_cry_3_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_4 ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVKZ0_cascade_ ;
    wire \b2v_inst11.N_236 ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ;
    wire \b2v_inst11.N_295 ;
    wire \b2v_inst11.mult1_un152_sum_i ;
    wire \b2v_inst11.N_3055_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_14Z0Z_0 ;
    wire \b2v_inst11.un1_dutycycle_172_m3_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_172_0 ;
    wire \b2v_inst11.N_19_i_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_172_m0_ns_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_172_m0 ;
    wire \b2v_inst11.g0_4_1_cascade_ ;
    wire \b2v_inst11.N_293_0 ;
    wire \b2v_inst11.g0_3_2_0 ;
    wire \b2v_inst11.un2_count_clk_17_0_a2_1_4_cascade_ ;
    wire \b2v_inst11.N_363_cascade_ ;
    wire \b2v_inst11.mult1_un145_sum_i ;
    wire \b2v_inst11.mult1_un131_sum_i ;
    wire bfn_7_14_0_;
    wire \b2v_inst11.mult1_un54_sum_s_3_sf ;
    wire \b2v_inst11.mult1_un54_sum_cry_2 ;
    wire \b2v_inst11.mult1_un54_sum_cry_3 ;
    wire \b2v_inst11.mult1_un54_sum_cry_4 ;
    wire \b2v_inst11.mult1_un54_sum_cry_5 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6 ;
    wire \b2v_inst11.mult1_un54_sum_cry_7 ;
    wire bfn_7_15_0_;
    wire \b2v_inst11.mult1_un47_sum_i_1 ;
    wire \b2v_inst11.mult1_un61_sum_cry_2 ;
    wire \b2v_inst11.mult1_un54_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_7_THRU_CO ;
    wire \b2v_inst11.mult1_un61_sum_cry_3 ;
    wire \b2v_inst11.mult1_un54_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_4 ;
    wire \b2v_inst11.mult1_un54_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_5 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_6 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6_THRU_CO ;
    wire \b2v_inst11.mult1_un61_sum_cry_7 ;
    wire \b2v_inst11.mult1_un54_sum_s_8 ;
    wire \b2v_inst11.mult1_un54_sum_i_8 ;
    wire bfn_7_16_0_;
    wire \b2v_inst11.mult1_un68_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_2 ;
    wire \b2v_inst11.mult1_un61_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_3 ;
    wire \b2v_inst11.mult1_un61_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_4 ;
    wire \b2v_inst11.mult1_un61_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_5 ;
    wire \b2v_inst11.mult1_un61_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un75_sum_axb_8 ;
    wire \b2v_inst11.mult1_un68_sum_cry_6 ;
    wire \b2v_inst11.mult1_un68_sum_axb_8 ;
    wire \b2v_inst11.mult1_un68_sum_cry_7 ;
    wire \b2v_inst11.mult1_un68_sum_s_8 ;
    wire \b2v_inst11.mult1_un61_sum_s_8 ;
    wire \b2v_inst11.mult1_un61_sum_i_0_8 ;
    wire \b2v_inst6.count_rst_11_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_3_cascade_ ;
    wire \b2v_inst6.count_rst_10_cascade_ ;
    wire \b2v_inst6.count_rst_11 ;
    wire \b2v_inst6.count_0_3 ;
    wire \b2v_inst6.count_rst_10 ;
    wire \b2v_inst6.countZ0Z_3_cascade_ ;
    wire \b2v_inst6.count_0_4 ;
    wire \b2v_inst5.un2_count_1_axb_11 ;
    wire \b2v_inst5.count_1_7 ;
    wire \b2v_inst5.un2_count_1_cry_6_c_RNIROVZ0Z9 ;
    wire \b2v_inst5.countZ0Z_7 ;
    wire \b2v_inst5.count_rst_3 ;
    wire \b2v_inst5.count_1_11 ;
    wire \b2v_inst5.countZ0Z_7_cascade_ ;
    wire \b2v_inst5.un2_count_1_cry_1_c_RNIMEQZ0Z9 ;
    wire \b2v_inst5.count_1_2 ;
    wire \b2v_inst5.countZ0Z_2 ;
    wire \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ;
    wire \b2v_inst5.count_1_3 ;
    wire \b2v_inst5.un2_count_1_axb_10_cascade_ ;
    wire \b2v_inst5.un12_clk_100khz_9 ;
    wire \b2v_inst5.countZ0Z_5 ;
    wire \b2v_inst5.un12_clk_100khz_1 ;
    wire \b2v_inst5.countZ0Z_6 ;
    wire \b2v_inst5.un2_count_1_axb_10 ;
    wire \b2v_inst5.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst5.count_rst_4 ;
    wire \b2v_inst5.count_1_10 ;
    wire \b2v_inst5.count_rst_4_cascade_ ;
    wire \b2v_inst5.un12_clk_100khz_4 ;
    wire \b2v_inst5.un12_clk_100khz_11 ;
    wire \b2v_inst5.un12_clk_100khz_5_cascade_ ;
    wire \b2v_inst5.un12_clk_100khz_12 ;
    wire \b2v_inst5.N_1_i_cascade_ ;
    wire \b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ;
    wire \b2v_inst5.count_1_9 ;
    wire \b2v_inst5.countZ0Z_13 ;
    wire \b2v_inst5.un2_count_1_cry_12_THRU_CO ;
    wire \b2v_inst5.count_rst_1 ;
    wire \b2v_inst5.N_1_i ;
    wire \b2v_inst5.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst5.countZ0Z_9 ;
    wire \b2v_inst5.count_0_sqmuxa ;
    wire \b2v_inst5.count_rst_5 ;
    wire v33a_ok;
    wire vccst_cpu_ok;
    wire v1p8a_ok;
    wire v5a_ok;
    wire vr_ready_vccinaux;
    wire vr_ready_vccin;
    wire \b2v_inst6.N_192_cascade_ ;
    wire \b2v_inst6.N_241_cascade_ ;
    wire \b2v_inst11.count_clk_RNIG8KAHZ0Z_7_cascade_ ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_ ;
    wire \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1 ;
    wire \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1_cascade_ ;
    wire \b2v_inst11.N_428_cascade_ ;
    wire \b2v_inst11.count_clk_RNITV5AUZ0Z_7 ;
    wire \b2v_inst11.count_clk_RNILG61T1Z0Z_5 ;
    wire \b2v_inst11.un1_func_state25_4_i_a2_sxZ0_cascade_ ;
    wire rsmrstn_cascade_;
    wire \b2v_inst11.dutycycle_1_0_iv_i_0_2 ;
    wire b2v_inst20_un4_counter_7_THRU_CO;
    wire \b2v_inst11.func_state_1_ss0_i_0_o3_0 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_331_N ;
    wire \b2v_inst11.un1_func_state25_6_0_a3_0_1_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_332_N ;
    wire \b2v_inst11.func_state_RNI_2Z0Z_1 ;
    wire \b2v_inst11.N_337_cascade_ ;
    wire \b2v_inst11.func_state_1_m2s2_i_1 ;
    wire \b2v_inst11.N_76 ;
    wire \b2v_inst11.func_state_RNI6IFF4_0Z0Z_1 ;
    wire \b2v_inst11.func_state_1_m2_0_cascade_ ;
    wire \b2v_inst11.func_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.func_state_1_m2_0 ;
    wire VCCST_EN_i_0_o3_0;
    wire \b2v_inst11.func_stateZ1Z_0 ;
    wire \b2v_inst11.count_clk_en_0 ;
    wire \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_3_1 ;
    wire \b2v_inst11.d_N_5 ;
    wire \b2v_inst11.dutycycleZ1Z_5_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_5_cascade_ ;
    wire \b2v_inst11.N_293 ;
    wire \b2v_inst11.N_365 ;
    wire \b2v_inst11.N_159_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_9Z0Z_0 ;
    wire \b2v_inst11.un1_dutycycle_172_m3_d_ns_1_0_cascade_ ;
    wire \b2v_inst11.g1_1 ;
    wire \b2v_inst11.dutycycle_RNIDQ4A1Z0Z_5 ;
    wire \b2v_inst11.un1_dutycycle_172_m4_rn_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_11Z0Z_0 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_5 ;
    wire \b2v_inst11.un1_dutycycle_172_m4_rn_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_172_m4 ;
    wire \b2v_inst11.N_3057_0 ;
    wire \b2v_inst11.g1_0_0_0 ;
    wire \b2v_inst11.N_3055_0_0 ;
    wire \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_1_cascade_ ;
    wire \b2v_inst11.g0_0_1 ;
    wire \b2v_inst11.g1_0_1_0 ;
    wire \b2v_inst11.g0_3_2 ;
    wire \b2v_inst11.g2_1_0_1_cascade_ ;
    wire \b2v_inst11.g2_1_0 ;
    wire \b2v_inst11.dutycycle_RNI_10Z0Z_0 ;
    wire \b2v_inst11.dutycycle_RNIPKS23Z0Z_4_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08UZ0 ;
    wire \b2v_inst11.dutycycleZ1Z_4 ;
    wire \b2v_inst11.dutycycle_RNI5AV24Z0Z_4 ;
    wire \b2v_inst11.dutycycle_RNIPKS23Z0Z_4 ;
    wire \b2v_inst11.dutycycleZ0Z_6_cascade_ ;
    wire \b2v_inst11.un1_i3_mux_cascade_ ;
    wire \b2v_inst11.d_i3_mux ;
    wire \b2v_inst11.un1_dutycycle_53_axb_0 ;
    wire bfn_8_14_0_;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_0 ;
    wire \b2v_inst11.mult1_un138_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_0 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_2 ;
    wire \b2v_inst11.mult1_un131_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_2 ;
    wire \b2v_inst11.mult1_un124_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_2 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_5 ;
    wire \b2v_inst11.mult1_un117_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_3 ;
    wire \b2v_inst11.mult1_un110_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_4 ;
    wire \b2v_inst11.mult1_un103_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_5 ;
    wire \b2v_inst11.mult1_un96_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_6 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_7 ;
    wire bfn_8_15_0_;
    wire \b2v_inst11.mult1_un82_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_8 ;
    wire \b2v_inst11.mult1_un75_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_9 ;
    wire \b2v_inst11.mult1_un68_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_10 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_11 ;
    wire \b2v_inst11.mult1_un47_sum_1 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_12 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15 ;
    wire bfn_8_16_0_;
    wire \b2v_inst11.CO2 ;
    wire \b2v_inst11.mult1_un61_sum ;
    wire \b2v_inst11.mult1_un61_sum_i ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_13 ;
    wire \b2v_inst11.mult1_un47_sum_6 ;
    wire \b2v_inst11.mult1_un89_sum ;
    wire \b2v_inst11.mult1_un89_sum_i ;
    wire \b2v_inst6.un2_count_1_axb_8_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_9_cascade_ ;
    wire \b2v_inst6.count_rst_6 ;
    wire \b2v_inst6.count_rst_5 ;
    wire \b2v_inst6.countZ0Z_8_cascade_ ;
    wire \b2v_inst6.count_0_9 ;
    wire \b2v_inst6.count_0_8 ;
    wire N_607_g;
    wire \b2v_inst6.N_394_cascade_ ;
    wire \b2v_inst6.curr_state_1_1 ;
    wire \b2v_inst6.m6_i_a3_cascade_ ;
    wire \b2v_inst6.curr_stateZ0Z_1 ;
    wire \b2v_inst6.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst6.curr_state_1_0 ;
    wire \b2v_inst6.curr_state_7_0_cascade_ ;
    wire \b2v_inst6.count_RNICV5H1Z0Z_0_cascade_ ;
    wire \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ;
    wire N_222;
    wire \b2v_inst6.N_2992_i_cascade_ ;
    wire SYNTHESIZED_WIRE_8;
    wire v5s_ok;
    wire v33s_ok;
    wire vccinaux_en;
    wire \b2v_inst6.curr_stateZ0Z_0 ;
    wire \b2v_inst6.curr_state_RNIKIRD1Z0Z_0 ;
    wire \b2v_inst6.N_276_0 ;
    wire \b2v_inst6.curr_state_RNIKIRD1Z0Z_0_cascade_ ;
    wire \b2v_inst6.delayed_vccin_vccinaux_ok_0 ;
    wire \b2v_inst6.N_2992_i ;
    wire \b2v_inst6.N_3011_i ;
    wire \b2v_inst6.N_192 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_clk_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst11.un1_count_clk_2_axb_1_cascade_ ;
    wire \b2v_inst11.count_clk_0_0 ;
    wire \b2v_inst11.count_clk_0_1 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_1 ;
    wire \b2v_inst11.count_clkZ0Z_1 ;
    wire \b2v_inst11.N_379 ;
    wire \b2v_inst11.count_clkZ0Z_3_cascade_ ;
    wire \b2v_inst11.N_190 ;
    wire \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_3 ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5Z0Z_0_cascade_ ;
    wire \b2v_inst11.count_clk_0_3 ;
    wire \b2v_inst11.N_428 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_ ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ;
    wire \b2v_inst11.func_state_1_m2_am_1_0_cascade_ ;
    wire \b2v_inst11.func_state_RNINCPR4Z0Z_0 ;
    wire \b2v_inst11.N_382 ;
    wire \b2v_inst11.N_315 ;
    wire vccst_en;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0 ;
    wire \b2v_inst11.count_clk_RNIG510TZ0Z_5 ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_1 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_ ;
    wire \b2v_inst11.count_off_enZ0 ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_ ;
    wire SYNTHESIZED_WIRE_1keep_3;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6_cascade_ ;
    wire \b2v_inst11.N_382_N ;
    wire SYNTHESIZED_WIRE_1keep_3_fast;
    wire RSMRSTn_0;
    wire \b2v_inst11.g0_4_sx_cascade_ ;
    wire curr_state_RNID8DP1_0_0;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0_0 ;
    wire \b2v_inst11.N_160_i ;
    wire \b2v_inst11.N_160_i_cascade_ ;
    wire \b2v_inst11.func_state_RNI5DLRZ0Z_0 ;
    wire \b2v_inst11.N_366 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_0 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_313_N ;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2BZ0_cascade_ ;
    wire \b2v_inst11.dutycycle_1_0_1 ;
    wire \b2v_inst11.dutycycle_1_0_1_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_1 ;
    wire \b2v_inst11.dutycycle_1_0_0 ;
    wire \b2v_inst11.dutycycleZ1Z_0 ;
    wire \b2v_inst11.dutycycle_1_0_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_8Z0Z_0 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_2 ;
    wire \b2v_inst11.N_19_i ;
    wire \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_0_cascade_ ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1 ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \b2v_inst11.N_186_i_cascade_ ;
    wire \b2v_inst11.N_309 ;
    wire \b2v_inst11.un1_dutycycle_96_0_a3_1 ;
    wire \b2v_inst11.dutycycle_eena_0 ;
    wire \b2v_inst11.un1_clk_100khz_25_and_i_0_1_0 ;
    wire \b2v_inst11.N_186_i ;
    wire \b2v_inst11.N_117_f0_1 ;
    wire v5s_enn;
    wire \b2v_inst11.N_117_f0_1_cascade_ ;
    wire \b2v_inst11.dutycycle_eena ;
    wire \b2v_inst11.dutycycleZ1Z_2 ;
    wire \b2v_inst11.N_73 ;
    wire \b2v_inst11.dutycycle_eena_1 ;
    wire \b2v_inst11.N_159 ;
    wire \b2v_inst11.dutycycleZ0Z_1_cascade_ ;
    wire \b2v_inst11.N_363 ;
    wire \b2v_inst11.func_state_RNI_1Z0Z_1 ;
    wire \b2v_inst11.dutycycle_eena_9_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_7_cascade_ ;
    wire \b2v_inst11.N_2943_i ;
    wire \b2v_inst11.func_state_RNIDQ4A1Z0Z_1 ;
    wire \b2v_inst11.N_360_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ;
    wire \b2v_inst11.N_234_N ;
    wire \b2v_inst11.dutycycle_eena_9 ;
    wire \b2v_inst11.dutycycleZ1Z_12 ;
    wire \b2v_inst11.dutycycleZ1Z_11 ;
    wire \b2v_inst11.dutycycle_eena_7 ;
    wire \b2v_inst11.N_6_0 ;
    wire \b2v_inst11.N_8_cascade_ ;
    wire \b2v_inst11.N_355 ;
    wire \b2v_inst11.g0_6_a5_0_0_cascade_ ;
    wire \b2v_inst11.g0_6_a5_2_1 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_7 ;
    wire \b2v_inst11.CO2_THRU_CO ;
    wire \b2v_inst11.mult1_un54_sum_axb_6_i_l_fx ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ;
    wire \b2v_inst11.mult1_un54_sum_axb_5_i_l_ofx ;
    wire \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0 ;
    wire \b2v_inst11.mult1_un40_sum_i_2 ;
    wire \b2v_inst11.mult1_un47_sum1_3 ;
    wire \b2v_inst11.un1_dutycycle_53_axb_12_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_15 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_6 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_11 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_15 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_14 ;
    wire \b2v_inst11.un1_dutycycle_53_44_0_0 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_7 ;
    wire \b2v_inst11.un1_dutycycle_53_axb_10 ;
    wire \b2v_inst11.N_11_cascade_ ;
    wire \b2v_inst11.N_35_0 ;
    wire \b2v_inst11.N_13_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_11 ;
    wire \b2v_inst11.g0_6_a5_1_0 ;
    wire \b2v_inst6.count_rst_7_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_7_cascade_ ;
    wire \b2v_inst6.count_rst_3_cascade_ ;
    wire \b2v_inst6.countZ0Z_11_cascade_ ;
    wire \b2v_inst6.count_0_11 ;
    wire \b2v_inst6.N_394 ;
    wire bfn_11_2_0_;
    wire \b2v_inst6.un2_count_1_cry_1 ;
    wire \b2v_inst6.un2_count_1_axb_3 ;
    wire \b2v_inst6.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_2 ;
    wire \b2v_inst6.un2_count_1_axb_4 ;
    wire \b2v_inst6.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_3 ;
    wire \b2v_inst6.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_4 ;
    wire \b2v_inst6.un2_count_1_cry_5 ;
    wire \b2v_inst6.un2_count_1_axb_7 ;
    wire \b2v_inst6.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_6 ;
    wire \b2v_inst6.un2_count_1_axb_8 ;
    wire \b2v_inst6.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_7 ;
    wire \b2v_inst6.un2_count_1_cry_8 ;
    wire \b2v_inst6.un2_count_1_axb_9 ;
    wire \b2v_inst6.un2_count_1_cry_8_THRU_CO ;
    wire bfn_11_3_0_;
    wire \b2v_inst6.un2_count_1_cry_9 ;
    wire \b2v_inst6.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_10 ;
    wire \b2v_inst6.un2_count_1_cry_11 ;
    wire \b2v_inst6.un2_count_1_cry_12 ;
    wire \b2v_inst6.un2_count_1_cry_13 ;
    wire \b2v_inst6.un2_count_1_cry_14 ;
    wire \b2v_inst6.un2_count_1_axb_13 ;
    wire \b2v_inst11.count_clkZ0Z_10 ;
    wire \b2v_inst11.count_clkZ0Z_12 ;
    wire \b2v_inst11.count_clkZ0Z_13_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_11 ;
    wire \b2v_inst11.un2_count_clk_17_0_o2_4_cascade_ ;
    wire \b2v_inst11.N_175 ;
    wire \b2v_inst11.count_clk_0_10 ;
    wire \b2v_inst11.un1_count_clk_2_axb_1 ;
    wire \b2v_inst11.count_clkZ0Z_0 ;
    wire bfn_11_5_0_;
    wire \b2v_inst11.un1_count_clk_2_cry_1 ;
    wire \b2v_inst11.un1_count_clk_2_axb_3 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_cZ0 ;
    wire bfn_11_6_0_;
    wire \b2v_inst11.un1_count_clk_2_axb_10 ;
    wire \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_9_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_axb_11 ;
    wire \b2v_inst11.un1_count_clk_2_cry_10_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_11 ;
    wire \b2v_inst11.un1_count_clk_2_cry_12 ;
    wire \b2v_inst11.un1_count_clk_2_cry_13 ;
    wire \b2v_inst11.func_state_RNIIGCET1_0_1 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14 ;
    wire \b2v_inst11.count_clk_1_11 ;
    wire \b2v_inst11.count_clk_0_11 ;
    wire \b2v_inst11.count_clkZ0Z_7 ;
    wire \b2v_inst11.count_clkZ0Z_8 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ;
    wire \b2v_inst11.count_clk_0_8 ;
    wire \b2v_inst11.count_clkZ0Z_9 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ;
    wire \b2v_inst11.count_clk_0_9 ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ;
    wire \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0_cascade_ ;
    wire \b2v_inst11.N_369 ;
    wire \b2v_inst11.count_clk_en_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_14 ;
    wire \b2v_inst11.N_417 ;
    wire \b2v_inst11.func_state_RNID7Q51Z0Z_0 ;
    wire \b2v_inst11.count_off_RNI_1Z0Z_1 ;
    wire \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0 ;
    wire \b2v_inst11.func_state_RNI6M5R2Z0Z_1 ;
    wire \b2v_inst11.func_state_RNIJGA54Z0Z_1 ;
    wire \b2v_inst11.count_clk_1_14 ;
    wire \b2v_inst11.count_clk_0_14 ;
    wire \b2v_inst11.func_stateZ0Z_0 ;
    wire \b2v_inst11.N_2904_i_cascade_ ;
    wire bfn_11_9_0_;
    wire \b2v_inst11.dutycycle_RNIZ0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_s1 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_2 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_2 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_s1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2_s1 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_4 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3_s1 ;
    wire CONSTANT_ONE_NET;
    wire \b2v_inst11.un1_dutycycle_94_cry_4_s1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_s1 ;
    wire \b2v_inst11.dutycycle_RNI_9Z0Z_7 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_s1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_s1 ;
    wire bfn_11_10_0_;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_s1 ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_10 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_s1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10_s1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11_s1 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_s1 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_14 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_s1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14_s1 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_6 ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_3 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_3 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EGZ0Z1 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_11 ;
    wire \b2v_inst11.dutycycle_rst_6 ;
    wire \b2v_inst11.dutycycle ;
    wire bfn_11_13_0_;
    wire \b2v_inst11.dutycycleZ0Z_2 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_s0 ;
    wire \b2v_inst11.dutycycleZ0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_2 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_2 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_s0 ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_3 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2_s0 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_4 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3_s0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_4_s0 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_6 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_s0 ;
    wire \b2v_inst11.dutycycle_RNI_10Z0Z_7 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_s0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_s0 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_8 ;
    wire bfn_11_14_0_;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_s0 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_10 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_s0 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_11 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10_s0 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_12 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11_s0 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_s0 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_14 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_s0 ;
    wire \b2v_inst11.un1_dutycycle_94_axb_15_s0 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_15 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14_s0 ;
    wire \b2v_inst11.un1_dutycycle_53_axb_12_1 ;
    wire \b2v_inst11.un1_dutycycle_53_3_1 ;
    wire \b2v_inst11.un1_dutycycle_53_31_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_53_31 ;
    wire \b2v_inst11.un1_dutycycle_53_55_0_tz ;
    wire \b2v_inst11.un1_dutycycle_53_axb_14_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_14_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_14 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_9 ;
    wire \b2v_inst11.N_2904_i ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_12 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_7 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_9_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_10 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_9 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_9 ;
    wire \b2v_inst11.i2_mux_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_5 ;
    wire \b2v_inst11.un1_N_5_cascade_ ;
    wire \b2v_inst11.un1_i2_mux_0_0 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_11 ;
    wire \b2v_inst6.count_rst_7 ;
    wire \b2v_inst6.count_0_7 ;
    wire \b2v_inst6.countZ0Z_5_cascade_ ;
    wire \b2v_inst6.count_RNICV5H1Z0Z_1_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_1 ;
    wire \b2v_inst6.un2_count_1_axb_1_cascade_ ;
    wire \b2v_inst6.count_RNICV5H1Z0Z_1 ;
    wire \b2v_inst6.countZ0Z_11 ;
    wire \b2v_inst6.count_0_1 ;
    wire \b2v_inst6.count_1_i_a3_4_0 ;
    wire \b2v_inst6.count_1_i_a3_6_0 ;
    wire \b2v_inst6.count_1_i_a3_3_0_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_5_0 ;
    wire \b2v_inst6.count_0_5 ;
    wire \b2v_inst6.count_rst_9 ;
    wire \b2v_inst6.un2_count_1_axb_5 ;
    wire \b2v_inst6.count_0_14 ;
    wire \b2v_inst6.un2_count_1_cry_13_c_RNIR6IOZ0Z5 ;
    wire \b2v_inst6.un2_count_1_axb_14 ;
    wire \b2v_inst6.countZ0Z_14 ;
    wire \b2v_inst6.count_rst_12_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_12_0 ;
    wire \b2v_inst6.count_1_i_a3_1_0_cascade_ ;
    wire \b2v_inst6.count_0_2 ;
    wire \b2v_inst6.un2_count_1_cry_1_c_RNIN2PZ0Z3 ;
    wire \b2v_inst6.un2_count_1_axb_2 ;
    wire \b2v_inst6.countZ0Z_6_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_0_0_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_7_0 ;
    wire \b2v_inst6.count_0_6 ;
    wire \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ;
    wire \b2v_inst6.un2_count_1_axb_6 ;
    wire \b2v_inst6.count_rst_2 ;
    wire \b2v_inst6.count_0_12 ;
    wire \b2v_inst6.un2_count_1_cry_11_c_RNI8RABZ0 ;
    wire \b2v_inst6.un2_count_1_axb_12 ;
    wire \b2v_inst6.un2_count_1_axb_10 ;
    wire \b2v_inst6.count_0_10 ;
    wire \b2v_inst6.un2_count_1_cry_9_c_RNIVIZ0Z14 ;
    wire \b2v_inst6.count_rst_4 ;
    wire \b2v_inst6.countZ0Z_15 ;
    wire \b2v_inst6.count_0_13 ;
    wire \b2v_inst6.countZ0Z_15_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_2_0 ;
    wire \b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0 ;
    wire \b2v_inst6.count_rst_1 ;
    wire \b2v_inst11.un1_count_clk_2_axb_12 ;
    wire \b2v_inst11.count_clk_1_12 ;
    wire \b2v_inst11.count_clk_0_12 ;
    wire \b2v_inst11.un1_count_clk_2_axb_13 ;
    wire \b2v_inst11.count_clk_1_13 ;
    wire \b2v_inst11.count_clk_0_13 ;
    wire \b2v_inst11.un1_count_clk_2_axb_5 ;
    wire \b2v_inst11.count_clk_0_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ;
    wire \b2v_inst11.count_clkZ0Z_5 ;
    wire \b2v_inst11.count_clk_0_7 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_axb_7 ;
    wire \b2v_inst11.count_clkZ0Z_4 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ;
    wire \b2v_inst11.count_clk_0_4 ;
    wire \b2v_inst11.un1_count_clk_2_axb_2 ;
    wire \b2v_inst11.count_clk_0_2 ;
    wire \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ;
    wire \b2v_inst11.count_clkZ0Z_2 ;
    wire \b2v_inst11.count_clkZ0Z_15 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ;
    wire \b2v_inst11.count_clk_0_15 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ;
    wire \b2v_inst11.count_clk_0_6 ;
    wire \b2v_inst11.count_clk_en ;
    wire \b2v_inst11.count_clkZ0Z_6 ;
    wire \b2v_inst6.N_241 ;
    wire \b2v_inst6.countZ0Z_0 ;
    wire \b2v_inst6.N_2994_i ;
    wire \b2v_inst6.N_2994_i_cascade_ ;
    wire \b2v_inst6.N_389 ;
    wire \b2v_inst6.count_0_0 ;
    wire \b2v_inst6.count_rst ;
    wire \b2v_inst6.count_0_15 ;
    wire \b2v_inst6.count_en ;
    wire \b2v_inst6.curr_state_RNICV5H1Z0Z_0 ;
    wire \b2v_inst11.func_state_RNI_4Z0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_s0_sf ;
    wire \b2v_inst11.count_clk_RNIG510TZ0Z_7 ;
    wire \b2v_inst11.N_305 ;
    wire \b2v_inst11.N_306 ;
    wire \b2v_inst11.N_231_N_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_13_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4 ;
    wire \b2v_inst11.dutycycle_0_6 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_13 ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ;
    wire \b2v_inst11.dutycycleZ1Z_6_cascade_ ;
    wire \b2v_inst11.dutycycle_RNILF063Z0Z_6 ;
    wire \b2v_inst11.N_172 ;
    wire \b2v_inst11.N_185 ;
    wire \b2v_inst11.dutycycle_set_1 ;
    wire \b2v_inst11.dutycycle_set_1_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_14_0 ;
    wire \b2v_inst11.dutycycle_0_5 ;
    wire \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJZ0Z9 ;
    wire \b2v_inst11.dutycycle_RNIM98E2Z0Z_3 ;
    wire \b2v_inst11.dutycycleZ1Z_3 ;
    wire \b2v_inst11.dutycycle_RNIM98E2Z0Z_3_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3 ;
    wire \b2v_inst11.dutycycleZ0Z_9 ;
    wire SYNTHESIZED_WIRE_1keep_3_rep1;
    wire \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_32_and_i_0_c_0_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_32_and_i_0_d ;
    wire \b2v_inst11.un1_clk_100khz_33_and_i_0_c_0_cascade_ ;
    wire \b2v_inst11.N_153_N ;
    wire \b2v_inst11.N_155_N_cascade_ ;
    wire \b2v_inst11.g0_0_1_0_cascade_ ;
    wire \b2v_inst11.g0_1_1 ;
    wire \b2v_inst11.g3_0_0 ;
    wire rsmrstn;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_7_cascade_ ;
    wire \b2v_inst11.g1_0_0 ;
    wire \b2v_inst11.un1_clk_100khz_36_and_i_0_0 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_7 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_7 ;
    wire \b2v_inst11.un1_dutycycle_94_0_7 ;
    wire \b2v_inst11.g0_0_1_0 ;
    wire \b2v_inst11.dutycycleZ1Z_7 ;
    wire \b2v_inst11.un1_dutycycle_94_0_7_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_s1_13 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_13 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0 ;
    wire \b2v_inst11.dutycycleZ0Z_13 ;
    wire \b2v_inst11.dutycycle_en_10 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_12 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_5 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_5 ;
    wire \b2v_inst11.N_302 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_6 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_6 ;
    wire \b2v_inst11.N_301 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_14 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_14 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0 ;
    wire \b2v_inst11.dutycycle_en_11 ;
    wire \b2v_inst11.dutycycleZ0Z_14 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_10 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_6 ;
    wire \b2v_inst11.un1_dutycycle_53_44_0_3_tz_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_44_1 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_10 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_10 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642 ;
    wire \b2v_inst11.dutycycleZ1Z_10 ;
    wire \b2v_inst11.dutycycle_eena_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_7 ;
    wire \b2v_inst11.dutycycleZ0Z_3_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_44_0_1 ;
    wire \b2v_inst11.dutycycleZ0Z_3 ;
    wire \b2v_inst11.g1_i_0 ;
    wire \b2v_inst11.dutycycle_eena_2 ;
    wire \b2v_inst11.dutycycleZ1Z_9 ;
    wire \b2v_inst11.dutycycle_eena_2_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1 ;
    wire \b2v_inst11.dutycycleZ0Z_0_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_30_and_i_0_0_1 ;
    wire \b2v_inst11.dutycycleZ0Z_10 ;
    wire \b2v_inst11.N_140_N ;
    wire \b2v_inst11.N_425 ;
    wire \b2v_inst11.N_158_N_cascade_ ;
    wire \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ;
    wire \b2v_inst11.dutycycle_en_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3AZ0Z64 ;
    wire \b2v_inst11.dutycycle_en_12_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_15 ;
    wire \b2v_inst11.N_326_N ;
    wire fpga_osc;
    wire \b2v_inst11.N_224_iZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_s1_8 ;
    wire \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_94_s0_8 ;
    wire \b2v_inst11.dutycycleZ1Z_5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1 ;
    wire \b2v_inst11.dutycycleZ1Z_8 ;
    wire \b2v_inst11.dutycycle_eena_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1_cascade_ ;
    wire G_149;
    wire \b2v_inst11.dutycycleZ0Z_4_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_6 ;
    wire \b2v_inst11.dutycycleZ0Z_0 ;
    wire \b2v_inst11.dutycycleZ0Z_7 ;
    wire \b2v_inst11.dutycycleZ0Z_4 ;
    wire \b2v_inst11.un1_i2_mux_0 ;
    wire \b2v_inst11.un1_N_5 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_12 ;
    wire \b2v_inst11.dutycycleZ0Z_8 ;
    wire \b2v_inst11.un1_dutycycle_53_s_9_sf_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_12 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_1 ;
    wire \b2v_inst11.N_371_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_cascade_ ;
    wire \b2v_inst11.func_state_RNIDUQ02Z0Z_1 ;
    wire \b2v_inst11.g2_0_0Z0Z_0 ;
    wire gpio_fpga_soc_4;
    wire \b2v_inst11.func_state ;
    wire \b2v_inst11.g2_3Z0Z_0_cascade_ ;
    wire \b2v_inst11.N_200_i ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_0 ;
    wire slp_s3n;
    wire slp_s4n;
    wire \b2v_inst11.N_161 ;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__39838),
            .DIN(N__39837),
            .DOUT(N__39836),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__39838),
            .PADOUT(N__39837),
            .PADIN(N__39836),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccinaux),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__39829),
            .DIN(N__39828),
            .DOUT(N__39827),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__39829),
            .PADOUT(N__39828),
            .PADIN(N__39827),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__39820),
            .DIN(N__39819),
            .DOUT(N__39818),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__39820),
            .PADOUT(N__39819),
            .PADIN(N__39818),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__39811),
            .DIN(N__39810),
            .DOUT(N__39809),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__39811),
            .PADOUT(N__39810),
            .PADIN(N__39809),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24846),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__39802),
            .DIN(N__39801),
            .DOUT(N__39800),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__39802),
            .PADOUT(N__39801),
            .PADIN(N__39800),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__39793),
            .DIN(N__39792),
            .DOUT(N__39791),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__39793),
            .PADOUT(N__39792),
            .PADIN(N__39791),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__39784),
            .DIN(N__39783),
            .DOUT(N__39782),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__39784),
            .PADOUT(N__39783),
            .PADIN(N__39782),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__39775),
            .DIN(N__39774),
            .DOUT(N__39773),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__39775),
            .PADOUT(N__39774),
            .PADIN(N__39773),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__39766),
            .DIN(N__39765),
            .DOUT(N__39764),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__39766),
            .PADOUT(N__39765),
            .PADIN(N__39764),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29116),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__39757),
            .DIN(N__39756),
            .DOUT(N__39755),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__39757),
            .PADOUT(N__39756),
            .PADIN(N__39755),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__39748),
            .DIN(N__39747),
            .DOUT(N__39746),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__39748),
            .PADOUT(N__39747),
            .PADIN(N__39746),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__39739),
            .DIN(N__39738),
            .DOUT(N__39737),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__39739),
            .PADOUT(N__39738),
            .PADIN(N__39737),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19878),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__39730),
            .DIN(N__39729),
            .DOUT(N__39728),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__39730),
            .PADOUT(N__39729),
            .PADIN(N__39728),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__39721),
            .DIN(N__39720),
            .DOUT(N__39719),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__39721),
            .PADOUT(N__39720),
            .PADIN(N__39719),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__39712),
            .DIN(N__39711),
            .DOUT(N__39710),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__39712),
            .PADOUT(N__39711),
            .PADIN(N__39710),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__39703),
            .DIN(N__39702),
            .DOUT(N__39701),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__39703),
            .PADOUT(N__39702),
            .PADIN(N__39701),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__39694),
            .DIN(N__39693),
            .DOUT(N__39692),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__39694),
            .PADOUT(N__39693),
            .PADIN(N__39692),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27984),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__39685),
            .DIN(N__39684),
            .DOUT(N__39683),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__39685),
            .PADOUT(N__39684),
            .PADIN(N__39683),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__39676),
            .DIN(N__39675),
            .DOUT(N__39674),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__39676),
            .PADOUT(N__39675),
            .PADIN(N__39674),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__39667),
            .DIN(N__39666),
            .DOUT(N__39665),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__39667),
            .PADOUT(N__39666),
            .PADIN(N__39665),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__39658),
            .DIN(N__39657),
            .DOUT(N__39656),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__39658),
            .PADOUT(N__39657),
            .PADIN(N__39656),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__39649),
            .DIN(N__39648),
            .DOUT(N__39647),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__39649),
            .PADOUT(N__39648),
            .PADIN(N__39647),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    defparam ipInertedIOPad_VR_READY_VCCIN_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__39640),
            .DIN(N__39639),
            .DOUT(N__39638),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__39640),
            .PADOUT(N__39639),
            .PADIN(N__39638),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__39631),
            .DIN(N__39630),
            .DOUT(N__39629),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__39631),
            .PADOUT(N__39630),
            .PADIN(N__39629),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__39622),
            .DIN(N__39621),
            .DOUT(N__39620),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__39622),
            .PADOUT(N__39621),
            .PADIN(N__39620),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34842),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__39613),
            .DIN(N__39612),
            .DOUT(N__39611),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__39613),
            .PADOUT(N__39612),
            .PADIN(N__39611),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__39604),
            .DIN(N__39603),
            .DOUT(N__39602),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__39604),
            .PADOUT(N__39603),
            .PADIN(N__39602),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23941),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__39595),
            .DIN(N__39594),
            .DOUT(N__39593),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__39595),
            .PADOUT(N__39594),
            .PADIN(N__39593),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23945),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__39586),
            .DIN(N__39585),
            .DOUT(N__39584),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__39586),
            .PADOUT(N__39585),
            .PADIN(N__39584),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__39577),
            .DIN(N__39576),
            .DOUT(N__39575),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__39577),
            .PADOUT(N__39576),
            .PADIN(N__39575),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__39568),
            .DIN(N__39567),
            .DOUT(N__39566),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__39568),
            .PADOUT(N__39567),
            .PADIN(N__39566),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__39559),
            .DIN(N__39558),
            .DOUT(N__39557),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__39559),
            .PADOUT(N__39558),
            .PADIN(N__39557),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__39550),
            .DIN(N__39549),
            .DOUT(N__39548),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__39550),
            .PADOUT(N__39549),
            .PADIN(N__39548),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__39541),
            .DIN(N__39540),
            .DOUT(N__39539),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__39541),
            .PADOUT(N__39540),
            .PADIN(N__39539),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21369),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__39532),
            .DIN(N__39531),
            .DOUT(N__39530),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__39532),
            .PADOUT(N__39531),
            .PADIN(N__39530),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__39523),
            .DIN(N__39522),
            .DOUT(N__39521),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__39523),
            .PADOUT(N__39522),
            .PADIN(N__39521),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19848),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__39514),
            .DIN(N__39513),
            .DOUT(N__39512),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__39514),
            .PADOUT(N__39513),
            .PADIN(N__39512),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__39505),
            .DIN(N__39504),
            .DOUT(N__39503),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__39505),
            .PADOUT(N__39504),
            .PADIN(N__39503),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__39496),
            .DIN(N__39495),
            .DOUT(N__39494),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__39496),
            .PADOUT(N__39495),
            .PADIN(N__39494),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__39487),
            .DIN(N__39486),
            .DOUT(N__39485),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__39487),
            .PADOUT(N__39486),
            .PADIN(N__39485),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__39478),
            .DIN(N__39477),
            .DOUT(N__39476),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__39478),
            .PADOUT(N__39477),
            .PADIN(N__39476),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27668),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__39469),
            .DIN(N__39468),
            .DOUT(N__39467),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__39469),
            .PADOUT(N__39468),
            .PADIN(N__39467),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__39460),
            .DIN(N__39459),
            .DOUT(N__39458),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__39460),
            .PADOUT(N__39459),
            .PADIN(N__39458),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29117),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__39451),
            .DIN(N__39450),
            .DOUT(N__39449),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__39451),
            .PADOUT(N__39450),
            .PADIN(N__39449),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__39442),
            .DIN(N__39441),
            .DOUT(N__39440),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__39442),
            .PADOUT(N__39441),
            .PADIN(N__39440),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24735),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__39433),
            .DIN(N__39432),
            .DOUT(N__39431),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__39433),
            .PADOUT(N__39432),
            .PADIN(N__39431),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30945),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__39424),
            .DIN(N__39423),
            .DOUT(N__39422),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__39424),
            .PADOUT(N__39423),
            .PADIN(N__39422),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__39415),
            .DIN(N__39414),
            .DOUT(N__39413),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__39415),
            .PADOUT(N__39414),
            .PADIN(N__39413),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__39406),
            .DIN(N__39405),
            .DOUT(N__39404),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__39406),
            .PADOUT(N__39405),
            .PADIN(N__39404),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__39397),
            .DIN(N__39396),
            .DOUT(N__39395),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__39397),
            .PADOUT(N__39396),
            .PADIN(N__39395),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__39388),
            .DIN(N__39387),
            .DOUT(N__39386),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__39388),
            .PADOUT(N__39387),
            .PADIN(N__39386),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27675),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__39379),
            .DIN(N__39378),
            .DOUT(N__39377),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__39379),
            .PADOUT(N__39378),
            .PADIN(N__39377),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__39370),
            .DIN(N__39369),
            .DOUT(N__39368),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__39370),
            .PADOUT(N__39369),
            .PADIN(N__39368),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__39361),
            .DIN(N__39360),
            .DOUT(N__39359),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__39361),
            .PADOUT(N__39360),
            .PADIN(N__39359),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__39352),
            .DIN(N__39351),
            .DOUT(N__39350),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__39352),
            .PADOUT(N__39351),
            .PADIN(N__39350),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__39343),
            .DIN(N__39342),
            .DOUT(N__39341),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__39343),
            .PADOUT(N__39342),
            .PADIN(N__39341),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__39334),
            .DIN(N__39333),
            .DOUT(N__39332),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__39334),
            .PADOUT(N__39333),
            .PADIN(N__39332),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__39325),
            .DIN(N__39324),
            .DOUT(N__39323),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__39325),
            .PADOUT(N__39324),
            .PADIN(N__39323),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23952),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__39316),
            .DIN(N__39315),
            .DOUT(N__39314),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__39316),
            .PADOUT(N__39315),
            .PADIN(N__39314),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__9172 (
            .O(N__39297),
            .I(N__39289));
    InMux I__9171 (
            .O(N__39296),
            .I(N__39289));
    InMux I__9170 (
            .O(N__39295),
            .I(N__39277));
    InMux I__9169 (
            .O(N__39294),
            .I(N__39274));
    LocalMux I__9168 (
            .O(N__39289),
            .I(N__39269));
    InMux I__9167 (
            .O(N__39288),
            .I(N__39266));
    InMux I__9166 (
            .O(N__39287),
            .I(N__39263));
    InMux I__9165 (
            .O(N__39286),
            .I(N__39256));
    InMux I__9164 (
            .O(N__39285),
            .I(N__39256));
    InMux I__9163 (
            .O(N__39284),
            .I(N__39256));
    InMux I__9162 (
            .O(N__39283),
            .I(N__39249));
    InMux I__9161 (
            .O(N__39282),
            .I(N__39249));
    InMux I__9160 (
            .O(N__39281),
            .I(N__39249));
    InMux I__9159 (
            .O(N__39280),
            .I(N__39246));
    LocalMux I__9158 (
            .O(N__39277),
            .I(N__39243));
    LocalMux I__9157 (
            .O(N__39274),
            .I(N__39240));
    InMux I__9156 (
            .O(N__39273),
            .I(N__39237));
    InMux I__9155 (
            .O(N__39272),
            .I(N__39234));
    Sp12to4 I__9154 (
            .O(N__39269),
            .I(N__39231));
    LocalMux I__9153 (
            .O(N__39266),
            .I(N__39224));
    LocalMux I__9152 (
            .O(N__39263),
            .I(N__39224));
    LocalMux I__9151 (
            .O(N__39256),
            .I(N__39224));
    LocalMux I__9150 (
            .O(N__39249),
            .I(N__39219));
    LocalMux I__9149 (
            .O(N__39246),
            .I(N__39219));
    Span4Mux_v I__9148 (
            .O(N__39243),
            .I(N__39214));
    Span4Mux_h I__9147 (
            .O(N__39240),
            .I(N__39214));
    LocalMux I__9146 (
            .O(N__39237),
            .I(N__39209));
    LocalMux I__9145 (
            .O(N__39234),
            .I(N__39209));
    Span12Mux_v I__9144 (
            .O(N__39231),
            .I(N__39206));
    Span4Mux_v I__9143 (
            .O(N__39224),
            .I(N__39203));
    Span12Mux_v I__9142 (
            .O(N__39219),
            .I(N__39200));
    Span4Mux_v I__9141 (
            .O(N__39214),
            .I(N__39195));
    Span4Mux_v I__9140 (
            .O(N__39209),
            .I(N__39195));
    Odrv12 I__9139 (
            .O(N__39206),
            .I(gpio_fpga_soc_4));
    Odrv4 I__9138 (
            .O(N__39203),
            .I(gpio_fpga_soc_4));
    Odrv12 I__9137 (
            .O(N__39200),
            .I(gpio_fpga_soc_4));
    Odrv4 I__9136 (
            .O(N__39195),
            .I(gpio_fpga_soc_4));
    InMux I__9135 (
            .O(N__39186),
            .I(N__39172));
    CascadeMux I__9134 (
            .O(N__39185),
            .I(N__39162));
    CascadeMux I__9133 (
            .O(N__39184),
            .I(N__39155));
    InMux I__9132 (
            .O(N__39183),
            .I(N__39147));
    InMux I__9131 (
            .O(N__39182),
            .I(N__39147));
    InMux I__9130 (
            .O(N__39181),
            .I(N__39147));
    CascadeMux I__9129 (
            .O(N__39180),
            .I(N__39143));
    CascadeMux I__9128 (
            .O(N__39179),
            .I(N__39140));
    CascadeMux I__9127 (
            .O(N__39178),
            .I(N__39136));
    CascadeMux I__9126 (
            .O(N__39177),
            .I(N__39133));
    CascadeMux I__9125 (
            .O(N__39176),
            .I(N__39129));
    InMux I__9124 (
            .O(N__39175),
            .I(N__39124));
    LocalMux I__9123 (
            .O(N__39172),
            .I(N__39121));
    InMux I__9122 (
            .O(N__39171),
            .I(N__39118));
    InMux I__9121 (
            .O(N__39170),
            .I(N__39102));
    InMux I__9120 (
            .O(N__39169),
            .I(N__39102));
    InMux I__9119 (
            .O(N__39168),
            .I(N__39102));
    InMux I__9118 (
            .O(N__39167),
            .I(N__39102));
    InMux I__9117 (
            .O(N__39166),
            .I(N__39102));
    InMux I__9116 (
            .O(N__39165),
            .I(N__39102));
    InMux I__9115 (
            .O(N__39162),
            .I(N__39102));
    CascadeMux I__9114 (
            .O(N__39161),
            .I(N__39099));
    CascadeMux I__9113 (
            .O(N__39160),
            .I(N__39096));
    CascadeMux I__9112 (
            .O(N__39159),
            .I(N__39088));
    InMux I__9111 (
            .O(N__39158),
            .I(N__39077));
    InMux I__9110 (
            .O(N__39155),
            .I(N__39077));
    InMux I__9109 (
            .O(N__39154),
            .I(N__39077));
    LocalMux I__9108 (
            .O(N__39147),
            .I(N__39074));
    InMux I__9107 (
            .O(N__39146),
            .I(N__39061));
    InMux I__9106 (
            .O(N__39143),
            .I(N__39061));
    InMux I__9105 (
            .O(N__39140),
            .I(N__39061));
    InMux I__9104 (
            .O(N__39139),
            .I(N__39061));
    InMux I__9103 (
            .O(N__39136),
            .I(N__39061));
    InMux I__9102 (
            .O(N__39133),
            .I(N__39061));
    InMux I__9101 (
            .O(N__39132),
            .I(N__39048));
    InMux I__9100 (
            .O(N__39129),
            .I(N__39048));
    InMux I__9099 (
            .O(N__39128),
            .I(N__39045));
    InMux I__9098 (
            .O(N__39127),
            .I(N__39042));
    LocalMux I__9097 (
            .O(N__39124),
            .I(N__39035));
    Span4Mux_s2_h I__9096 (
            .O(N__39121),
            .I(N__39035));
    LocalMux I__9095 (
            .O(N__39118),
            .I(N__39035));
    InMux I__9094 (
            .O(N__39117),
            .I(N__39032));
    LocalMux I__9093 (
            .O(N__39102),
            .I(N__39029));
    InMux I__9092 (
            .O(N__39099),
            .I(N__39022));
    InMux I__9091 (
            .O(N__39096),
            .I(N__39022));
    InMux I__9090 (
            .O(N__39095),
            .I(N__39022));
    InMux I__9089 (
            .O(N__39094),
            .I(N__39019));
    CascadeMux I__9088 (
            .O(N__39093),
            .I(N__39016));
    CascadeMux I__9087 (
            .O(N__39092),
            .I(N__39013));
    InMux I__9086 (
            .O(N__39091),
            .I(N__39007));
    InMux I__9085 (
            .O(N__39088),
            .I(N__39007));
    InMux I__9084 (
            .O(N__39087),
            .I(N__39002));
    InMux I__9083 (
            .O(N__39086),
            .I(N__39002));
    CascadeMux I__9082 (
            .O(N__39085),
            .I(N__38998));
    InMux I__9081 (
            .O(N__39084),
            .I(N__38995));
    LocalMux I__9080 (
            .O(N__39077),
            .I(N__38992));
    Span4Mux_s2_v I__9079 (
            .O(N__39074),
            .I(N__38987));
    LocalMux I__9078 (
            .O(N__39061),
            .I(N__38987));
    CascadeMux I__9077 (
            .O(N__39060),
            .I(N__38984));
    InMux I__9076 (
            .O(N__39059),
            .I(N__38971));
    InMux I__9075 (
            .O(N__39058),
            .I(N__38971));
    InMux I__9074 (
            .O(N__39057),
            .I(N__38971));
    InMux I__9073 (
            .O(N__39056),
            .I(N__38971));
    InMux I__9072 (
            .O(N__39055),
            .I(N__38968));
    InMux I__9071 (
            .O(N__39054),
            .I(N__38964));
    InMux I__9070 (
            .O(N__39053),
            .I(N__38961));
    LocalMux I__9069 (
            .O(N__39048),
            .I(N__38958));
    LocalMux I__9068 (
            .O(N__39045),
            .I(N__38945));
    LocalMux I__9067 (
            .O(N__39042),
            .I(N__38945));
    Span4Mux_v I__9066 (
            .O(N__39035),
            .I(N__38945));
    LocalMux I__9065 (
            .O(N__39032),
            .I(N__38945));
    Span4Mux_s2_h I__9064 (
            .O(N__39029),
            .I(N__38945));
    LocalMux I__9063 (
            .O(N__39022),
            .I(N__38945));
    LocalMux I__9062 (
            .O(N__39019),
            .I(N__38942));
    InMux I__9061 (
            .O(N__39016),
            .I(N__38935));
    InMux I__9060 (
            .O(N__39013),
            .I(N__38935));
    InMux I__9059 (
            .O(N__39012),
            .I(N__38935));
    LocalMux I__9058 (
            .O(N__39007),
            .I(N__38930));
    LocalMux I__9057 (
            .O(N__39002),
            .I(N__38930));
    InMux I__9056 (
            .O(N__39001),
            .I(N__38925));
    InMux I__9055 (
            .O(N__38998),
            .I(N__38925));
    LocalMux I__9054 (
            .O(N__38995),
            .I(N__38918));
    Span4Mux_v I__9053 (
            .O(N__38992),
            .I(N__38918));
    Span4Mux_v I__9052 (
            .O(N__38987),
            .I(N__38918));
    InMux I__9051 (
            .O(N__38984),
            .I(N__38913));
    InMux I__9050 (
            .O(N__38983),
            .I(N__38913));
    InMux I__9049 (
            .O(N__38982),
            .I(N__38910));
    InMux I__9048 (
            .O(N__38981),
            .I(N__38905));
    InMux I__9047 (
            .O(N__38980),
            .I(N__38905));
    LocalMux I__9046 (
            .O(N__38971),
            .I(N__38900));
    LocalMux I__9045 (
            .O(N__38968),
            .I(N__38900));
    InMux I__9044 (
            .O(N__38967),
            .I(N__38897));
    LocalMux I__9043 (
            .O(N__38964),
            .I(N__38888));
    LocalMux I__9042 (
            .O(N__38961),
            .I(N__38888));
    Span4Mux_s2_h I__9041 (
            .O(N__38958),
            .I(N__38888));
    Span4Mux_v I__9040 (
            .O(N__38945),
            .I(N__38888));
    Span4Mux_v I__9039 (
            .O(N__38942),
            .I(N__38877));
    LocalMux I__9038 (
            .O(N__38935),
            .I(N__38877));
    Span4Mux_h I__9037 (
            .O(N__38930),
            .I(N__38877));
    LocalMux I__9036 (
            .O(N__38925),
            .I(N__38877));
    Span4Mux_h I__9035 (
            .O(N__38918),
            .I(N__38877));
    LocalMux I__9034 (
            .O(N__38913),
            .I(\b2v_inst11.func_state ));
    LocalMux I__9033 (
            .O(N__38910),
            .I(\b2v_inst11.func_state ));
    LocalMux I__9032 (
            .O(N__38905),
            .I(\b2v_inst11.func_state ));
    Odrv12 I__9031 (
            .O(N__38900),
            .I(\b2v_inst11.func_state ));
    LocalMux I__9030 (
            .O(N__38897),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__9029 (
            .O(N__38888),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__9028 (
            .O(N__38877),
            .I(\b2v_inst11.func_state ));
    CascadeMux I__9027 (
            .O(N__38862),
            .I(\b2v_inst11.g2_3Z0Z_0_cascade_ ));
    CascadeMux I__9026 (
            .O(N__38859),
            .I(N__38855));
    CascadeMux I__9025 (
            .O(N__38858),
            .I(N__38852));
    InMux I__9024 (
            .O(N__38855),
            .I(N__38839));
    InMux I__9023 (
            .O(N__38852),
            .I(N__38839));
    InMux I__9022 (
            .O(N__38851),
            .I(N__38839));
    InMux I__9021 (
            .O(N__38850),
            .I(N__38836));
    CascadeMux I__9020 (
            .O(N__38849),
            .I(N__38833));
    InMux I__9019 (
            .O(N__38848),
            .I(N__38828));
    InMux I__9018 (
            .O(N__38847),
            .I(N__38825));
    InMux I__9017 (
            .O(N__38846),
            .I(N__38822));
    LocalMux I__9016 (
            .O(N__38839),
            .I(N__38819));
    LocalMux I__9015 (
            .O(N__38836),
            .I(N__38816));
    InMux I__9014 (
            .O(N__38833),
            .I(N__38809));
    InMux I__9013 (
            .O(N__38832),
            .I(N__38804));
    InMux I__9012 (
            .O(N__38831),
            .I(N__38804));
    LocalMux I__9011 (
            .O(N__38828),
            .I(N__38798));
    LocalMux I__9010 (
            .O(N__38825),
            .I(N__38791));
    LocalMux I__9009 (
            .O(N__38822),
            .I(N__38791));
    Span4Mux_v I__9008 (
            .O(N__38819),
            .I(N__38791));
    Span4Mux_h I__9007 (
            .O(N__38816),
            .I(N__38788));
    InMux I__9006 (
            .O(N__38815),
            .I(N__38781));
    InMux I__9005 (
            .O(N__38814),
            .I(N__38781));
    InMux I__9004 (
            .O(N__38813),
            .I(N__38781));
    InMux I__9003 (
            .O(N__38812),
            .I(N__38778));
    LocalMux I__9002 (
            .O(N__38809),
            .I(N__38773));
    LocalMux I__9001 (
            .O(N__38804),
            .I(N__38773));
    InMux I__9000 (
            .O(N__38803),
            .I(N__38766));
    InMux I__8999 (
            .O(N__38802),
            .I(N__38766));
    InMux I__8998 (
            .O(N__38801),
            .I(N__38766));
    Span4Mux_h I__8997 (
            .O(N__38798),
            .I(N__38761));
    Span4Mux_h I__8996 (
            .O(N__38791),
            .I(N__38761));
    Span4Mux_v I__8995 (
            .O(N__38788),
            .I(N__38758));
    LocalMux I__8994 (
            .O(N__38781),
            .I(N__38749));
    LocalMux I__8993 (
            .O(N__38778),
            .I(N__38749));
    Span12Mux_s2_v I__8992 (
            .O(N__38773),
            .I(N__38749));
    LocalMux I__8991 (
            .O(N__38766),
            .I(N__38749));
    Odrv4 I__8990 (
            .O(N__38761),
            .I(\b2v_inst11.N_200_i ));
    Odrv4 I__8989 (
            .O(N__38758),
            .I(\b2v_inst11.N_200_i ));
    Odrv12 I__8988 (
            .O(N__38749),
            .I(\b2v_inst11.N_200_i ));
    CascadeMux I__8987 (
            .O(N__38742),
            .I(N__38739));
    InMux I__8986 (
            .O(N__38739),
            .I(N__38736));
    LocalMux I__8985 (
            .O(N__38736),
            .I(N__38733));
    Odrv12 I__8984 (
            .O(N__38733),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_0 ));
    InMux I__8983 (
            .O(N__38730),
            .I(N__38726));
    CascadeMux I__8982 (
            .O(N__38729),
            .I(N__38719));
    LocalMux I__8981 (
            .O(N__38726),
            .I(N__38714));
    InMux I__8980 (
            .O(N__38725),
            .I(N__38711));
    InMux I__8979 (
            .O(N__38724),
            .I(N__38708));
    CascadeMux I__8978 (
            .O(N__38723),
            .I(N__38705));
    InMux I__8977 (
            .O(N__38722),
            .I(N__38697));
    InMux I__8976 (
            .O(N__38719),
            .I(N__38697));
    InMux I__8975 (
            .O(N__38718),
            .I(N__38697));
    CascadeMux I__8974 (
            .O(N__38717),
            .I(N__38694));
    Span4Mux_v I__8973 (
            .O(N__38714),
            .I(N__38688));
    LocalMux I__8972 (
            .O(N__38711),
            .I(N__38688));
    LocalMux I__8971 (
            .O(N__38708),
            .I(N__38685));
    InMux I__8970 (
            .O(N__38705),
            .I(N__38680));
    InMux I__8969 (
            .O(N__38704),
            .I(N__38680));
    LocalMux I__8968 (
            .O(N__38697),
            .I(N__38671));
    InMux I__8967 (
            .O(N__38694),
            .I(N__38666));
    InMux I__8966 (
            .O(N__38693),
            .I(N__38666));
    Span4Mux_h I__8965 (
            .O(N__38688),
            .I(N__38659));
    Span4Mux_h I__8964 (
            .O(N__38685),
            .I(N__38659));
    LocalMux I__8963 (
            .O(N__38680),
            .I(N__38659));
    InMux I__8962 (
            .O(N__38679),
            .I(N__38652));
    InMux I__8961 (
            .O(N__38678),
            .I(N__38652));
    InMux I__8960 (
            .O(N__38677),
            .I(N__38652));
    CascadeMux I__8959 (
            .O(N__38676),
            .I(N__38649));
    CascadeMux I__8958 (
            .O(N__38675),
            .I(N__38646));
    CascadeMux I__8957 (
            .O(N__38674),
            .I(N__38642));
    Span4Mux_v I__8956 (
            .O(N__38671),
            .I(N__38632));
    LocalMux I__8955 (
            .O(N__38666),
            .I(N__38632));
    Span4Mux_s3_h I__8954 (
            .O(N__38659),
            .I(N__38632));
    LocalMux I__8953 (
            .O(N__38652),
            .I(N__38632));
    InMux I__8952 (
            .O(N__38649),
            .I(N__38627));
    InMux I__8951 (
            .O(N__38646),
            .I(N__38627));
    InMux I__8950 (
            .O(N__38645),
            .I(N__38622));
    InMux I__8949 (
            .O(N__38642),
            .I(N__38622));
    InMux I__8948 (
            .O(N__38641),
            .I(N__38619));
    Span4Mux_v I__8947 (
            .O(N__38632),
            .I(N__38616));
    LocalMux I__8946 (
            .O(N__38627),
            .I(N__38608));
    LocalMux I__8945 (
            .O(N__38622),
            .I(N__38608));
    LocalMux I__8944 (
            .O(N__38619),
            .I(N__38608));
    IoSpan4Mux I__8943 (
            .O(N__38616),
            .I(N__38605));
    InMux I__8942 (
            .O(N__38615),
            .I(N__38602));
    Span4Mux_v I__8941 (
            .O(N__38608),
            .I(N__38595));
    Span4Mux_s1_h I__8940 (
            .O(N__38605),
            .I(N__38595));
    LocalMux I__8939 (
            .O(N__38602),
            .I(N__38595));
    Span4Mux_h I__8938 (
            .O(N__38595),
            .I(N__38592));
    Span4Mux_v I__8937 (
            .O(N__38592),
            .I(N__38584));
    InMux I__8936 (
            .O(N__38591),
            .I(N__38579));
    InMux I__8935 (
            .O(N__38590),
            .I(N__38579));
    InMux I__8934 (
            .O(N__38589),
            .I(N__38572));
    InMux I__8933 (
            .O(N__38588),
            .I(N__38572));
    InMux I__8932 (
            .O(N__38587),
            .I(N__38572));
    Odrv4 I__8931 (
            .O(N__38584),
            .I(slp_s3n));
    LocalMux I__8930 (
            .O(N__38579),
            .I(slp_s3n));
    LocalMux I__8929 (
            .O(N__38572),
            .I(slp_s3n));
    CascadeMux I__8928 (
            .O(N__38565),
            .I(N__38557));
    InMux I__8927 (
            .O(N__38564),
            .I(N__38547));
    InMux I__8926 (
            .O(N__38563),
            .I(N__38547));
    InMux I__8925 (
            .O(N__38562),
            .I(N__38544));
    InMux I__8924 (
            .O(N__38561),
            .I(N__38539));
    InMux I__8923 (
            .O(N__38560),
            .I(N__38539));
    InMux I__8922 (
            .O(N__38557),
            .I(N__38530));
    InMux I__8921 (
            .O(N__38556),
            .I(N__38530));
    InMux I__8920 (
            .O(N__38555),
            .I(N__38530));
    InMux I__8919 (
            .O(N__38554),
            .I(N__38530));
    InMux I__8918 (
            .O(N__38553),
            .I(N__38518));
    InMux I__8917 (
            .O(N__38552),
            .I(N__38518));
    LocalMux I__8916 (
            .O(N__38547),
            .I(N__38510));
    LocalMux I__8915 (
            .O(N__38544),
            .I(N__38510));
    LocalMux I__8914 (
            .O(N__38539),
            .I(N__38505));
    LocalMux I__8913 (
            .O(N__38530),
            .I(N__38505));
    InMux I__8912 (
            .O(N__38529),
            .I(N__38502));
    InMux I__8911 (
            .O(N__38528),
            .I(N__38499));
    InMux I__8910 (
            .O(N__38527),
            .I(N__38488));
    InMux I__8909 (
            .O(N__38526),
            .I(N__38488));
    InMux I__8908 (
            .O(N__38525),
            .I(N__38488));
    InMux I__8907 (
            .O(N__38524),
            .I(N__38488));
    InMux I__8906 (
            .O(N__38523),
            .I(N__38488));
    LocalMux I__8905 (
            .O(N__38518),
            .I(N__38485));
    InMux I__8904 (
            .O(N__38517),
            .I(N__38477));
    InMux I__8903 (
            .O(N__38516),
            .I(N__38477));
    InMux I__8902 (
            .O(N__38515),
            .I(N__38477));
    Span4Mux_v I__8901 (
            .O(N__38510),
            .I(N__38472));
    Span4Mux_v I__8900 (
            .O(N__38505),
            .I(N__38472));
    LocalMux I__8899 (
            .O(N__38502),
            .I(N__38469));
    LocalMux I__8898 (
            .O(N__38499),
            .I(N__38466));
    LocalMux I__8897 (
            .O(N__38488),
            .I(N__38463));
    Span4Mux_v I__8896 (
            .O(N__38485),
            .I(N__38460));
    InMux I__8895 (
            .O(N__38484),
            .I(N__38457));
    LocalMux I__8894 (
            .O(N__38477),
            .I(N__38454));
    Span4Mux_h I__8893 (
            .O(N__38472),
            .I(N__38447));
    Span4Mux_s3_h I__8892 (
            .O(N__38469),
            .I(N__38447));
    Span4Mux_h I__8891 (
            .O(N__38466),
            .I(N__38447));
    IoSpan4Mux I__8890 (
            .O(N__38463),
            .I(N__38444));
    Sp12to4 I__8889 (
            .O(N__38460),
            .I(N__38439));
    LocalMux I__8888 (
            .O(N__38457),
            .I(N__38439));
    Span12Mux_s8_h I__8887 (
            .O(N__38454),
            .I(N__38436));
    Span4Mux_v I__8886 (
            .O(N__38447),
            .I(N__38433));
    IoSpan4Mux I__8885 (
            .O(N__38444),
            .I(N__38430));
    Span12Mux_s8_h I__8884 (
            .O(N__38439),
            .I(N__38427));
    Odrv12 I__8883 (
            .O(N__38436),
            .I(slp_s4n));
    Odrv4 I__8882 (
            .O(N__38433),
            .I(slp_s4n));
    Odrv4 I__8881 (
            .O(N__38430),
            .I(slp_s4n));
    Odrv12 I__8880 (
            .O(N__38427),
            .I(slp_s4n));
    CascadeMux I__8879 (
            .O(N__38418),
            .I(N__38413));
    CascadeMux I__8878 (
            .O(N__38417),
            .I(N__38410));
    CascadeMux I__8877 (
            .O(N__38416),
            .I(N__38405));
    InMux I__8876 (
            .O(N__38413),
            .I(N__38399));
    InMux I__8875 (
            .O(N__38410),
            .I(N__38399));
    InMux I__8874 (
            .O(N__38409),
            .I(N__38392));
    InMux I__8873 (
            .O(N__38408),
            .I(N__38392));
    InMux I__8872 (
            .O(N__38405),
            .I(N__38392));
    InMux I__8871 (
            .O(N__38404),
            .I(N__38388));
    LocalMux I__8870 (
            .O(N__38399),
            .I(N__38383));
    LocalMux I__8869 (
            .O(N__38392),
            .I(N__38383));
    CascadeMux I__8868 (
            .O(N__38391),
            .I(N__38380));
    LocalMux I__8867 (
            .O(N__38388),
            .I(N__38377));
    Span4Mux_h I__8866 (
            .O(N__38383),
            .I(N__38374));
    InMux I__8865 (
            .O(N__38380),
            .I(N__38371));
    Span4Mux_v I__8864 (
            .O(N__38377),
            .I(N__38368));
    Sp12to4 I__8863 (
            .O(N__38374),
            .I(N__38363));
    LocalMux I__8862 (
            .O(N__38371),
            .I(N__38363));
    Span4Mux_h I__8861 (
            .O(N__38368),
            .I(N__38360));
    Span12Mux_s10_v I__8860 (
            .O(N__38363),
            .I(N__38357));
    Odrv4 I__8859 (
            .O(N__38360),
            .I(\b2v_inst11.N_161 ));
    Odrv12 I__8858 (
            .O(N__38357),
            .I(\b2v_inst11.N_161 ));
    CascadeMux I__8857 (
            .O(N__38352),
            .I(N__38348));
    CascadeMux I__8856 (
            .O(N__38351),
            .I(N__38333));
    InMux I__8855 (
            .O(N__38348),
            .I(N__38321));
    InMux I__8854 (
            .O(N__38347),
            .I(N__38321));
    InMux I__8853 (
            .O(N__38346),
            .I(N__38321));
    InMux I__8852 (
            .O(N__38345),
            .I(N__38316));
    InMux I__8851 (
            .O(N__38344),
            .I(N__38316));
    CascadeMux I__8850 (
            .O(N__38343),
            .I(N__38313));
    InMux I__8849 (
            .O(N__38342),
            .I(N__38306));
    CascadeMux I__8848 (
            .O(N__38341),
            .I(N__38303));
    InMux I__8847 (
            .O(N__38340),
            .I(N__38296));
    InMux I__8846 (
            .O(N__38339),
            .I(N__38296));
    InMux I__8845 (
            .O(N__38338),
            .I(N__38296));
    InMux I__8844 (
            .O(N__38337),
            .I(N__38292));
    InMux I__8843 (
            .O(N__38336),
            .I(N__38287));
    InMux I__8842 (
            .O(N__38333),
            .I(N__38287));
    InMux I__8841 (
            .O(N__38332),
            .I(N__38280));
    InMux I__8840 (
            .O(N__38331),
            .I(N__38280));
    InMux I__8839 (
            .O(N__38330),
            .I(N__38280));
    InMux I__8838 (
            .O(N__38329),
            .I(N__38275));
    InMux I__8837 (
            .O(N__38328),
            .I(N__38275));
    LocalMux I__8836 (
            .O(N__38321),
            .I(N__38271));
    LocalMux I__8835 (
            .O(N__38316),
            .I(N__38268));
    InMux I__8834 (
            .O(N__38313),
            .I(N__38259));
    InMux I__8833 (
            .O(N__38312),
            .I(N__38259));
    InMux I__8832 (
            .O(N__38311),
            .I(N__38259));
    InMux I__8831 (
            .O(N__38310),
            .I(N__38259));
    InMux I__8830 (
            .O(N__38309),
            .I(N__38254));
    LocalMux I__8829 (
            .O(N__38306),
            .I(N__38251));
    InMux I__8828 (
            .O(N__38303),
            .I(N__38248));
    LocalMux I__8827 (
            .O(N__38296),
            .I(N__38245));
    InMux I__8826 (
            .O(N__38295),
            .I(N__38242));
    LocalMux I__8825 (
            .O(N__38292),
            .I(N__38237));
    LocalMux I__8824 (
            .O(N__38287),
            .I(N__38237));
    LocalMux I__8823 (
            .O(N__38280),
            .I(N__38232));
    LocalMux I__8822 (
            .O(N__38275),
            .I(N__38232));
    InMux I__8821 (
            .O(N__38274),
            .I(N__38229));
    Span4Mux_h I__8820 (
            .O(N__38271),
            .I(N__38220));
    Span4Mux_v I__8819 (
            .O(N__38268),
            .I(N__38220));
    LocalMux I__8818 (
            .O(N__38259),
            .I(N__38220));
    InMux I__8817 (
            .O(N__38258),
            .I(N__38215));
    InMux I__8816 (
            .O(N__38257),
            .I(N__38215));
    LocalMux I__8815 (
            .O(N__38254),
            .I(N__38204));
    Span4Mux_h I__8814 (
            .O(N__38251),
            .I(N__38204));
    LocalMux I__8813 (
            .O(N__38248),
            .I(N__38204));
    Span4Mux_s1_v I__8812 (
            .O(N__38245),
            .I(N__38204));
    LocalMux I__8811 (
            .O(N__38242),
            .I(N__38204));
    Span4Mux_v I__8810 (
            .O(N__38237),
            .I(N__38197));
    Span4Mux_v I__8809 (
            .O(N__38232),
            .I(N__38197));
    LocalMux I__8808 (
            .O(N__38229),
            .I(N__38197));
    InMux I__8807 (
            .O(N__38228),
            .I(N__38194));
    InMux I__8806 (
            .O(N__38227),
            .I(N__38191));
    Span4Mux_v I__8805 (
            .O(N__38220),
            .I(N__38188));
    LocalMux I__8804 (
            .O(N__38215),
            .I(N__38183));
    Span4Mux_v I__8803 (
            .O(N__38204),
            .I(N__38183));
    Span4Mux_v I__8802 (
            .O(N__38197),
            .I(N__38180));
    LocalMux I__8801 (
            .O(N__38194),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    LocalMux I__8800 (
            .O(N__38191),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__8799 (
            .O(N__38188),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__8798 (
            .O(N__38183),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__8797 (
            .O(N__38180),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    CascadeMux I__8796 (
            .O(N__38169),
            .I(N__38163));
    InMux I__8795 (
            .O(N__38168),
            .I(N__38155));
    InMux I__8794 (
            .O(N__38167),
            .I(N__38145));
    InMux I__8793 (
            .O(N__38166),
            .I(N__38145));
    InMux I__8792 (
            .O(N__38163),
            .I(N__38145));
    InMux I__8791 (
            .O(N__38162),
            .I(N__38145));
    InMux I__8790 (
            .O(N__38161),
            .I(N__38140));
    InMux I__8789 (
            .O(N__38160),
            .I(N__38140));
    InMux I__8788 (
            .O(N__38159),
            .I(N__38137));
    InMux I__8787 (
            .O(N__38158),
            .I(N__38132));
    LocalMux I__8786 (
            .O(N__38155),
            .I(N__38127));
    InMux I__8785 (
            .O(N__38154),
            .I(N__38124));
    LocalMux I__8784 (
            .O(N__38145),
            .I(N__38118));
    LocalMux I__8783 (
            .O(N__38140),
            .I(N__38115));
    LocalMux I__8782 (
            .O(N__38137),
            .I(N__38112));
    InMux I__8781 (
            .O(N__38136),
            .I(N__38109));
    CascadeMux I__8780 (
            .O(N__38135),
            .I(N__38103));
    LocalMux I__8779 (
            .O(N__38132),
            .I(N__38100));
    InMux I__8778 (
            .O(N__38131),
            .I(N__38095));
    InMux I__8777 (
            .O(N__38130),
            .I(N__38095));
    Span4Mux_h I__8776 (
            .O(N__38127),
            .I(N__38092));
    LocalMux I__8775 (
            .O(N__38124),
            .I(N__38089));
    InMux I__8774 (
            .O(N__38123),
            .I(N__38086));
    InMux I__8773 (
            .O(N__38122),
            .I(N__38081));
    InMux I__8772 (
            .O(N__38121),
            .I(N__38081));
    Span4Mux_s2_v I__8771 (
            .O(N__38118),
            .I(N__38076));
    Span4Mux_v I__8770 (
            .O(N__38115),
            .I(N__38076));
    Span12Mux_v I__8769 (
            .O(N__38112),
            .I(N__38071));
    LocalMux I__8768 (
            .O(N__38109),
            .I(N__38071));
    InMux I__8767 (
            .O(N__38108),
            .I(N__38064));
    InMux I__8766 (
            .O(N__38107),
            .I(N__38064));
    InMux I__8765 (
            .O(N__38106),
            .I(N__38064));
    InMux I__8764 (
            .O(N__38103),
            .I(N__38061));
    Span4Mux_v I__8763 (
            .O(N__38100),
            .I(N__38054));
    LocalMux I__8762 (
            .O(N__38095),
            .I(N__38054));
    Span4Mux_h I__8761 (
            .O(N__38092),
            .I(N__38054));
    Odrv4 I__8760 (
            .O(N__38089),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__8759 (
            .O(N__38086),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__8758 (
            .O(N__38081),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__8757 (
            .O(N__38076),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv12 I__8756 (
            .O(N__38071),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__8755 (
            .O(N__38064),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__8754 (
            .O(N__38061),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__8753 (
            .O(N__38054),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    CascadeMux I__8752 (
            .O(N__38037),
            .I(N__38024));
    InMux I__8751 (
            .O(N__38036),
            .I(N__38019));
    InMux I__8750 (
            .O(N__38035),
            .I(N__38014));
    InMux I__8749 (
            .O(N__38034),
            .I(N__38014));
    CascadeMux I__8748 (
            .O(N__38033),
            .I(N__38011));
    InMux I__8747 (
            .O(N__38032),
            .I(N__38008));
    InMux I__8746 (
            .O(N__38031),
            .I(N__38003));
    InMux I__8745 (
            .O(N__38030),
            .I(N__38003));
    InMux I__8744 (
            .O(N__38029),
            .I(N__37994));
    InMux I__8743 (
            .O(N__38028),
            .I(N__37994));
    InMux I__8742 (
            .O(N__38027),
            .I(N__37994));
    InMux I__8741 (
            .O(N__38024),
            .I(N__37994));
    InMux I__8740 (
            .O(N__38023),
            .I(N__37991));
    CascadeMux I__8739 (
            .O(N__38022),
            .I(N__37988));
    LocalMux I__8738 (
            .O(N__38019),
            .I(N__37985));
    LocalMux I__8737 (
            .O(N__38014),
            .I(N__37982));
    InMux I__8736 (
            .O(N__38011),
            .I(N__37977));
    LocalMux I__8735 (
            .O(N__38008),
            .I(N__37974));
    LocalMux I__8734 (
            .O(N__38003),
            .I(N__37969));
    LocalMux I__8733 (
            .O(N__37994),
            .I(N__37969));
    LocalMux I__8732 (
            .O(N__37991),
            .I(N__37966));
    InMux I__8731 (
            .O(N__37988),
            .I(N__37963));
    Span12Mux_s10_v I__8730 (
            .O(N__37985),
            .I(N__37958));
    Span12Mux_s5_v I__8729 (
            .O(N__37982),
            .I(N__37958));
    InMux I__8728 (
            .O(N__37981),
            .I(N__37953));
    InMux I__8727 (
            .O(N__37980),
            .I(N__37953));
    LocalMux I__8726 (
            .O(N__37977),
            .I(N__37942));
    Span4Mux_h I__8725 (
            .O(N__37974),
            .I(N__37942));
    Span4Mux_s3_v I__8724 (
            .O(N__37969),
            .I(N__37942));
    Span4Mux_h I__8723 (
            .O(N__37966),
            .I(N__37942));
    LocalMux I__8722 (
            .O(N__37963),
            .I(N__37942));
    Odrv12 I__8721 (
            .O(N__37958),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    LocalMux I__8720 (
            .O(N__37953),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__8719 (
            .O(N__37942),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    CascadeMux I__8718 (
            .O(N__37935),
            .I(N__37931));
    CascadeMux I__8717 (
            .O(N__37934),
            .I(N__37924));
    InMux I__8716 (
            .O(N__37931),
            .I(N__37920));
    InMux I__8715 (
            .O(N__37930),
            .I(N__37917));
    CascadeMux I__8714 (
            .O(N__37929),
            .I(N__37912));
    InMux I__8713 (
            .O(N__37928),
            .I(N__37907));
    InMux I__8712 (
            .O(N__37927),
            .I(N__37904));
    InMux I__8711 (
            .O(N__37924),
            .I(N__37899));
    InMux I__8710 (
            .O(N__37923),
            .I(N__37899));
    LocalMux I__8709 (
            .O(N__37920),
            .I(N__37896));
    LocalMux I__8708 (
            .O(N__37917),
            .I(N__37893));
    InMux I__8707 (
            .O(N__37916),
            .I(N__37888));
    InMux I__8706 (
            .O(N__37915),
            .I(N__37888));
    InMux I__8705 (
            .O(N__37912),
            .I(N__37885));
    InMux I__8704 (
            .O(N__37911),
            .I(N__37882));
    CascadeMux I__8703 (
            .O(N__37910),
            .I(N__37878));
    LocalMux I__8702 (
            .O(N__37907),
            .I(N__37865));
    LocalMux I__8701 (
            .O(N__37904),
            .I(N__37865));
    LocalMux I__8700 (
            .O(N__37899),
            .I(N__37862));
    Span4Mux_v I__8699 (
            .O(N__37896),
            .I(N__37855));
    Span4Mux_v I__8698 (
            .O(N__37893),
            .I(N__37855));
    LocalMux I__8697 (
            .O(N__37888),
            .I(N__37855));
    LocalMux I__8696 (
            .O(N__37885),
            .I(N__37850));
    LocalMux I__8695 (
            .O(N__37882),
            .I(N__37850));
    InMux I__8694 (
            .O(N__37881),
            .I(N__37843));
    InMux I__8693 (
            .O(N__37878),
            .I(N__37843));
    InMux I__8692 (
            .O(N__37877),
            .I(N__37843));
    InMux I__8691 (
            .O(N__37876),
            .I(N__37840));
    CascadeMux I__8690 (
            .O(N__37875),
            .I(N__37837));
    InMux I__8689 (
            .O(N__37874),
            .I(N__37832));
    InMux I__8688 (
            .O(N__37873),
            .I(N__37832));
    InMux I__8687 (
            .O(N__37872),
            .I(N__37825));
    InMux I__8686 (
            .O(N__37871),
            .I(N__37825));
    InMux I__8685 (
            .O(N__37870),
            .I(N__37825));
    Span4Mux_s1_v I__8684 (
            .O(N__37865),
            .I(N__37820));
    Span4Mux_v I__8683 (
            .O(N__37862),
            .I(N__37820));
    Span4Mux_h I__8682 (
            .O(N__37855),
            .I(N__37817));
    Span4Mux_v I__8681 (
            .O(N__37850),
            .I(N__37812));
    LocalMux I__8680 (
            .O(N__37843),
            .I(N__37812));
    LocalMux I__8679 (
            .O(N__37840),
            .I(N__37809));
    InMux I__8678 (
            .O(N__37837),
            .I(N__37806));
    LocalMux I__8677 (
            .O(N__37832),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__8676 (
            .O(N__37825),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__8675 (
            .O(N__37820),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__8674 (
            .O(N__37817),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__8673 (
            .O(N__37812),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv12 I__8672 (
            .O(N__37809),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__8671 (
            .O(N__37806),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    InMux I__8670 (
            .O(N__37791),
            .I(N__37788));
    LocalMux I__8669 (
            .O(N__37788),
            .I(\b2v_inst11.un1_i2_mux_0 ));
    InMux I__8668 (
            .O(N__37785),
            .I(N__37782));
    LocalMux I__8667 (
            .O(N__37782),
            .I(\b2v_inst11.un1_N_5 ));
    CascadeMux I__8666 (
            .O(N__37779),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_ ));
    InMux I__8665 (
            .O(N__37776),
            .I(N__37773));
    LocalMux I__8664 (
            .O(N__37773),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_12 ));
    CascadeMux I__8663 (
            .O(N__37770),
            .I(N__37758));
    CascadeMux I__8662 (
            .O(N__37769),
            .I(N__37753));
    InMux I__8661 (
            .O(N__37768),
            .I(N__37750));
    InMux I__8660 (
            .O(N__37767),
            .I(N__37743));
    InMux I__8659 (
            .O(N__37766),
            .I(N__37740));
    InMux I__8658 (
            .O(N__37765),
            .I(N__37731));
    InMux I__8657 (
            .O(N__37764),
            .I(N__37731));
    InMux I__8656 (
            .O(N__37763),
            .I(N__37731));
    InMux I__8655 (
            .O(N__37762),
            .I(N__37731));
    InMux I__8654 (
            .O(N__37761),
            .I(N__37724));
    InMux I__8653 (
            .O(N__37758),
            .I(N__37724));
    InMux I__8652 (
            .O(N__37757),
            .I(N__37724));
    InMux I__8651 (
            .O(N__37756),
            .I(N__37721));
    InMux I__8650 (
            .O(N__37753),
            .I(N__37718));
    LocalMux I__8649 (
            .O(N__37750),
            .I(N__37715));
    InMux I__8648 (
            .O(N__37749),
            .I(N__37706));
    InMux I__8647 (
            .O(N__37748),
            .I(N__37706));
    InMux I__8646 (
            .O(N__37747),
            .I(N__37706));
    InMux I__8645 (
            .O(N__37746),
            .I(N__37706));
    LocalMux I__8644 (
            .O(N__37743),
            .I(N__37701));
    LocalMux I__8643 (
            .O(N__37740),
            .I(N__37698));
    LocalMux I__8642 (
            .O(N__37731),
            .I(N__37693));
    LocalMux I__8641 (
            .O(N__37724),
            .I(N__37693));
    LocalMux I__8640 (
            .O(N__37721),
            .I(N__37690));
    LocalMux I__8639 (
            .O(N__37718),
            .I(N__37687));
    Span4Mux_v I__8638 (
            .O(N__37715),
            .I(N__37682));
    LocalMux I__8637 (
            .O(N__37706),
            .I(N__37682));
    InMux I__8636 (
            .O(N__37705),
            .I(N__37677));
    InMux I__8635 (
            .O(N__37704),
            .I(N__37677));
    Span4Mux_v I__8634 (
            .O(N__37701),
            .I(N__37670));
    Span4Mux_v I__8633 (
            .O(N__37698),
            .I(N__37670));
    Span4Mux_v I__8632 (
            .O(N__37693),
            .I(N__37670));
    Span4Mux_s2_v I__8631 (
            .O(N__37690),
            .I(N__37665));
    Span4Mux_s2_h I__8630 (
            .O(N__37687),
            .I(N__37665));
    Odrv4 I__8629 (
            .O(N__37682),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__8628 (
            .O(N__37677),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__8627 (
            .O(N__37670),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__8626 (
            .O(N__37665),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    CascadeMux I__8625 (
            .O(N__37656),
            .I(\b2v_inst11.un1_dutycycle_53_s_9_sf_cascade_ ));
    CascadeMux I__8624 (
            .O(N__37653),
            .I(N__37650));
    InMux I__8623 (
            .O(N__37650),
            .I(N__37647));
    LocalMux I__8622 (
            .O(N__37647),
            .I(N__37644));
    Odrv12 I__8621 (
            .O(N__37644),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_12 ));
    InMux I__8620 (
            .O(N__37641),
            .I(N__37638));
    LocalMux I__8619 (
            .O(N__37638),
            .I(N__37635));
    Span4Mux_h I__8618 (
            .O(N__37635),
            .I(N__37632));
    Span4Mux_v I__8617 (
            .O(N__37632),
            .I(N__37629));
    Span4Mux_v I__8616 (
            .O(N__37629),
            .I(N__37626));
    Odrv4 I__8615 (
            .O(N__37626),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_1 ));
    CascadeMux I__8614 (
            .O(N__37623),
            .I(\b2v_inst11.N_371_cascade_ ));
    CascadeMux I__8613 (
            .O(N__37620),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_cascade_ ));
    InMux I__8612 (
            .O(N__37617),
            .I(N__37614));
    LocalMux I__8611 (
            .O(N__37614),
            .I(N__37611));
    Span4Mux_v I__8610 (
            .O(N__37611),
            .I(N__37608));
    Span4Mux_v I__8609 (
            .O(N__37608),
            .I(N__37605));
    Odrv4 I__8608 (
            .O(N__37605),
            .I(\b2v_inst11.func_state_RNIDUQ02Z0Z_1 ));
    InMux I__8607 (
            .O(N__37602),
            .I(N__37599));
    LocalMux I__8606 (
            .O(N__37599),
            .I(\b2v_inst11.g2_0_0Z0Z_0 ));
    InMux I__8605 (
            .O(N__37596),
            .I(N__37590));
    CascadeMux I__8604 (
            .O(N__37595),
            .I(N__37585));
    InMux I__8603 (
            .O(N__37594),
            .I(N__37579));
    InMux I__8602 (
            .O(N__37593),
            .I(N__37576));
    LocalMux I__8601 (
            .O(N__37590),
            .I(N__37573));
    InMux I__8600 (
            .O(N__37589),
            .I(N__37570));
    InMux I__8599 (
            .O(N__37588),
            .I(N__37565));
    InMux I__8598 (
            .O(N__37585),
            .I(N__37565));
    InMux I__8597 (
            .O(N__37584),
            .I(N__37560));
    InMux I__8596 (
            .O(N__37583),
            .I(N__37560));
    CascadeMux I__8595 (
            .O(N__37582),
            .I(N__37557));
    LocalMux I__8594 (
            .O(N__37579),
            .I(N__37554));
    LocalMux I__8593 (
            .O(N__37576),
            .I(N__37549));
    Span4Mux_s3_h I__8592 (
            .O(N__37573),
            .I(N__37549));
    LocalMux I__8591 (
            .O(N__37570),
            .I(N__37544));
    LocalMux I__8590 (
            .O(N__37565),
            .I(N__37544));
    LocalMux I__8589 (
            .O(N__37560),
            .I(N__37541));
    InMux I__8588 (
            .O(N__37557),
            .I(N__37537));
    Span4Mux_v I__8587 (
            .O(N__37554),
            .I(N__37534));
    Span4Mux_v I__8586 (
            .O(N__37549),
            .I(N__37527));
    Span4Mux_s2_v I__8585 (
            .O(N__37544),
            .I(N__37527));
    Span4Mux_s2_v I__8584 (
            .O(N__37541),
            .I(N__37527));
    InMux I__8583 (
            .O(N__37540),
            .I(N__37524));
    LocalMux I__8582 (
            .O(N__37537),
            .I(N__37519));
    Span4Mux_h I__8581 (
            .O(N__37534),
            .I(N__37519));
    Odrv4 I__8580 (
            .O(N__37527),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    LocalMux I__8579 (
            .O(N__37524),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    Odrv4 I__8578 (
            .O(N__37519),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    CascadeMux I__8577 (
            .O(N__37512),
            .I(N__37503));
    InMux I__8576 (
            .O(N__37511),
            .I(N__37495));
    InMux I__8575 (
            .O(N__37510),
            .I(N__37495));
    InMux I__8574 (
            .O(N__37509),
            .I(N__37492));
    InMux I__8573 (
            .O(N__37508),
            .I(N__37489));
    InMux I__8572 (
            .O(N__37507),
            .I(N__37486));
    InMux I__8571 (
            .O(N__37506),
            .I(N__37477));
    InMux I__8570 (
            .O(N__37503),
            .I(N__37477));
    InMux I__8569 (
            .O(N__37502),
            .I(N__37477));
    InMux I__8568 (
            .O(N__37501),
            .I(N__37477));
    InMux I__8567 (
            .O(N__37500),
            .I(N__37474));
    LocalMux I__8566 (
            .O(N__37495),
            .I(N__37471));
    LocalMux I__8565 (
            .O(N__37492),
            .I(N__37468));
    LocalMux I__8564 (
            .O(N__37489),
            .I(N__37465));
    LocalMux I__8563 (
            .O(N__37486),
            .I(N__37462));
    LocalMux I__8562 (
            .O(N__37477),
            .I(N__37459));
    LocalMux I__8561 (
            .O(N__37474),
            .I(N__37454));
    Span4Mux_s2_h I__8560 (
            .O(N__37471),
            .I(N__37454));
    Span4Mux_v I__8559 (
            .O(N__37468),
            .I(N__37449));
    Span4Mux_v I__8558 (
            .O(N__37465),
            .I(N__37449));
    Span4Mux_s2_h I__8557 (
            .O(N__37462),
            .I(N__37446));
    Span4Mux_s2_h I__8556 (
            .O(N__37459),
            .I(N__37441));
    Span4Mux_v I__8555 (
            .O(N__37454),
            .I(N__37441));
    Odrv4 I__8554 (
            .O(N__37449),
            .I(\b2v_inst11.N_140_N ));
    Odrv4 I__8553 (
            .O(N__37446),
            .I(\b2v_inst11.N_140_N ));
    Odrv4 I__8552 (
            .O(N__37441),
            .I(\b2v_inst11.N_140_N ));
    InMux I__8551 (
            .O(N__37434),
            .I(N__37417));
    InMux I__8550 (
            .O(N__37433),
            .I(N__37417));
    InMux I__8549 (
            .O(N__37432),
            .I(N__37417));
    InMux I__8548 (
            .O(N__37431),
            .I(N__37417));
    InMux I__8547 (
            .O(N__37430),
            .I(N__37412));
    InMux I__8546 (
            .O(N__37429),
            .I(N__37412));
    InMux I__8545 (
            .O(N__37428),
            .I(N__37409));
    InMux I__8544 (
            .O(N__37427),
            .I(N__37403));
    InMux I__8543 (
            .O(N__37426),
            .I(N__37403));
    LocalMux I__8542 (
            .O(N__37417),
            .I(N__37399));
    LocalMux I__8541 (
            .O(N__37412),
            .I(N__37394));
    LocalMux I__8540 (
            .O(N__37409),
            .I(N__37394));
    InMux I__8539 (
            .O(N__37408),
            .I(N__37391));
    LocalMux I__8538 (
            .O(N__37403),
            .I(N__37388));
    InMux I__8537 (
            .O(N__37402),
            .I(N__37385));
    Span4Mux_s0_h I__8536 (
            .O(N__37399),
            .I(N__37380));
    Span4Mux_v I__8535 (
            .O(N__37394),
            .I(N__37380));
    LocalMux I__8534 (
            .O(N__37391),
            .I(N__37375));
    Span4Mux_s3_h I__8533 (
            .O(N__37388),
            .I(N__37375));
    LocalMux I__8532 (
            .O(N__37385),
            .I(N__37372));
    Odrv4 I__8531 (
            .O(N__37380),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__8530 (
            .O(N__37375),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__8529 (
            .O(N__37372),
            .I(\b2v_inst11.N_425 ));
    CascadeMux I__8528 (
            .O(N__37365),
            .I(\b2v_inst11.N_158_N_cascade_ ));
    CascadeMux I__8527 (
            .O(N__37362),
            .I(N__37358));
    InMux I__8526 (
            .O(N__37361),
            .I(N__37351));
    InMux I__8525 (
            .O(N__37358),
            .I(N__37351));
    CascadeMux I__8524 (
            .O(N__37357),
            .I(N__37347));
    InMux I__8523 (
            .O(N__37356),
            .I(N__37337));
    LocalMux I__8522 (
            .O(N__37351),
            .I(N__37334));
    InMux I__8521 (
            .O(N__37350),
            .I(N__37327));
    InMux I__8520 (
            .O(N__37347),
            .I(N__37327));
    InMux I__8519 (
            .O(N__37346),
            .I(N__37327));
    InMux I__8518 (
            .O(N__37345),
            .I(N__37324));
    InMux I__8517 (
            .O(N__37344),
            .I(N__37320));
    InMux I__8516 (
            .O(N__37343),
            .I(N__37317));
    InMux I__8515 (
            .O(N__37342),
            .I(N__37311));
    InMux I__8514 (
            .O(N__37341),
            .I(N__37311));
    InMux I__8513 (
            .O(N__37340),
            .I(N__37308));
    LocalMux I__8512 (
            .O(N__37337),
            .I(N__37305));
    Span4Mux_v I__8511 (
            .O(N__37334),
            .I(N__37300));
    LocalMux I__8510 (
            .O(N__37327),
            .I(N__37300));
    LocalMux I__8509 (
            .O(N__37324),
            .I(N__37297));
    CascadeMux I__8508 (
            .O(N__37323),
            .I(N__37294));
    LocalMux I__8507 (
            .O(N__37320),
            .I(N__37284));
    LocalMux I__8506 (
            .O(N__37317),
            .I(N__37284));
    CascadeMux I__8505 (
            .O(N__37316),
            .I(N__37279));
    LocalMux I__8504 (
            .O(N__37311),
            .I(N__37272));
    LocalMux I__8503 (
            .O(N__37308),
            .I(N__37272));
    Span4Mux_v I__8502 (
            .O(N__37305),
            .I(N__37265));
    Span4Mux_v I__8501 (
            .O(N__37300),
            .I(N__37265));
    Span4Mux_h I__8500 (
            .O(N__37297),
            .I(N__37265));
    InMux I__8499 (
            .O(N__37294),
            .I(N__37262));
    InMux I__8498 (
            .O(N__37293),
            .I(N__37257));
    InMux I__8497 (
            .O(N__37292),
            .I(N__37257));
    InMux I__8496 (
            .O(N__37291),
            .I(N__37254));
    InMux I__8495 (
            .O(N__37290),
            .I(N__37249));
    InMux I__8494 (
            .O(N__37289),
            .I(N__37249));
    Span4Mux_h I__8493 (
            .O(N__37284),
            .I(N__37246));
    InMux I__8492 (
            .O(N__37283),
            .I(N__37241));
    InMux I__8491 (
            .O(N__37282),
            .I(N__37241));
    InMux I__8490 (
            .O(N__37279),
            .I(N__37234));
    InMux I__8489 (
            .O(N__37278),
            .I(N__37234));
    InMux I__8488 (
            .O(N__37277),
            .I(N__37234));
    Span4Mux_h I__8487 (
            .O(N__37272),
            .I(N__37229));
    Span4Mux_h I__8486 (
            .O(N__37265),
            .I(N__37229));
    LocalMux I__8485 (
            .O(N__37262),
            .I(N__37224));
    LocalMux I__8484 (
            .O(N__37257),
            .I(N__37224));
    LocalMux I__8483 (
            .O(N__37254),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    LocalMux I__8482 (
            .O(N__37249),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv4 I__8481 (
            .O(N__37246),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    LocalMux I__8480 (
            .O(N__37241),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    LocalMux I__8479 (
            .O(N__37234),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv4 I__8478 (
            .O(N__37229),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv12 I__8477 (
            .O(N__37224),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    InMux I__8476 (
            .O(N__37209),
            .I(N__37206));
    LocalMux I__8475 (
            .O(N__37206),
            .I(\b2v_inst11.dutycycle_en_12 ));
    InMux I__8474 (
            .O(N__37203),
            .I(N__37197));
    InMux I__8473 (
            .O(N__37202),
            .I(N__37197));
    LocalMux I__8472 (
            .O(N__37197),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3AZ0Z64 ));
    CascadeMux I__8471 (
            .O(N__37194),
            .I(\b2v_inst11.dutycycle_en_12_cascade_ ));
    CascadeMux I__8470 (
            .O(N__37191),
            .I(N__37187));
    InMux I__8469 (
            .O(N__37190),
            .I(N__37182));
    InMux I__8468 (
            .O(N__37187),
            .I(N__37182));
    LocalMux I__8467 (
            .O(N__37182),
            .I(\b2v_inst11.dutycycleZ0Z_15 ));
    CascadeMux I__8466 (
            .O(N__37179),
            .I(N__37175));
    InMux I__8465 (
            .O(N__37178),
            .I(N__37172));
    InMux I__8464 (
            .O(N__37175),
            .I(N__37169));
    LocalMux I__8463 (
            .O(N__37172),
            .I(N__37165));
    LocalMux I__8462 (
            .O(N__37169),
            .I(N__37162));
    InMux I__8461 (
            .O(N__37168),
            .I(N__37159));
    Span12Mux_s8_v I__8460 (
            .O(N__37165),
            .I(N__37154));
    Span12Mux_s0_h I__8459 (
            .O(N__37162),
            .I(N__37154));
    LocalMux I__8458 (
            .O(N__37159),
            .I(\b2v_inst11.N_326_N ));
    Odrv12 I__8457 (
            .O(N__37154),
            .I(\b2v_inst11.N_326_N ));
    ClkMux I__8456 (
            .O(N__37149),
            .I(N__37145));
    ClkMux I__8455 (
            .O(N__37148),
            .I(N__37136));
    LocalMux I__8454 (
            .O(N__37145),
            .I(N__37131));
    ClkMux I__8453 (
            .O(N__37144),
            .I(N__37128));
    ClkMux I__8452 (
            .O(N__37143),
            .I(N__37122));
    ClkMux I__8451 (
            .O(N__37142),
            .I(N__37119));
    ClkMux I__8450 (
            .O(N__37141),
            .I(N__37116));
    ClkMux I__8449 (
            .O(N__37140),
            .I(N__37113));
    ClkMux I__8448 (
            .O(N__37139),
            .I(N__37110));
    LocalMux I__8447 (
            .O(N__37136),
            .I(N__37105));
    ClkMux I__8446 (
            .O(N__37135),
            .I(N__37102));
    ClkMux I__8445 (
            .O(N__37134),
            .I(N__37096));
    Span4Mux_s1_h I__8444 (
            .O(N__37131),
            .I(N__37092));
    LocalMux I__8443 (
            .O(N__37128),
            .I(N__37089));
    ClkMux I__8442 (
            .O(N__37127),
            .I(N__37082));
    ClkMux I__8441 (
            .O(N__37126),
            .I(N__37079));
    ClkMux I__8440 (
            .O(N__37125),
            .I(N__37076));
    LocalMux I__8439 (
            .O(N__37122),
            .I(N__37073));
    LocalMux I__8438 (
            .O(N__37119),
            .I(N__37064));
    LocalMux I__8437 (
            .O(N__37116),
            .I(N__37055));
    LocalMux I__8436 (
            .O(N__37113),
            .I(N__37055));
    LocalMux I__8435 (
            .O(N__37110),
            .I(N__37055));
    ClkMux I__8434 (
            .O(N__37109),
            .I(N__37052));
    ClkMux I__8433 (
            .O(N__37108),
            .I(N__37049));
    Span4Mux_v I__8432 (
            .O(N__37105),
            .I(N__37044));
    LocalMux I__8431 (
            .O(N__37102),
            .I(N__37044));
    ClkMux I__8430 (
            .O(N__37101),
            .I(N__37041));
    ClkMux I__8429 (
            .O(N__37100),
            .I(N__37038));
    ClkMux I__8428 (
            .O(N__37099),
            .I(N__37035));
    LocalMux I__8427 (
            .O(N__37096),
            .I(N__37031));
    ClkMux I__8426 (
            .O(N__37095),
            .I(N__37028));
    Span4Mux_v I__8425 (
            .O(N__37092),
            .I(N__37022));
    Span4Mux_s1_h I__8424 (
            .O(N__37089),
            .I(N__37022));
    ClkMux I__8423 (
            .O(N__37088),
            .I(N__37019));
    ClkMux I__8422 (
            .O(N__37087),
            .I(N__37015));
    ClkMux I__8421 (
            .O(N__37086),
            .I(N__37011));
    ClkMux I__8420 (
            .O(N__37085),
            .I(N__37008));
    LocalMux I__8419 (
            .O(N__37082),
            .I(N__37003));
    LocalMux I__8418 (
            .O(N__37079),
            .I(N__36998));
    LocalMux I__8417 (
            .O(N__37076),
            .I(N__36993));
    Span4Mux_v I__8416 (
            .O(N__37073),
            .I(N__36990));
    ClkMux I__8415 (
            .O(N__37072),
            .I(N__36987));
    ClkMux I__8414 (
            .O(N__37071),
            .I(N__36984));
    ClkMux I__8413 (
            .O(N__37070),
            .I(N__36981));
    ClkMux I__8412 (
            .O(N__37069),
            .I(N__36977));
    ClkMux I__8411 (
            .O(N__37068),
            .I(N__36974));
    ClkMux I__8410 (
            .O(N__37067),
            .I(N__36970));
    Span4Mux_s2_h I__8409 (
            .O(N__37064),
            .I(N__36962));
    ClkMux I__8408 (
            .O(N__37063),
            .I(N__36959));
    ClkMux I__8407 (
            .O(N__37062),
            .I(N__36956));
    Span4Mux_v I__8406 (
            .O(N__37055),
            .I(N__36948));
    LocalMux I__8405 (
            .O(N__37052),
            .I(N__36948));
    LocalMux I__8404 (
            .O(N__37049),
            .I(N__36948));
    Span4Mux_v I__8403 (
            .O(N__37044),
            .I(N__36943));
    LocalMux I__8402 (
            .O(N__37041),
            .I(N__36943));
    LocalMux I__8401 (
            .O(N__37038),
            .I(N__36939));
    LocalMux I__8400 (
            .O(N__37035),
            .I(N__36936));
    ClkMux I__8399 (
            .O(N__37034),
            .I(N__36933));
    Span4Mux_v I__8398 (
            .O(N__37031),
            .I(N__36928));
    LocalMux I__8397 (
            .O(N__37028),
            .I(N__36928));
    ClkMux I__8396 (
            .O(N__37027),
            .I(N__36925));
    Span4Mux_h I__8395 (
            .O(N__37022),
            .I(N__36922));
    LocalMux I__8394 (
            .O(N__37019),
            .I(N__36919));
    ClkMux I__8393 (
            .O(N__37018),
            .I(N__36916));
    LocalMux I__8392 (
            .O(N__37015),
            .I(N__36913));
    ClkMux I__8391 (
            .O(N__37014),
            .I(N__36910));
    LocalMux I__8390 (
            .O(N__37011),
            .I(N__36906));
    LocalMux I__8389 (
            .O(N__37008),
            .I(N__36903));
    ClkMux I__8388 (
            .O(N__37007),
            .I(N__36900));
    ClkMux I__8387 (
            .O(N__37006),
            .I(N__36895));
    Span4Mux_s1_h I__8386 (
            .O(N__37003),
            .I(N__36892));
    ClkMux I__8385 (
            .O(N__37002),
            .I(N__36886));
    ClkMux I__8384 (
            .O(N__37001),
            .I(N__36883));
    Span4Mux_v I__8383 (
            .O(N__36998),
            .I(N__36880));
    ClkMux I__8382 (
            .O(N__36997),
            .I(N__36877));
    ClkMux I__8381 (
            .O(N__36996),
            .I(N__36874));
    Span4Mux_h I__8380 (
            .O(N__36993),
            .I(N__36863));
    Span4Mux_h I__8379 (
            .O(N__36990),
            .I(N__36863));
    LocalMux I__8378 (
            .O(N__36987),
            .I(N__36863));
    LocalMux I__8377 (
            .O(N__36984),
            .I(N__36863));
    LocalMux I__8376 (
            .O(N__36981),
            .I(N__36858));
    ClkMux I__8375 (
            .O(N__36980),
            .I(N__36855));
    LocalMux I__8374 (
            .O(N__36977),
            .I(N__36850));
    LocalMux I__8373 (
            .O(N__36974),
            .I(N__36850));
    ClkMux I__8372 (
            .O(N__36973),
            .I(N__36847));
    LocalMux I__8371 (
            .O(N__36970),
            .I(N__36844));
    ClkMux I__8370 (
            .O(N__36969),
            .I(N__36841));
    ClkMux I__8369 (
            .O(N__36968),
            .I(N__36837));
    ClkMux I__8368 (
            .O(N__36967),
            .I(N__36831));
    ClkMux I__8367 (
            .O(N__36966),
            .I(N__36827));
    ClkMux I__8366 (
            .O(N__36965),
            .I(N__36824));
    Span4Mux_h I__8365 (
            .O(N__36962),
            .I(N__36817));
    LocalMux I__8364 (
            .O(N__36959),
            .I(N__36817));
    LocalMux I__8363 (
            .O(N__36956),
            .I(N__36814));
    ClkMux I__8362 (
            .O(N__36955),
            .I(N__36811));
    Span4Mux_v I__8361 (
            .O(N__36948),
            .I(N__36805));
    Span4Mux_v I__8360 (
            .O(N__36943),
            .I(N__36805));
    ClkMux I__8359 (
            .O(N__36942),
            .I(N__36802));
    Span4Mux_s1_h I__8358 (
            .O(N__36939),
            .I(N__36793));
    Span4Mux_v I__8357 (
            .O(N__36936),
            .I(N__36793));
    LocalMux I__8356 (
            .O(N__36933),
            .I(N__36793));
    Span4Mux_v I__8355 (
            .O(N__36928),
            .I(N__36788));
    LocalMux I__8354 (
            .O(N__36925),
            .I(N__36788));
    Span4Mux_v I__8353 (
            .O(N__36922),
            .I(N__36781));
    Span4Mux_v I__8352 (
            .O(N__36919),
            .I(N__36781));
    LocalMux I__8351 (
            .O(N__36916),
            .I(N__36781));
    Span4Mux_v I__8350 (
            .O(N__36913),
            .I(N__36776));
    LocalMux I__8349 (
            .O(N__36910),
            .I(N__36776));
    ClkMux I__8348 (
            .O(N__36909),
            .I(N__36771));
    Span4Mux_s1_h I__8347 (
            .O(N__36906),
            .I(N__36768));
    Span4Mux_s1_h I__8346 (
            .O(N__36903),
            .I(N__36765));
    LocalMux I__8345 (
            .O(N__36900),
            .I(N__36762));
    ClkMux I__8344 (
            .O(N__36899),
            .I(N__36759));
    ClkMux I__8343 (
            .O(N__36898),
            .I(N__36756));
    LocalMux I__8342 (
            .O(N__36895),
            .I(N__36752));
    Span4Mux_h I__8341 (
            .O(N__36892),
            .I(N__36749));
    ClkMux I__8340 (
            .O(N__36891),
            .I(N__36746));
    ClkMux I__8339 (
            .O(N__36890),
            .I(N__36741));
    ClkMux I__8338 (
            .O(N__36889),
            .I(N__36738));
    LocalMux I__8337 (
            .O(N__36886),
            .I(N__36733));
    LocalMux I__8336 (
            .O(N__36883),
            .I(N__36733));
    Span4Mux_h I__8335 (
            .O(N__36880),
            .I(N__36726));
    LocalMux I__8334 (
            .O(N__36877),
            .I(N__36726));
    LocalMux I__8333 (
            .O(N__36874),
            .I(N__36726));
    ClkMux I__8332 (
            .O(N__36873),
            .I(N__36723));
    ClkMux I__8331 (
            .O(N__36872),
            .I(N__36720));
    Span4Mux_v I__8330 (
            .O(N__36863),
            .I(N__36716));
    ClkMux I__8329 (
            .O(N__36862),
            .I(N__36713));
    ClkMux I__8328 (
            .O(N__36861),
            .I(N__36710));
    Span4Mux_s3_h I__8327 (
            .O(N__36858),
            .I(N__36704));
    LocalMux I__8326 (
            .O(N__36855),
            .I(N__36704));
    Span4Mux_v I__8325 (
            .O(N__36850),
            .I(N__36695));
    LocalMux I__8324 (
            .O(N__36847),
            .I(N__36695));
    Span4Mux_s3_h I__8323 (
            .O(N__36844),
            .I(N__36695));
    LocalMux I__8322 (
            .O(N__36841),
            .I(N__36695));
    ClkMux I__8321 (
            .O(N__36840),
            .I(N__36692));
    LocalMux I__8320 (
            .O(N__36837),
            .I(N__36689));
    ClkMux I__8319 (
            .O(N__36836),
            .I(N__36686));
    ClkMux I__8318 (
            .O(N__36835),
            .I(N__36683));
    ClkMux I__8317 (
            .O(N__36834),
            .I(N__36680));
    LocalMux I__8316 (
            .O(N__36831),
            .I(N__36677));
    ClkMux I__8315 (
            .O(N__36830),
            .I(N__36674));
    LocalMux I__8314 (
            .O(N__36827),
            .I(N__36668));
    LocalMux I__8313 (
            .O(N__36824),
            .I(N__36668));
    ClkMux I__8312 (
            .O(N__36823),
            .I(N__36665));
    ClkMux I__8311 (
            .O(N__36822),
            .I(N__36662));
    Span4Mux_v I__8310 (
            .O(N__36817),
            .I(N__36655));
    Span4Mux_h I__8309 (
            .O(N__36814),
            .I(N__36655));
    LocalMux I__8308 (
            .O(N__36811),
            .I(N__36655));
    ClkMux I__8307 (
            .O(N__36810),
            .I(N__36652));
    IoSpan4Mux I__8306 (
            .O(N__36805),
            .I(N__36647));
    LocalMux I__8305 (
            .O(N__36802),
            .I(N__36647));
    ClkMux I__8304 (
            .O(N__36801),
            .I(N__36644));
    ClkMux I__8303 (
            .O(N__36800),
            .I(N__36641));
    Span4Mux_v I__8302 (
            .O(N__36793),
            .I(N__36636));
    Span4Mux_v I__8301 (
            .O(N__36788),
            .I(N__36633));
    Span4Mux_v I__8300 (
            .O(N__36781),
            .I(N__36628));
    Span4Mux_h I__8299 (
            .O(N__36776),
            .I(N__36628));
    ClkMux I__8298 (
            .O(N__36775),
            .I(N__36625));
    ClkMux I__8297 (
            .O(N__36774),
            .I(N__36622));
    LocalMux I__8296 (
            .O(N__36771),
            .I(N__36619));
    Span4Mux_h I__8295 (
            .O(N__36768),
            .I(N__36612));
    Span4Mux_h I__8294 (
            .O(N__36765),
            .I(N__36612));
    Span4Mux_h I__8293 (
            .O(N__36762),
            .I(N__36612));
    LocalMux I__8292 (
            .O(N__36759),
            .I(N__36608));
    LocalMux I__8291 (
            .O(N__36756),
            .I(N__36605));
    ClkMux I__8290 (
            .O(N__36755),
            .I(N__36602));
    Span4Mux_s1_h I__8289 (
            .O(N__36752),
            .I(N__36599));
    Span4Mux_v I__8288 (
            .O(N__36749),
            .I(N__36594));
    LocalMux I__8287 (
            .O(N__36746),
            .I(N__36594));
    ClkMux I__8286 (
            .O(N__36745),
            .I(N__36591));
    ClkMux I__8285 (
            .O(N__36744),
            .I(N__36588));
    LocalMux I__8284 (
            .O(N__36741),
            .I(N__36585));
    LocalMux I__8283 (
            .O(N__36738),
            .I(N__36582));
    Span4Mux_v I__8282 (
            .O(N__36733),
            .I(N__36573));
    Span4Mux_v I__8281 (
            .O(N__36726),
            .I(N__36573));
    LocalMux I__8280 (
            .O(N__36723),
            .I(N__36573));
    LocalMux I__8279 (
            .O(N__36720),
            .I(N__36573));
    ClkMux I__8278 (
            .O(N__36719),
            .I(N__36570));
    Span4Mux_h I__8277 (
            .O(N__36716),
            .I(N__36565));
    LocalMux I__8276 (
            .O(N__36713),
            .I(N__36565));
    LocalMux I__8275 (
            .O(N__36710),
            .I(N__36562));
    ClkMux I__8274 (
            .O(N__36709),
            .I(N__36559));
    Span4Mux_v I__8273 (
            .O(N__36704),
            .I(N__36544));
    Span4Mux_v I__8272 (
            .O(N__36695),
            .I(N__36544));
    LocalMux I__8271 (
            .O(N__36692),
            .I(N__36544));
    Span4Mux_s3_h I__8270 (
            .O(N__36689),
            .I(N__36544));
    LocalMux I__8269 (
            .O(N__36686),
            .I(N__36544));
    LocalMux I__8268 (
            .O(N__36683),
            .I(N__36544));
    LocalMux I__8267 (
            .O(N__36680),
            .I(N__36544));
    Span4Mux_s2_h I__8266 (
            .O(N__36677),
            .I(N__36541));
    LocalMux I__8265 (
            .O(N__36674),
            .I(N__36538));
    ClkMux I__8264 (
            .O(N__36673),
            .I(N__36535));
    Span4Mux_h I__8263 (
            .O(N__36668),
            .I(N__36528));
    LocalMux I__8262 (
            .O(N__36665),
            .I(N__36528));
    LocalMux I__8261 (
            .O(N__36662),
            .I(N__36528));
    Span4Mux_v I__8260 (
            .O(N__36655),
            .I(N__36523));
    LocalMux I__8259 (
            .O(N__36652),
            .I(N__36523));
    Span4Mux_s0_v I__8258 (
            .O(N__36647),
            .I(N__36516));
    LocalMux I__8257 (
            .O(N__36644),
            .I(N__36516));
    LocalMux I__8256 (
            .O(N__36641),
            .I(N__36516));
    ClkMux I__8255 (
            .O(N__36640),
            .I(N__36513));
    ClkMux I__8254 (
            .O(N__36639),
            .I(N__36509));
    Span4Mux_h I__8253 (
            .O(N__36636),
            .I(N__36498));
    Span4Mux_h I__8252 (
            .O(N__36633),
            .I(N__36498));
    Span4Mux_h I__8251 (
            .O(N__36628),
            .I(N__36498));
    LocalMux I__8250 (
            .O(N__36625),
            .I(N__36498));
    LocalMux I__8249 (
            .O(N__36622),
            .I(N__36498));
    Span4Mux_v I__8248 (
            .O(N__36619),
            .I(N__36493));
    Span4Mux_v I__8247 (
            .O(N__36612),
            .I(N__36493));
    ClkMux I__8246 (
            .O(N__36611),
            .I(N__36490));
    Span4Mux_s1_h I__8245 (
            .O(N__36608),
            .I(N__36487));
    Span4Mux_s2_h I__8244 (
            .O(N__36605),
            .I(N__36482));
    LocalMux I__8243 (
            .O(N__36602),
            .I(N__36482));
    Span4Mux_h I__8242 (
            .O(N__36599),
            .I(N__36473));
    Span4Mux_v I__8241 (
            .O(N__36594),
            .I(N__36473));
    LocalMux I__8240 (
            .O(N__36591),
            .I(N__36473));
    LocalMux I__8239 (
            .O(N__36588),
            .I(N__36473));
    IoSpan4Mux I__8238 (
            .O(N__36585),
            .I(N__36470));
    Span4Mux_h I__8237 (
            .O(N__36582),
            .I(N__36463));
    Span4Mux_v I__8236 (
            .O(N__36573),
            .I(N__36463));
    LocalMux I__8235 (
            .O(N__36570),
            .I(N__36463));
    Span4Mux_v I__8234 (
            .O(N__36565),
            .I(N__36454));
    Span4Mux_s3_h I__8233 (
            .O(N__36562),
            .I(N__36454));
    LocalMux I__8232 (
            .O(N__36559),
            .I(N__36454));
    Span4Mux_v I__8231 (
            .O(N__36544),
            .I(N__36454));
    Span4Mux_v I__8230 (
            .O(N__36541),
            .I(N__36447));
    Span4Mux_s2_h I__8229 (
            .O(N__36538),
            .I(N__36447));
    LocalMux I__8228 (
            .O(N__36535),
            .I(N__36447));
    Span4Mux_v I__8227 (
            .O(N__36528),
            .I(N__36438));
    Span4Mux_v I__8226 (
            .O(N__36523),
            .I(N__36438));
    Span4Mux_h I__8225 (
            .O(N__36516),
            .I(N__36438));
    LocalMux I__8224 (
            .O(N__36513),
            .I(N__36438));
    ClkMux I__8223 (
            .O(N__36512),
            .I(N__36433));
    LocalMux I__8222 (
            .O(N__36509),
            .I(N__36428));
    Span4Mux_s2_v I__8221 (
            .O(N__36498),
            .I(N__36428));
    Span4Mux_v I__8220 (
            .O(N__36493),
            .I(N__36424));
    LocalMux I__8219 (
            .O(N__36490),
            .I(N__36421));
    Span4Mux_h I__8218 (
            .O(N__36487),
            .I(N__36414));
    Span4Mux_h I__8217 (
            .O(N__36482),
            .I(N__36414));
    Span4Mux_v I__8216 (
            .O(N__36473),
            .I(N__36414));
    IoSpan4Mux I__8215 (
            .O(N__36470),
            .I(N__36407));
    IoSpan4Mux I__8214 (
            .O(N__36463),
            .I(N__36407));
    IoSpan4Mux I__8213 (
            .O(N__36454),
            .I(N__36407));
    IoSpan4Mux I__8212 (
            .O(N__36447),
            .I(N__36402));
    IoSpan4Mux I__8211 (
            .O(N__36438),
            .I(N__36402));
    ClkMux I__8210 (
            .O(N__36437),
            .I(N__36399));
    ClkMux I__8209 (
            .O(N__36436),
            .I(N__36396));
    LocalMux I__8208 (
            .O(N__36433),
            .I(N__36391));
    Span4Mux_v I__8207 (
            .O(N__36428),
            .I(N__36391));
    ClkMux I__8206 (
            .O(N__36427),
            .I(N__36388));
    Odrv4 I__8205 (
            .O(N__36424),
            .I(fpga_osc));
    Odrv12 I__8204 (
            .O(N__36421),
            .I(fpga_osc));
    Odrv4 I__8203 (
            .O(N__36414),
            .I(fpga_osc));
    Odrv4 I__8202 (
            .O(N__36407),
            .I(fpga_osc));
    Odrv4 I__8201 (
            .O(N__36402),
            .I(fpga_osc));
    LocalMux I__8200 (
            .O(N__36399),
            .I(fpga_osc));
    LocalMux I__8199 (
            .O(N__36396),
            .I(fpga_osc));
    Odrv4 I__8198 (
            .O(N__36391),
            .I(fpga_osc));
    LocalMux I__8197 (
            .O(N__36388),
            .I(fpga_osc));
    SRMux I__8196 (
            .O(N__36369),
            .I(N__36363));
    SRMux I__8195 (
            .O(N__36368),
            .I(N__36358));
    SRMux I__8194 (
            .O(N__36367),
            .I(N__36355));
    SRMux I__8193 (
            .O(N__36366),
            .I(N__36352));
    LocalMux I__8192 (
            .O(N__36363),
            .I(N__36349));
    SRMux I__8191 (
            .O(N__36362),
            .I(N__36345));
    SRMux I__8190 (
            .O(N__36361),
            .I(N__36342));
    LocalMux I__8189 (
            .O(N__36358),
            .I(N__36338));
    LocalMux I__8188 (
            .O(N__36355),
            .I(N__36333));
    LocalMux I__8187 (
            .O(N__36352),
            .I(N__36333));
    Span4Mux_s0_h I__8186 (
            .O(N__36349),
            .I(N__36330));
    SRMux I__8185 (
            .O(N__36348),
            .I(N__36327));
    LocalMux I__8184 (
            .O(N__36345),
            .I(N__36321));
    LocalMux I__8183 (
            .O(N__36342),
            .I(N__36318));
    SRMux I__8182 (
            .O(N__36341),
            .I(N__36315));
    Span4Mux_v I__8181 (
            .O(N__36338),
            .I(N__36310));
    Span4Mux_v I__8180 (
            .O(N__36333),
            .I(N__36310));
    Span4Mux_s2_v I__8179 (
            .O(N__36330),
            .I(N__36305));
    LocalMux I__8178 (
            .O(N__36327),
            .I(N__36305));
    SRMux I__8177 (
            .O(N__36326),
            .I(N__36302));
    SRMux I__8176 (
            .O(N__36325),
            .I(N__36299));
    SRMux I__8175 (
            .O(N__36324),
            .I(N__36296));
    Span4Mux_s3_h I__8174 (
            .O(N__36321),
            .I(N__36291));
    Span4Mux_s3_h I__8173 (
            .O(N__36318),
            .I(N__36291));
    LocalMux I__8172 (
            .O(N__36315),
            .I(N__36288));
    Span4Mux_h I__8171 (
            .O(N__36310),
            .I(N__36285));
    Span4Mux_v I__8170 (
            .O(N__36305),
            .I(N__36282));
    LocalMux I__8169 (
            .O(N__36302),
            .I(N__36279));
    LocalMux I__8168 (
            .O(N__36299),
            .I(N__36274));
    LocalMux I__8167 (
            .O(N__36296),
            .I(N__36274));
    Span4Mux_v I__8166 (
            .O(N__36291),
            .I(N__36271));
    Span4Mux_v I__8165 (
            .O(N__36288),
            .I(N__36266));
    Span4Mux_h I__8164 (
            .O(N__36285),
            .I(N__36266));
    Span4Mux_v I__8163 (
            .O(N__36282),
            .I(N__36263));
    Span4Mux_v I__8162 (
            .O(N__36279),
            .I(N__36256));
    Span4Mux_v I__8161 (
            .O(N__36274),
            .I(N__36256));
    Span4Mux_s3_h I__8160 (
            .O(N__36271),
            .I(N__36256));
    Span4Mux_v I__8159 (
            .O(N__36266),
            .I(N__36253));
    Odrv4 I__8158 (
            .O(N__36263),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv4 I__8157 (
            .O(N__36256),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv4 I__8156 (
            .O(N__36253),
            .I(\b2v_inst11.N_224_iZ0 ));
    InMux I__8155 (
            .O(N__36246),
            .I(N__36243));
    LocalMux I__8154 (
            .O(N__36243),
            .I(N__36240));
    Span4Mux_s1_h I__8153 (
            .O(N__36240),
            .I(N__36237));
    Span4Mux_v I__8152 (
            .O(N__36237),
            .I(N__36234));
    Odrv4 I__8151 (
            .O(N__36234),
            .I(\b2v_inst11.un1_dutycycle_94_s1_8 ));
    CascadeMux I__8150 (
            .O(N__36231),
            .I(N__36217));
    CascadeMux I__8149 (
            .O(N__36230),
            .I(N__36212));
    InMux I__8148 (
            .O(N__36229),
            .I(N__36200));
    InMux I__8147 (
            .O(N__36228),
            .I(N__36191));
    InMux I__8146 (
            .O(N__36227),
            .I(N__36191));
    InMux I__8145 (
            .O(N__36226),
            .I(N__36191));
    InMux I__8144 (
            .O(N__36225),
            .I(N__36191));
    InMux I__8143 (
            .O(N__36224),
            .I(N__36188));
    InMux I__8142 (
            .O(N__36223),
            .I(N__36185));
    InMux I__8141 (
            .O(N__36222),
            .I(N__36182));
    CascadeMux I__8140 (
            .O(N__36221),
            .I(N__36179));
    InMux I__8139 (
            .O(N__36220),
            .I(N__36170));
    InMux I__8138 (
            .O(N__36217),
            .I(N__36163));
    InMux I__8137 (
            .O(N__36216),
            .I(N__36163));
    InMux I__8136 (
            .O(N__36215),
            .I(N__36163));
    InMux I__8135 (
            .O(N__36212),
            .I(N__36158));
    InMux I__8134 (
            .O(N__36211),
            .I(N__36158));
    InMux I__8133 (
            .O(N__36210),
            .I(N__36151));
    InMux I__8132 (
            .O(N__36209),
            .I(N__36151));
    InMux I__8131 (
            .O(N__36208),
            .I(N__36151));
    InMux I__8130 (
            .O(N__36207),
            .I(N__36140));
    InMux I__8129 (
            .O(N__36206),
            .I(N__36140));
    InMux I__8128 (
            .O(N__36205),
            .I(N__36140));
    InMux I__8127 (
            .O(N__36204),
            .I(N__36140));
    InMux I__8126 (
            .O(N__36203),
            .I(N__36140));
    LocalMux I__8125 (
            .O(N__36200),
            .I(N__36129));
    LocalMux I__8124 (
            .O(N__36191),
            .I(N__36129));
    LocalMux I__8123 (
            .O(N__36188),
            .I(N__36129));
    LocalMux I__8122 (
            .O(N__36185),
            .I(N__36129));
    LocalMux I__8121 (
            .O(N__36182),
            .I(N__36129));
    InMux I__8120 (
            .O(N__36179),
            .I(N__36126));
    InMux I__8119 (
            .O(N__36178),
            .I(N__36117));
    InMux I__8118 (
            .O(N__36177),
            .I(N__36117));
    InMux I__8117 (
            .O(N__36176),
            .I(N__36117));
    InMux I__8116 (
            .O(N__36175),
            .I(N__36117));
    InMux I__8115 (
            .O(N__36174),
            .I(N__36114));
    InMux I__8114 (
            .O(N__36173),
            .I(N__36111));
    LocalMux I__8113 (
            .O(N__36170),
            .I(N__36096));
    LocalMux I__8112 (
            .O(N__36163),
            .I(N__36096));
    LocalMux I__8111 (
            .O(N__36158),
            .I(N__36096));
    LocalMux I__8110 (
            .O(N__36151),
            .I(N__36096));
    LocalMux I__8109 (
            .O(N__36140),
            .I(N__36096));
    Span4Mux_v I__8108 (
            .O(N__36129),
            .I(N__36096));
    LocalMux I__8107 (
            .O(N__36126),
            .I(N__36096));
    LocalMux I__8106 (
            .O(N__36117),
            .I(N__36091));
    LocalMux I__8105 (
            .O(N__36114),
            .I(N__36091));
    LocalMux I__8104 (
            .O(N__36111),
            .I(N__36088));
    Span4Mux_v I__8103 (
            .O(N__36096),
            .I(N__36085));
    Odrv4 I__8102 (
            .O(N__36091),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    Odrv12 I__8101 (
            .O(N__36088),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    Odrv4 I__8100 (
            .O(N__36085),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ));
    CascadeMux I__8099 (
            .O(N__36078),
            .I(N__36075));
    InMux I__8098 (
            .O(N__36075),
            .I(N__36072));
    LocalMux I__8097 (
            .O(N__36072),
            .I(\b2v_inst11.un1_dutycycle_94_s0_8 ));
    CascadeMux I__8096 (
            .O(N__36069),
            .I(N__36065));
    CascadeMux I__8095 (
            .O(N__36068),
            .I(N__36062));
    InMux I__8094 (
            .O(N__36065),
            .I(N__36054));
    InMux I__8093 (
            .O(N__36062),
            .I(N__36051));
    CascadeMux I__8092 (
            .O(N__36061),
            .I(N__36046));
    CascadeMux I__8091 (
            .O(N__36060),
            .I(N__36043));
    CascadeMux I__8090 (
            .O(N__36059),
            .I(N__36038));
    InMux I__8089 (
            .O(N__36058),
            .I(N__36032));
    InMux I__8088 (
            .O(N__36057),
            .I(N__36032));
    LocalMux I__8087 (
            .O(N__36054),
            .I(N__36027));
    LocalMux I__8086 (
            .O(N__36051),
            .I(N__36027));
    InMux I__8085 (
            .O(N__36050),
            .I(N__36024));
    InMux I__8084 (
            .O(N__36049),
            .I(N__36021));
    InMux I__8083 (
            .O(N__36046),
            .I(N__36016));
    InMux I__8082 (
            .O(N__36043),
            .I(N__36013));
    CascadeMux I__8081 (
            .O(N__36042),
            .I(N__36006));
    CascadeMux I__8080 (
            .O(N__36041),
            .I(N__36001));
    InMux I__8079 (
            .O(N__36038),
            .I(N__35998));
    InMux I__8078 (
            .O(N__36037),
            .I(N__35995));
    LocalMux I__8077 (
            .O(N__36032),
            .I(N__35992));
    Span4Mux_s3_v I__8076 (
            .O(N__36027),
            .I(N__35985));
    LocalMux I__8075 (
            .O(N__36024),
            .I(N__35985));
    LocalMux I__8074 (
            .O(N__36021),
            .I(N__35985));
    InMux I__8073 (
            .O(N__36020),
            .I(N__35980));
    InMux I__8072 (
            .O(N__36019),
            .I(N__35980));
    LocalMux I__8071 (
            .O(N__36016),
            .I(N__35975));
    LocalMux I__8070 (
            .O(N__36013),
            .I(N__35975));
    InMux I__8069 (
            .O(N__36012),
            .I(N__35970));
    InMux I__8068 (
            .O(N__36011),
            .I(N__35970));
    InMux I__8067 (
            .O(N__36010),
            .I(N__35967));
    InMux I__8066 (
            .O(N__36009),
            .I(N__35964));
    InMux I__8065 (
            .O(N__36006),
            .I(N__35959));
    InMux I__8064 (
            .O(N__36005),
            .I(N__35959));
    InMux I__8063 (
            .O(N__36004),
            .I(N__35956));
    InMux I__8062 (
            .O(N__36001),
            .I(N__35953));
    LocalMux I__8061 (
            .O(N__35998),
            .I(N__35948));
    LocalMux I__8060 (
            .O(N__35995),
            .I(N__35948));
    Span4Mux_v I__8059 (
            .O(N__35992),
            .I(N__35941));
    Span4Mux_v I__8058 (
            .O(N__35985),
            .I(N__35941));
    LocalMux I__8057 (
            .O(N__35980),
            .I(N__35932));
    Span4Mux_s3_v I__8056 (
            .O(N__35975),
            .I(N__35932));
    LocalMux I__8055 (
            .O(N__35970),
            .I(N__35932));
    LocalMux I__8054 (
            .O(N__35967),
            .I(N__35932));
    LocalMux I__8053 (
            .O(N__35964),
            .I(N__35921));
    LocalMux I__8052 (
            .O(N__35959),
            .I(N__35921));
    LocalMux I__8051 (
            .O(N__35956),
            .I(N__35921));
    LocalMux I__8050 (
            .O(N__35953),
            .I(N__35921));
    Span4Mux_s3_v I__8049 (
            .O(N__35948),
            .I(N__35921));
    InMux I__8048 (
            .O(N__35947),
            .I(N__35914));
    InMux I__8047 (
            .O(N__35946),
            .I(N__35914));
    Span4Mux_s0_h I__8046 (
            .O(N__35941),
            .I(N__35907));
    Span4Mux_v I__8045 (
            .O(N__35932),
            .I(N__35907));
    Span4Mux_v I__8044 (
            .O(N__35921),
            .I(N__35907));
    InMux I__8043 (
            .O(N__35920),
            .I(N__35902));
    InMux I__8042 (
            .O(N__35919),
            .I(N__35902));
    LocalMux I__8041 (
            .O(N__35914),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    Odrv4 I__8040 (
            .O(N__35907),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    LocalMux I__8039 (
            .O(N__35902),
            .I(\b2v_inst11.dutycycleZ1Z_5 ));
    InMux I__8038 (
            .O(N__35895),
            .I(N__35892));
    LocalMux I__8037 (
            .O(N__35892),
            .I(\b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1 ));
    InMux I__8036 (
            .O(N__35889),
            .I(N__35883));
    InMux I__8035 (
            .O(N__35888),
            .I(N__35883));
    LocalMux I__8034 (
            .O(N__35883),
            .I(\b2v_inst11.dutycycleZ1Z_8 ));
    InMux I__8033 (
            .O(N__35880),
            .I(N__35874));
    InMux I__8032 (
            .O(N__35879),
            .I(N__35874));
    LocalMux I__8031 (
            .O(N__35874),
            .I(N__35871));
    Odrv12 I__8030 (
            .O(N__35871),
            .I(\b2v_inst11.dutycycle_eena_3 ));
    CascadeMux I__8029 (
            .O(N__35868),
            .I(\b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1_cascade_ ));
    CascadeMux I__8028 (
            .O(N__35865),
            .I(N__35861));
    InMux I__8027 (
            .O(N__35864),
            .I(N__35853));
    InMux I__8026 (
            .O(N__35861),
            .I(N__35849));
    InMux I__8025 (
            .O(N__35860),
            .I(N__35846));
    InMux I__8024 (
            .O(N__35859),
            .I(N__35838));
    InMux I__8023 (
            .O(N__35858),
            .I(N__35838));
    InMux I__8022 (
            .O(N__35857),
            .I(N__35838));
    CascadeMux I__8021 (
            .O(N__35856),
            .I(N__35824));
    LocalMux I__8020 (
            .O(N__35853),
            .I(N__35821));
    CascadeMux I__8019 (
            .O(N__35852),
            .I(N__35818));
    LocalMux I__8018 (
            .O(N__35849),
            .I(N__35812));
    LocalMux I__8017 (
            .O(N__35846),
            .I(N__35812));
    InMux I__8016 (
            .O(N__35845),
            .I(N__35809));
    LocalMux I__8015 (
            .O(N__35838),
            .I(N__35805));
    InMux I__8014 (
            .O(N__35837),
            .I(N__35800));
    InMux I__8013 (
            .O(N__35836),
            .I(N__35800));
    InMux I__8012 (
            .O(N__35835),
            .I(N__35793));
    InMux I__8011 (
            .O(N__35834),
            .I(N__35793));
    InMux I__8010 (
            .O(N__35833),
            .I(N__35783));
    InMux I__8009 (
            .O(N__35832),
            .I(N__35783));
    CascadeMux I__8008 (
            .O(N__35831),
            .I(N__35776));
    InMux I__8007 (
            .O(N__35830),
            .I(N__35771));
    InMux I__8006 (
            .O(N__35829),
            .I(N__35771));
    IoInMux I__8005 (
            .O(N__35828),
            .I(N__35768));
    InMux I__8004 (
            .O(N__35827),
            .I(N__35765));
    InMux I__8003 (
            .O(N__35824),
            .I(N__35762));
    Span4Mux_s1_h I__8002 (
            .O(N__35821),
            .I(N__35759));
    InMux I__8001 (
            .O(N__35818),
            .I(N__35754));
    InMux I__8000 (
            .O(N__35817),
            .I(N__35754));
    Span4Mux_s1_h I__7999 (
            .O(N__35812),
            .I(N__35751));
    LocalMux I__7998 (
            .O(N__35809),
            .I(N__35748));
    InMux I__7997 (
            .O(N__35808),
            .I(N__35745));
    Span4Mux_s2_h I__7996 (
            .O(N__35805),
            .I(N__35742));
    LocalMux I__7995 (
            .O(N__35800),
            .I(N__35739));
    InMux I__7994 (
            .O(N__35799),
            .I(N__35736));
    InMux I__7993 (
            .O(N__35798),
            .I(N__35733));
    LocalMux I__7992 (
            .O(N__35793),
            .I(N__35730));
    InMux I__7991 (
            .O(N__35792),
            .I(N__35723));
    InMux I__7990 (
            .O(N__35791),
            .I(N__35723));
    InMux I__7989 (
            .O(N__35790),
            .I(N__35723));
    InMux I__7988 (
            .O(N__35789),
            .I(N__35720));
    InMux I__7987 (
            .O(N__35788),
            .I(N__35717));
    LocalMux I__7986 (
            .O(N__35783),
            .I(N__35714));
    InMux I__7985 (
            .O(N__35782),
            .I(N__35711));
    InMux I__7984 (
            .O(N__35781),
            .I(N__35708));
    InMux I__7983 (
            .O(N__35780),
            .I(N__35701));
    InMux I__7982 (
            .O(N__35779),
            .I(N__35701));
    InMux I__7981 (
            .O(N__35776),
            .I(N__35701));
    LocalMux I__7980 (
            .O(N__35771),
            .I(N__35698));
    LocalMux I__7979 (
            .O(N__35768),
            .I(N__35695));
    LocalMux I__7978 (
            .O(N__35765),
            .I(N__35692));
    LocalMux I__7977 (
            .O(N__35762),
            .I(N__35681));
    Span4Mux_v I__7976 (
            .O(N__35759),
            .I(N__35681));
    LocalMux I__7975 (
            .O(N__35754),
            .I(N__35681));
    Span4Mux_v I__7974 (
            .O(N__35751),
            .I(N__35681));
    Span4Mux_s1_h I__7973 (
            .O(N__35748),
            .I(N__35681));
    LocalMux I__7972 (
            .O(N__35745),
            .I(N__35678));
    Span4Mux_h I__7971 (
            .O(N__35742),
            .I(N__35675));
    Span4Mux_s2_h I__7970 (
            .O(N__35739),
            .I(N__35670));
    LocalMux I__7969 (
            .O(N__35736),
            .I(N__35670));
    LocalMux I__7968 (
            .O(N__35733),
            .I(N__35661));
    Span4Mux_s2_h I__7967 (
            .O(N__35730),
            .I(N__35661));
    LocalMux I__7966 (
            .O(N__35723),
            .I(N__35661));
    LocalMux I__7965 (
            .O(N__35720),
            .I(N__35661));
    LocalMux I__7964 (
            .O(N__35717),
            .I(N__35658));
    Span4Mux_v I__7963 (
            .O(N__35714),
            .I(N__35653));
    LocalMux I__7962 (
            .O(N__35711),
            .I(N__35653));
    LocalMux I__7961 (
            .O(N__35708),
            .I(N__35646));
    LocalMux I__7960 (
            .O(N__35701),
            .I(N__35646));
    Span4Mux_s2_h I__7959 (
            .O(N__35698),
            .I(N__35646));
    Span4Mux_s3_v I__7958 (
            .O(N__35695),
            .I(N__35643));
    Span4Mux_v I__7957 (
            .O(N__35692),
            .I(N__35638));
    Span4Mux_h I__7956 (
            .O(N__35681),
            .I(N__35638));
    Span12Mux_s5_h I__7955 (
            .O(N__35678),
            .I(N__35633));
    Sp12to4 I__7954 (
            .O(N__35675),
            .I(N__35633));
    Span4Mux_h I__7953 (
            .O(N__35670),
            .I(N__35628));
    Span4Mux_h I__7952 (
            .O(N__35661),
            .I(N__35628));
    Span4Mux_s2_h I__7951 (
            .O(N__35658),
            .I(N__35621));
    Span4Mux_v I__7950 (
            .O(N__35653),
            .I(N__35621));
    Span4Mux_v I__7949 (
            .O(N__35646),
            .I(N__35621));
    Odrv4 I__7948 (
            .O(N__35643),
            .I(G_149));
    Odrv4 I__7947 (
            .O(N__35638),
            .I(G_149));
    Odrv12 I__7946 (
            .O(N__35633),
            .I(G_149));
    Odrv4 I__7945 (
            .O(N__35628),
            .I(G_149));
    Odrv4 I__7944 (
            .O(N__35621),
            .I(G_149));
    CascadeMux I__7943 (
            .O(N__35610),
            .I(\b2v_inst11.dutycycleZ0Z_4_cascade_ ));
    InMux I__7942 (
            .O(N__35607),
            .I(N__35604));
    LocalMux I__7941 (
            .O(N__35604),
            .I(N__35601));
    Span4Mux_s1_h I__7940 (
            .O(N__35601),
            .I(N__35598));
    Odrv4 I__7939 (
            .O(N__35598),
            .I(\b2v_inst11.un1_dutycycle_94_s1_10 ));
    InMux I__7938 (
            .O(N__35595),
            .I(N__35592));
    LocalMux I__7937 (
            .O(N__35592),
            .I(\b2v_inst11.un1_dutycycle_94_s0_10 ));
    InMux I__7936 (
            .O(N__35589),
            .I(N__35586));
    LocalMux I__7935 (
            .O(N__35586),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642 ));
    CascadeMux I__7934 (
            .O(N__35583),
            .I(N__35580));
    InMux I__7933 (
            .O(N__35580),
            .I(N__35574));
    InMux I__7932 (
            .O(N__35579),
            .I(N__35574));
    LocalMux I__7931 (
            .O(N__35574),
            .I(\b2v_inst11.dutycycleZ1Z_10 ));
    InMux I__7930 (
            .O(N__35571),
            .I(N__35565));
    InMux I__7929 (
            .O(N__35570),
            .I(N__35565));
    LocalMux I__7928 (
            .O(N__35565),
            .I(N__35562));
    Odrv4 I__7927 (
            .O(N__35562),
            .I(\b2v_inst11.dutycycle_eena_4 ));
    CascadeMux I__7926 (
            .O(N__35559),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642_cascade_ ));
    InMux I__7925 (
            .O(N__35556),
            .I(N__35549));
    InMux I__7924 (
            .O(N__35555),
            .I(N__35549));
    CascadeMux I__7923 (
            .O(N__35554),
            .I(N__35546));
    LocalMux I__7922 (
            .O(N__35549),
            .I(N__35541));
    InMux I__7921 (
            .O(N__35546),
            .I(N__35538));
    InMux I__7920 (
            .O(N__35545),
            .I(N__35531));
    InMux I__7919 (
            .O(N__35544),
            .I(N__35531));
    Span4Mux_s1_v I__7918 (
            .O(N__35541),
            .I(N__35527));
    LocalMux I__7917 (
            .O(N__35538),
            .I(N__35524));
    InMux I__7916 (
            .O(N__35537),
            .I(N__35519));
    InMux I__7915 (
            .O(N__35536),
            .I(N__35519));
    LocalMux I__7914 (
            .O(N__35531),
            .I(N__35516));
    InMux I__7913 (
            .O(N__35530),
            .I(N__35513));
    Span4Mux_v I__7912 (
            .O(N__35527),
            .I(N__35510));
    Span4Mux_h I__7911 (
            .O(N__35524),
            .I(N__35507));
    LocalMux I__7910 (
            .O(N__35519),
            .I(N__35502));
    Span4Mux_h I__7909 (
            .O(N__35516),
            .I(N__35502));
    LocalMux I__7908 (
            .O(N__35513),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    Odrv4 I__7907 (
            .O(N__35510),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    Odrv4 I__7906 (
            .O(N__35507),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    Odrv4 I__7905 (
            .O(N__35502),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ));
    CascadeMux I__7904 (
            .O(N__35493),
            .I(\b2v_inst11.dutycycleZ0Z_3_cascade_ ));
    CascadeMux I__7903 (
            .O(N__35490),
            .I(N__35487));
    InMux I__7902 (
            .O(N__35487),
            .I(N__35481));
    InMux I__7901 (
            .O(N__35486),
            .I(N__35481));
    LocalMux I__7900 (
            .O(N__35481),
            .I(N__35478));
    Span4Mux_s3_v I__7899 (
            .O(N__35478),
            .I(N__35475));
    Odrv4 I__7898 (
            .O(N__35475),
            .I(\b2v_inst11.un1_dutycycle_53_44_0_1 ));
    InMux I__7897 (
            .O(N__35472),
            .I(N__35469));
    LocalMux I__7896 (
            .O(N__35469),
            .I(N__35458));
    InMux I__7895 (
            .O(N__35468),
            .I(N__35455));
    InMux I__7894 (
            .O(N__35467),
            .I(N__35450));
    InMux I__7893 (
            .O(N__35466),
            .I(N__35450));
    InMux I__7892 (
            .O(N__35465),
            .I(N__35445));
    InMux I__7891 (
            .O(N__35464),
            .I(N__35445));
    InMux I__7890 (
            .O(N__35463),
            .I(N__35442));
    CascadeMux I__7889 (
            .O(N__35462),
            .I(N__35439));
    CascadeMux I__7888 (
            .O(N__35461),
            .I(N__35436));
    Span4Mux_v I__7887 (
            .O(N__35458),
            .I(N__35429));
    LocalMux I__7886 (
            .O(N__35455),
            .I(N__35429));
    LocalMux I__7885 (
            .O(N__35450),
            .I(N__35424));
    LocalMux I__7884 (
            .O(N__35445),
            .I(N__35424));
    LocalMux I__7883 (
            .O(N__35442),
            .I(N__35419));
    InMux I__7882 (
            .O(N__35439),
            .I(N__35416));
    InMux I__7881 (
            .O(N__35436),
            .I(N__35413));
    CascadeMux I__7880 (
            .O(N__35435),
            .I(N__35410));
    InMux I__7879 (
            .O(N__35434),
            .I(N__35407));
    Span4Mux_s3_v I__7878 (
            .O(N__35429),
            .I(N__35404));
    Span4Mux_s3_v I__7877 (
            .O(N__35424),
            .I(N__35401));
    InMux I__7876 (
            .O(N__35423),
            .I(N__35398));
    InMux I__7875 (
            .O(N__35422),
            .I(N__35395));
    Span4Mux_s3_v I__7874 (
            .O(N__35419),
            .I(N__35388));
    LocalMux I__7873 (
            .O(N__35416),
            .I(N__35388));
    LocalMux I__7872 (
            .O(N__35413),
            .I(N__35388));
    InMux I__7871 (
            .O(N__35410),
            .I(N__35385));
    LocalMux I__7870 (
            .O(N__35407),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__7869 (
            .O(N__35404),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__7868 (
            .O(N__35401),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__7867 (
            .O(N__35398),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__7866 (
            .O(N__35395),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__7865 (
            .O(N__35388),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__7864 (
            .O(N__35385),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    InMux I__7863 (
            .O(N__35370),
            .I(N__35367));
    LocalMux I__7862 (
            .O(N__35367),
            .I(N__35364));
    Odrv4 I__7861 (
            .O(N__35364),
            .I(\b2v_inst11.g1_i_0 ));
    InMux I__7860 (
            .O(N__35361),
            .I(N__35358));
    LocalMux I__7859 (
            .O(N__35358),
            .I(N__35355));
    Span4Mux_v I__7858 (
            .O(N__35355),
            .I(N__35352));
    Odrv4 I__7857 (
            .O(N__35352),
            .I(\b2v_inst11.dutycycle_eena_2 ));
    InMux I__7856 (
            .O(N__35349),
            .I(N__35346));
    LocalMux I__7855 (
            .O(N__35346),
            .I(N__35342));
    InMux I__7854 (
            .O(N__35345),
            .I(N__35339));
    Span4Mux_v I__7853 (
            .O(N__35342),
            .I(N__35336));
    LocalMux I__7852 (
            .O(N__35339),
            .I(N__35331));
    Span4Mux_s0_h I__7851 (
            .O(N__35336),
            .I(N__35331));
    Odrv4 I__7850 (
            .O(N__35331),
            .I(\b2v_inst11.dutycycleZ1Z_9 ));
    CascadeMux I__7849 (
            .O(N__35328),
            .I(\b2v_inst11.dutycycle_eena_2_cascade_ ));
    InMux I__7848 (
            .O(N__35325),
            .I(N__35322));
    LocalMux I__7847 (
            .O(N__35322),
            .I(N__35319));
    Span4Mux_h I__7846 (
            .O(N__35319),
            .I(N__35315));
    InMux I__7845 (
            .O(N__35318),
            .I(N__35312));
    Span4Mux_v I__7844 (
            .O(N__35315),
            .I(N__35309));
    LocalMux I__7843 (
            .O(N__35312),
            .I(N__35306));
    Odrv4 I__7842 (
            .O(N__35309),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1 ));
    Odrv4 I__7841 (
            .O(N__35306),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1 ));
    CascadeMux I__7840 (
            .O(N__35301),
            .I(\b2v_inst11.dutycycleZ0Z_0_cascade_ ));
    CascadeMux I__7839 (
            .O(N__35298),
            .I(N__35295));
    InMux I__7838 (
            .O(N__35295),
            .I(N__35292));
    LocalMux I__7837 (
            .O(N__35292),
            .I(\b2v_inst11.un1_clk_100khz_30_and_i_0_0_1 ));
    CascadeMux I__7836 (
            .O(N__35289),
            .I(N__35286));
    InMux I__7835 (
            .O(N__35286),
            .I(N__35283));
    LocalMux I__7834 (
            .O(N__35283),
            .I(\b2v_inst11.un1_dutycycle_94_s0_5 ));
    InMux I__7833 (
            .O(N__35280),
            .I(N__35277));
    LocalMux I__7832 (
            .O(N__35277),
            .I(N__35274));
    Odrv4 I__7831 (
            .O(N__35274),
            .I(\b2v_inst11.un1_dutycycle_94_s1_5 ));
    InMux I__7830 (
            .O(N__35271),
            .I(N__35268));
    LocalMux I__7829 (
            .O(N__35268),
            .I(N__35265));
    Odrv12 I__7828 (
            .O(N__35265),
            .I(\b2v_inst11.N_302 ));
    InMux I__7827 (
            .O(N__35262),
            .I(N__35259));
    LocalMux I__7826 (
            .O(N__35259),
            .I(N__35256));
    Span4Mux_v I__7825 (
            .O(N__35256),
            .I(N__35253));
    Odrv4 I__7824 (
            .O(N__35253),
            .I(\b2v_inst11.un1_dutycycle_94_s1_6 ));
    InMux I__7823 (
            .O(N__35250),
            .I(N__35247));
    LocalMux I__7822 (
            .O(N__35247),
            .I(\b2v_inst11.un1_dutycycle_94_s0_6 ));
    InMux I__7821 (
            .O(N__35244),
            .I(N__35241));
    LocalMux I__7820 (
            .O(N__35241),
            .I(N__35238));
    Span4Mux_s0_h I__7819 (
            .O(N__35238),
            .I(N__35235));
    Odrv4 I__7818 (
            .O(N__35235),
            .I(\b2v_inst11.N_301 ));
    InMux I__7817 (
            .O(N__35232),
            .I(N__35229));
    LocalMux I__7816 (
            .O(N__35229),
            .I(N__35226));
    Odrv4 I__7815 (
            .O(N__35226),
            .I(\b2v_inst11.un1_dutycycle_94_s1_14 ));
    InMux I__7814 (
            .O(N__35223),
            .I(N__35220));
    LocalMux I__7813 (
            .O(N__35220),
            .I(N__35217));
    Odrv4 I__7812 (
            .O(N__35217),
            .I(\b2v_inst11.un1_dutycycle_94_s0_14 ));
    CascadeMux I__7811 (
            .O(N__35214),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0_cascade_ ));
    InMux I__7810 (
            .O(N__35211),
            .I(N__35206));
    CascadeMux I__7809 (
            .O(N__35210),
            .I(N__35200));
    CascadeMux I__7808 (
            .O(N__35209),
            .I(N__35196));
    LocalMux I__7807 (
            .O(N__35206),
            .I(N__35190));
    InMux I__7806 (
            .O(N__35205),
            .I(N__35185));
    InMux I__7805 (
            .O(N__35204),
            .I(N__35182));
    InMux I__7804 (
            .O(N__35203),
            .I(N__35177));
    InMux I__7803 (
            .O(N__35200),
            .I(N__35177));
    InMux I__7802 (
            .O(N__35199),
            .I(N__35170));
    InMux I__7801 (
            .O(N__35196),
            .I(N__35170));
    InMux I__7800 (
            .O(N__35195),
            .I(N__35170));
    CascadeMux I__7799 (
            .O(N__35194),
            .I(N__35166));
    InMux I__7798 (
            .O(N__35193),
            .I(N__35163));
    Span4Mux_v I__7797 (
            .O(N__35190),
            .I(N__35160));
    InMux I__7796 (
            .O(N__35189),
            .I(N__35157));
    InMux I__7795 (
            .O(N__35188),
            .I(N__35154));
    LocalMux I__7794 (
            .O(N__35185),
            .I(N__35149));
    LocalMux I__7793 (
            .O(N__35182),
            .I(N__35149));
    LocalMux I__7792 (
            .O(N__35177),
            .I(N__35146));
    LocalMux I__7791 (
            .O(N__35170),
            .I(N__35143));
    InMux I__7790 (
            .O(N__35169),
            .I(N__35138));
    InMux I__7789 (
            .O(N__35166),
            .I(N__35138));
    LocalMux I__7788 (
            .O(N__35163),
            .I(N__35135));
    Span4Mux_h I__7787 (
            .O(N__35160),
            .I(N__35120));
    LocalMux I__7786 (
            .O(N__35157),
            .I(N__35120));
    LocalMux I__7785 (
            .O(N__35154),
            .I(N__35120));
    Span4Mux_v I__7784 (
            .O(N__35149),
            .I(N__35120));
    Span4Mux_h I__7783 (
            .O(N__35146),
            .I(N__35120));
    Span4Mux_h I__7782 (
            .O(N__35143),
            .I(N__35120));
    LocalMux I__7781 (
            .O(N__35138),
            .I(N__35120));
    Odrv12 I__7780 (
            .O(N__35135),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    Odrv4 I__7779 (
            .O(N__35120),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    InMux I__7778 (
            .O(N__35115),
            .I(N__35112));
    LocalMux I__7777 (
            .O(N__35112),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0 ));
    InMux I__7776 (
            .O(N__35109),
            .I(N__35103));
    InMux I__7775 (
            .O(N__35108),
            .I(N__35103));
    LocalMux I__7774 (
            .O(N__35103),
            .I(N__35100));
    Odrv12 I__7773 (
            .O(N__35100),
            .I(\b2v_inst11.dutycycle_en_11 ));
    CascadeMux I__7772 (
            .O(N__35097),
            .I(N__35094));
    InMux I__7771 (
            .O(N__35094),
            .I(N__35088));
    InMux I__7770 (
            .O(N__35093),
            .I(N__35088));
    LocalMux I__7769 (
            .O(N__35088),
            .I(\b2v_inst11.dutycycleZ0Z_14 ));
    CascadeMux I__7768 (
            .O(N__35085),
            .I(N__35080));
    InMux I__7767 (
            .O(N__35084),
            .I(N__35077));
    CascadeMux I__7766 (
            .O(N__35083),
            .I(N__35074));
    InMux I__7765 (
            .O(N__35080),
            .I(N__35071));
    LocalMux I__7764 (
            .O(N__35077),
            .I(N__35066));
    InMux I__7763 (
            .O(N__35074),
            .I(N__35063));
    LocalMux I__7762 (
            .O(N__35071),
            .I(N__35060));
    InMux I__7761 (
            .O(N__35070),
            .I(N__35057));
    InMux I__7760 (
            .O(N__35069),
            .I(N__35054));
    Span4Mux_v I__7759 (
            .O(N__35066),
            .I(N__35049));
    LocalMux I__7758 (
            .O(N__35063),
            .I(N__35049));
    Span4Mux_s3_v I__7757 (
            .O(N__35060),
            .I(N__35046));
    LocalMux I__7756 (
            .O(N__35057),
            .I(N__35043));
    LocalMux I__7755 (
            .O(N__35054),
            .I(N__35038));
    Span4Mux_h I__7754 (
            .O(N__35049),
            .I(N__35038));
    Odrv4 I__7753 (
            .O(N__35046),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_10 ));
    Odrv12 I__7752 (
            .O(N__35043),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_10 ));
    Odrv4 I__7751 (
            .O(N__35038),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_10 ));
    CascadeMux I__7750 (
            .O(N__35031),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_ ));
    InMux I__7749 (
            .O(N__35028),
            .I(N__35020));
    InMux I__7748 (
            .O(N__35027),
            .I(N__35020));
    CascadeMux I__7747 (
            .O(N__35026),
            .I(N__35017));
    InMux I__7746 (
            .O(N__35025),
            .I(N__35012));
    LocalMux I__7745 (
            .O(N__35020),
            .I(N__35003));
    InMux I__7744 (
            .O(N__35017),
            .I(N__34997));
    InMux I__7743 (
            .O(N__35016),
            .I(N__34997));
    InMux I__7742 (
            .O(N__35015),
            .I(N__34994));
    LocalMux I__7741 (
            .O(N__35012),
            .I(N__34990));
    InMux I__7740 (
            .O(N__35011),
            .I(N__34987));
    CascadeMux I__7739 (
            .O(N__35010),
            .I(N__34983));
    CascadeMux I__7738 (
            .O(N__35009),
            .I(N__34979));
    InMux I__7737 (
            .O(N__35008),
            .I(N__34969));
    InMux I__7736 (
            .O(N__35007),
            .I(N__34969));
    InMux I__7735 (
            .O(N__35006),
            .I(N__34969));
    Span4Mux_h I__7734 (
            .O(N__35003),
            .I(N__34966));
    InMux I__7733 (
            .O(N__35002),
            .I(N__34963));
    LocalMux I__7732 (
            .O(N__34997),
            .I(N__34959));
    LocalMux I__7731 (
            .O(N__34994),
            .I(N__34956));
    CascadeMux I__7730 (
            .O(N__34993),
            .I(N__34950));
    Span4Mux_s3_h I__7729 (
            .O(N__34990),
            .I(N__34947));
    LocalMux I__7728 (
            .O(N__34987),
            .I(N__34944));
    InMux I__7727 (
            .O(N__34986),
            .I(N__34941));
    InMux I__7726 (
            .O(N__34983),
            .I(N__34936));
    InMux I__7725 (
            .O(N__34982),
            .I(N__34936));
    InMux I__7724 (
            .O(N__34979),
            .I(N__34933));
    InMux I__7723 (
            .O(N__34978),
            .I(N__34926));
    InMux I__7722 (
            .O(N__34977),
            .I(N__34926));
    InMux I__7721 (
            .O(N__34976),
            .I(N__34926));
    LocalMux I__7720 (
            .O(N__34969),
            .I(N__34923));
    Sp12to4 I__7719 (
            .O(N__34966),
            .I(N__34918));
    LocalMux I__7718 (
            .O(N__34963),
            .I(N__34918));
    InMux I__7717 (
            .O(N__34962),
            .I(N__34915));
    Span4Mux_s3_v I__7716 (
            .O(N__34959),
            .I(N__34910));
    Span4Mux_s0_h I__7715 (
            .O(N__34956),
            .I(N__34910));
    InMux I__7714 (
            .O(N__34955),
            .I(N__34901));
    InMux I__7713 (
            .O(N__34954),
            .I(N__34901));
    InMux I__7712 (
            .O(N__34953),
            .I(N__34901));
    InMux I__7711 (
            .O(N__34950),
            .I(N__34901));
    Odrv4 I__7710 (
            .O(N__34947),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv12 I__7709 (
            .O(N__34944),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__7708 (
            .O(N__34941),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__7707 (
            .O(N__34936),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__7706 (
            .O(N__34933),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__7705 (
            .O(N__34926),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__7704 (
            .O(N__34923),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv12 I__7703 (
            .O(N__34918),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__7702 (
            .O(N__34915),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__7701 (
            .O(N__34910),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__7700 (
            .O(N__34901),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    CascadeMux I__7699 (
            .O(N__34878),
            .I(\b2v_inst11.un1_dutycycle_53_44_0_3_tz_1_cascade_ ));
    InMux I__7698 (
            .O(N__34875),
            .I(N__34871));
    InMux I__7697 (
            .O(N__34874),
            .I(N__34868));
    LocalMux I__7696 (
            .O(N__34871),
            .I(N__34865));
    LocalMux I__7695 (
            .O(N__34868),
            .I(N__34862));
    Span4Mux_s3_v I__7694 (
            .O(N__34865),
            .I(N__34859));
    Odrv4 I__7693 (
            .O(N__34862),
            .I(\b2v_inst11.un1_dutycycle_53_44_1 ));
    Odrv4 I__7692 (
            .O(N__34859),
            .I(\b2v_inst11.un1_dutycycle_53_44_1 ));
    InMux I__7691 (
            .O(N__34854),
            .I(N__34851));
    LocalMux I__7690 (
            .O(N__34851),
            .I(N__34848));
    Span4Mux_s3_h I__7689 (
            .O(N__34848),
            .I(N__34845));
    Odrv4 I__7688 (
            .O(N__34845),
            .I(\b2v_inst11.g3_0_0 ));
    IoInMux I__7687 (
            .O(N__34842),
            .I(N__34839));
    LocalMux I__7686 (
            .O(N__34839),
            .I(N__34834));
    InMux I__7685 (
            .O(N__34838),
            .I(N__34830));
    CascadeMux I__7684 (
            .O(N__34837),
            .I(N__34827));
    IoSpan4Mux I__7683 (
            .O(N__34834),
            .I(N__34824));
    InMux I__7682 (
            .O(N__34833),
            .I(N__34820));
    LocalMux I__7681 (
            .O(N__34830),
            .I(N__34814));
    InMux I__7680 (
            .O(N__34827),
            .I(N__34811));
    IoSpan4Mux I__7679 (
            .O(N__34824),
            .I(N__34808));
    InMux I__7678 (
            .O(N__34823),
            .I(N__34805));
    LocalMux I__7677 (
            .O(N__34820),
            .I(N__34802));
    InMux I__7676 (
            .O(N__34819),
            .I(N__34797));
    CascadeMux I__7675 (
            .O(N__34818),
            .I(N__34794));
    InMux I__7674 (
            .O(N__34817),
            .I(N__34791));
    Span4Mux_v I__7673 (
            .O(N__34814),
            .I(N__34786));
    LocalMux I__7672 (
            .O(N__34811),
            .I(N__34786));
    Span4Mux_s3_v I__7671 (
            .O(N__34808),
            .I(N__34781));
    LocalMux I__7670 (
            .O(N__34805),
            .I(N__34781));
    Span4Mux_s3_h I__7669 (
            .O(N__34802),
            .I(N__34778));
    InMux I__7668 (
            .O(N__34801),
            .I(N__34775));
    InMux I__7667 (
            .O(N__34800),
            .I(N__34772));
    LocalMux I__7666 (
            .O(N__34797),
            .I(N__34766));
    InMux I__7665 (
            .O(N__34794),
            .I(N__34763));
    LocalMux I__7664 (
            .O(N__34791),
            .I(N__34760));
    Span4Mux_v I__7663 (
            .O(N__34786),
            .I(N__34757));
    Span4Mux_v I__7662 (
            .O(N__34781),
            .I(N__34748));
    Span4Mux_h I__7661 (
            .O(N__34778),
            .I(N__34748));
    LocalMux I__7660 (
            .O(N__34775),
            .I(N__34748));
    LocalMux I__7659 (
            .O(N__34772),
            .I(N__34748));
    InMux I__7658 (
            .O(N__34771),
            .I(N__34741));
    InMux I__7657 (
            .O(N__34770),
            .I(N__34741));
    InMux I__7656 (
            .O(N__34769),
            .I(N__34741));
    Span4Mux_s3_h I__7655 (
            .O(N__34766),
            .I(N__34738));
    LocalMux I__7654 (
            .O(N__34763),
            .I(rsmrstn));
    Odrv4 I__7653 (
            .O(N__34760),
            .I(rsmrstn));
    Odrv4 I__7652 (
            .O(N__34757),
            .I(rsmrstn));
    Odrv4 I__7651 (
            .O(N__34748),
            .I(rsmrstn));
    LocalMux I__7650 (
            .O(N__34741),
            .I(rsmrstn));
    Odrv4 I__7649 (
            .O(N__34738),
            .I(rsmrstn));
    CascadeMux I__7648 (
            .O(N__34725),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_7_cascade_ ));
    InMux I__7647 (
            .O(N__34722),
            .I(N__34719));
    LocalMux I__7646 (
            .O(N__34719),
            .I(\b2v_inst11.g1_0_0 ));
    InMux I__7645 (
            .O(N__34716),
            .I(N__34713));
    LocalMux I__7644 (
            .O(N__34713),
            .I(\b2v_inst11.un1_clk_100khz_36_and_i_0_0 ));
    InMux I__7643 (
            .O(N__34710),
            .I(N__34707));
    LocalMux I__7642 (
            .O(N__34707),
            .I(N__34704));
    Span4Mux_s1_h I__7641 (
            .O(N__34704),
            .I(N__34701));
    Odrv4 I__7640 (
            .O(N__34701),
            .I(\b2v_inst11.un1_dutycycle_94_s1_7 ));
    InMux I__7639 (
            .O(N__34698),
            .I(N__34695));
    LocalMux I__7638 (
            .O(N__34695),
            .I(N__34692));
    Span4Mux_s0_h I__7637 (
            .O(N__34692),
            .I(N__34689));
    Odrv4 I__7636 (
            .O(N__34689),
            .I(\b2v_inst11.un1_dutycycle_94_s0_7 ));
    InMux I__7635 (
            .O(N__34686),
            .I(N__34683));
    LocalMux I__7634 (
            .O(N__34683),
            .I(\b2v_inst11.un1_dutycycle_94_0_7 ));
    InMux I__7633 (
            .O(N__34680),
            .I(N__34677));
    LocalMux I__7632 (
            .O(N__34677),
            .I(\b2v_inst11.g0_0_1_0 ));
    InMux I__7631 (
            .O(N__34674),
            .I(N__34668));
    InMux I__7630 (
            .O(N__34673),
            .I(N__34668));
    LocalMux I__7629 (
            .O(N__34668),
            .I(\b2v_inst11.dutycycleZ1Z_7 ));
    CascadeMux I__7628 (
            .O(N__34665),
            .I(\b2v_inst11.un1_dutycycle_94_0_7_cascade_ ));
    InMux I__7627 (
            .O(N__34662),
            .I(N__34659));
    LocalMux I__7626 (
            .O(N__34659),
            .I(N__34656));
    Span4Mux_s1_h I__7625 (
            .O(N__34656),
            .I(N__34653));
    Odrv4 I__7624 (
            .O(N__34653),
            .I(\b2v_inst11.un1_dutycycle_94_s1_13 ));
    InMux I__7623 (
            .O(N__34650),
            .I(N__34647));
    LocalMux I__7622 (
            .O(N__34647),
            .I(N__34644));
    Odrv4 I__7621 (
            .O(N__34644),
            .I(\b2v_inst11.un1_dutycycle_94_s0_13 ));
    InMux I__7620 (
            .O(N__34641),
            .I(N__34638));
    LocalMux I__7619 (
            .O(N__34638),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0 ));
    CascadeMux I__7618 (
            .O(N__34635),
            .I(N__34632));
    InMux I__7617 (
            .O(N__34632),
            .I(N__34626));
    InMux I__7616 (
            .O(N__34631),
            .I(N__34626));
    LocalMux I__7615 (
            .O(N__34626),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    InMux I__7614 (
            .O(N__34623),
            .I(N__34617));
    InMux I__7613 (
            .O(N__34622),
            .I(N__34617));
    LocalMux I__7612 (
            .O(N__34617),
            .I(N__34614));
    Odrv12 I__7611 (
            .O(N__34614),
            .I(\b2v_inst11.dutycycle_en_10 ));
    CascadeMux I__7610 (
            .O(N__34611),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0_cascade_ ));
    CascadeMux I__7609 (
            .O(N__34608),
            .I(N__34601));
    InMux I__7608 (
            .O(N__34607),
            .I(N__34595));
    InMux I__7607 (
            .O(N__34606),
            .I(N__34592));
    InMux I__7606 (
            .O(N__34605),
            .I(N__34588));
    InMux I__7605 (
            .O(N__34604),
            .I(N__34585));
    InMux I__7604 (
            .O(N__34601),
            .I(N__34580));
    InMux I__7603 (
            .O(N__34600),
            .I(N__34580));
    InMux I__7602 (
            .O(N__34599),
            .I(N__34575));
    InMux I__7601 (
            .O(N__34598),
            .I(N__34575));
    LocalMux I__7600 (
            .O(N__34595),
            .I(N__34570));
    LocalMux I__7599 (
            .O(N__34592),
            .I(N__34570));
    InMux I__7598 (
            .O(N__34591),
            .I(N__34564));
    LocalMux I__7597 (
            .O(N__34588),
            .I(N__34560));
    LocalMux I__7596 (
            .O(N__34585),
            .I(N__34557));
    LocalMux I__7595 (
            .O(N__34580),
            .I(N__34552));
    LocalMux I__7594 (
            .O(N__34575),
            .I(N__34552));
    Span4Mux_v I__7593 (
            .O(N__34570),
            .I(N__34549));
    InMux I__7592 (
            .O(N__34569),
            .I(N__34544));
    InMux I__7591 (
            .O(N__34568),
            .I(N__34544));
    InMux I__7590 (
            .O(N__34567),
            .I(N__34541));
    LocalMux I__7589 (
            .O(N__34564),
            .I(N__34538));
    InMux I__7588 (
            .O(N__34563),
            .I(N__34535));
    Span4Mux_v I__7587 (
            .O(N__34560),
            .I(N__34528));
    Span4Mux_v I__7586 (
            .O(N__34557),
            .I(N__34528));
    Span4Mux_v I__7585 (
            .O(N__34552),
            .I(N__34528));
    Span4Mux_s0_h I__7584 (
            .O(N__34549),
            .I(N__34521));
    LocalMux I__7583 (
            .O(N__34544),
            .I(N__34521));
    LocalMux I__7582 (
            .O(N__34541),
            .I(N__34521));
    Odrv12 I__7581 (
            .O(N__34538),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__7580 (
            .O(N__34535),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__7579 (
            .O(N__34528),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__7578 (
            .O(N__34521),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    CascadeMux I__7577 (
            .O(N__34512),
            .I(\b2v_inst11.un1_clk_100khz_32_and_i_0_c_0_cascade_ ));
    InMux I__7576 (
            .O(N__34509),
            .I(N__34503));
    InMux I__7575 (
            .O(N__34508),
            .I(N__34503));
    LocalMux I__7574 (
            .O(N__34503),
            .I(\b2v_inst11.un1_clk_100khz_32_and_i_0_d ));
    CascadeMux I__7573 (
            .O(N__34500),
            .I(\b2v_inst11.un1_clk_100khz_33_and_i_0_c_0_cascade_ ));
    InMux I__7572 (
            .O(N__34497),
            .I(N__34494));
    LocalMux I__7571 (
            .O(N__34494),
            .I(\b2v_inst11.N_153_N ));
    CascadeMux I__7570 (
            .O(N__34491),
            .I(\b2v_inst11.N_155_N_cascade_ ));
    CascadeMux I__7569 (
            .O(N__34488),
            .I(\b2v_inst11.g0_0_1_0_cascade_ ));
    InMux I__7568 (
            .O(N__34485),
            .I(N__34482));
    LocalMux I__7567 (
            .O(N__34482),
            .I(\b2v_inst11.g0_1_1 ));
    CascadeMux I__7566 (
            .O(N__34479),
            .I(\b2v_inst11.dutycycle_set_1_cascade_ ));
    InMux I__7565 (
            .O(N__34476),
            .I(N__34473));
    LocalMux I__7564 (
            .O(N__34473),
            .I(N__34470));
    Span4Mux_s0_h I__7563 (
            .O(N__34470),
            .I(N__34467));
    Span4Mux_h I__7562 (
            .O(N__34467),
            .I(N__34463));
    InMux I__7561 (
            .O(N__34466),
            .I(N__34460));
    Odrv4 I__7560 (
            .O(N__34463),
            .I(\b2v_inst11.dutycycle_eena_14_0 ));
    LocalMux I__7559 (
            .O(N__34460),
            .I(\b2v_inst11.dutycycle_eena_14_0 ));
    InMux I__7558 (
            .O(N__34455),
            .I(N__34452));
    LocalMux I__7557 (
            .O(N__34452),
            .I(N__34448));
    InMux I__7556 (
            .O(N__34451),
            .I(N__34445));
    Span4Mux_h I__7555 (
            .O(N__34448),
            .I(N__34442));
    LocalMux I__7554 (
            .O(N__34445),
            .I(\b2v_inst11.dutycycle_0_5 ));
    Odrv4 I__7553 (
            .O(N__34442),
            .I(\b2v_inst11.dutycycle_0_5 ));
    CascadeMux I__7552 (
            .O(N__34437),
            .I(\b2v_inst11.dutycycle_RNIOFQO2Z0Z_3_cascade_ ));
    InMux I__7551 (
            .O(N__34434),
            .I(N__34431));
    LocalMux I__7550 (
            .O(N__34431),
            .I(N__34428));
    Span4Mux_v I__7549 (
            .O(N__34428),
            .I(N__34425));
    Odrv4 I__7548 (
            .O(N__34425),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJZ0Z9 ));
    InMux I__7547 (
            .O(N__34422),
            .I(N__34419));
    LocalMux I__7546 (
            .O(N__34419),
            .I(\b2v_inst11.dutycycle_RNIM98E2Z0Z_3 ));
    CascadeMux I__7545 (
            .O(N__34416),
            .I(N__34413));
    InMux I__7544 (
            .O(N__34413),
            .I(N__34408));
    InMux I__7543 (
            .O(N__34412),
            .I(N__34403));
    InMux I__7542 (
            .O(N__34411),
            .I(N__34403));
    LocalMux I__7541 (
            .O(N__34408),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    LocalMux I__7540 (
            .O(N__34403),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    CascadeMux I__7539 (
            .O(N__34398),
            .I(\b2v_inst11.dutycycle_RNIM98E2Z0Z_3_cascade_ ));
    InMux I__7538 (
            .O(N__34395),
            .I(N__34392));
    LocalMux I__7537 (
            .O(N__34392),
            .I(\b2v_inst11.dutycycle_RNIOFQO2Z0Z_3 ));
    InMux I__7536 (
            .O(N__34389),
            .I(N__34384));
    InMux I__7535 (
            .O(N__34388),
            .I(N__34373));
    InMux I__7534 (
            .O(N__34387),
            .I(N__34373));
    LocalMux I__7533 (
            .O(N__34384),
            .I(N__34370));
    InMux I__7532 (
            .O(N__34383),
            .I(N__34363));
    InMux I__7531 (
            .O(N__34382),
            .I(N__34363));
    InMux I__7530 (
            .O(N__34381),
            .I(N__34357));
    InMux I__7529 (
            .O(N__34380),
            .I(N__34357));
    CascadeMux I__7528 (
            .O(N__34379),
            .I(N__34351));
    InMux I__7527 (
            .O(N__34378),
            .I(N__34348));
    LocalMux I__7526 (
            .O(N__34373),
            .I(N__34343));
    Span4Mux_v I__7525 (
            .O(N__34370),
            .I(N__34343));
    InMux I__7524 (
            .O(N__34369),
            .I(N__34338));
    InMux I__7523 (
            .O(N__34368),
            .I(N__34338));
    LocalMux I__7522 (
            .O(N__34363),
            .I(N__34335));
    InMux I__7521 (
            .O(N__34362),
            .I(N__34332));
    LocalMux I__7520 (
            .O(N__34357),
            .I(N__34329));
    InMux I__7519 (
            .O(N__34356),
            .I(N__34324));
    InMux I__7518 (
            .O(N__34355),
            .I(N__34324));
    InMux I__7517 (
            .O(N__34354),
            .I(N__34319));
    InMux I__7516 (
            .O(N__34351),
            .I(N__34316));
    LocalMux I__7515 (
            .O(N__34348),
            .I(N__34309));
    Span4Mux_h I__7514 (
            .O(N__34343),
            .I(N__34309));
    LocalMux I__7513 (
            .O(N__34338),
            .I(N__34309));
    Span4Mux_s3_v I__7512 (
            .O(N__34335),
            .I(N__34306));
    LocalMux I__7511 (
            .O(N__34332),
            .I(N__34303));
    Span4Mux_h I__7510 (
            .O(N__34329),
            .I(N__34298));
    LocalMux I__7509 (
            .O(N__34324),
            .I(N__34298));
    CascadeMux I__7508 (
            .O(N__34323),
            .I(N__34295));
    InMux I__7507 (
            .O(N__34322),
            .I(N__34292));
    LocalMux I__7506 (
            .O(N__34319),
            .I(N__34285));
    LocalMux I__7505 (
            .O(N__34316),
            .I(N__34285));
    Span4Mux_v I__7504 (
            .O(N__34309),
            .I(N__34285));
    Span4Mux_v I__7503 (
            .O(N__34306),
            .I(N__34278));
    Span4Mux_h I__7502 (
            .O(N__34303),
            .I(N__34278));
    Span4Mux_v I__7501 (
            .O(N__34298),
            .I(N__34278));
    InMux I__7500 (
            .O(N__34295),
            .I(N__34275));
    LocalMux I__7499 (
            .O(N__34292),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__7498 (
            .O(N__34285),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__7497 (
            .O(N__34278),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__7496 (
            .O(N__34275),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    InMux I__7495 (
            .O(N__34266),
            .I(N__34262));
    InMux I__7494 (
            .O(N__34265),
            .I(N__34255));
    LocalMux I__7493 (
            .O(N__34262),
            .I(N__34252));
    InMux I__7492 (
            .O(N__34261),
            .I(N__34242));
    InMux I__7491 (
            .O(N__34260),
            .I(N__34242));
    InMux I__7490 (
            .O(N__34259),
            .I(N__34242));
    InMux I__7489 (
            .O(N__34258),
            .I(N__34242));
    LocalMux I__7488 (
            .O(N__34255),
            .I(N__34235));
    Span4Mux_s1_h I__7487 (
            .O(N__34252),
            .I(N__34235));
    InMux I__7486 (
            .O(N__34251),
            .I(N__34232));
    LocalMux I__7485 (
            .O(N__34242),
            .I(N__34229));
    InMux I__7484 (
            .O(N__34241),
            .I(N__34224));
    InMux I__7483 (
            .O(N__34240),
            .I(N__34224));
    Span4Mux_h I__7482 (
            .O(N__34235),
            .I(N__34221));
    LocalMux I__7481 (
            .O(N__34232),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    Odrv4 I__7480 (
            .O(N__34229),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    LocalMux I__7479 (
            .O(N__34224),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    Odrv4 I__7478 (
            .O(N__34221),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    CascadeMux I__7477 (
            .O(N__34212),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3_cascade_ ));
    CascadeMux I__7476 (
            .O(N__34209),
            .I(N__34206));
    InMux I__7475 (
            .O(N__34206),
            .I(N__34203));
    LocalMux I__7474 (
            .O(N__34203),
            .I(N__34200));
    Span4Mux_v I__7473 (
            .O(N__34200),
            .I(N__34197));
    Odrv4 I__7472 (
            .O(N__34197),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_s0_sf ));
    CascadeMux I__7471 (
            .O(N__34194),
            .I(N__34190));
    CascadeMux I__7470 (
            .O(N__34193),
            .I(N__34184));
    InMux I__7469 (
            .O(N__34190),
            .I(N__34178));
    InMux I__7468 (
            .O(N__34189),
            .I(N__34178));
    InMux I__7467 (
            .O(N__34188),
            .I(N__34175));
    InMux I__7466 (
            .O(N__34187),
            .I(N__34170));
    InMux I__7465 (
            .O(N__34184),
            .I(N__34170));
    InMux I__7464 (
            .O(N__34183),
            .I(N__34167));
    LocalMux I__7463 (
            .O(N__34178),
            .I(N__34156));
    LocalMux I__7462 (
            .O(N__34175),
            .I(N__34156));
    LocalMux I__7461 (
            .O(N__34170),
            .I(N__34156));
    LocalMux I__7460 (
            .O(N__34167),
            .I(N__34156));
    InMux I__7459 (
            .O(N__34166),
            .I(N__34153));
    InMux I__7458 (
            .O(N__34165),
            .I(N__34150));
    Span4Mux_v I__7457 (
            .O(N__34156),
            .I(N__34147));
    LocalMux I__7456 (
            .O(N__34153),
            .I(N__34144));
    LocalMux I__7455 (
            .O(N__34150),
            .I(N__34141));
    Span4Mux_v I__7454 (
            .O(N__34147),
            .I(N__34136));
    Span4Mux_v I__7453 (
            .O(N__34144),
            .I(N__34136));
    Odrv12 I__7452 (
            .O(N__34141),
            .I(\b2v_inst11.count_clk_RNIG510TZ0Z_7 ));
    Odrv4 I__7451 (
            .O(N__34136),
            .I(\b2v_inst11.count_clk_RNIG510TZ0Z_7 ));
    InMux I__7450 (
            .O(N__34131),
            .I(N__34128));
    LocalMux I__7449 (
            .O(N__34128),
            .I(N__34125));
    Span4Mux_s0_h I__7448 (
            .O(N__34125),
            .I(N__34122));
    Odrv4 I__7447 (
            .O(N__34122),
            .I(\b2v_inst11.N_305 ));
    InMux I__7446 (
            .O(N__34119),
            .I(N__34116));
    LocalMux I__7445 (
            .O(N__34116),
            .I(N__34113));
    Odrv12 I__7444 (
            .O(N__34113),
            .I(\b2v_inst11.N_306 ));
    CascadeMux I__7443 (
            .O(N__34110),
            .I(\b2v_inst11.N_231_N_cascade_ ));
    CascadeMux I__7442 (
            .O(N__34107),
            .I(\b2v_inst11.dutycycle_eena_13_cascade_ ));
    InMux I__7441 (
            .O(N__34104),
            .I(N__34101));
    LocalMux I__7440 (
            .O(N__34101),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4 ));
    InMux I__7439 (
            .O(N__34098),
            .I(N__34092));
    InMux I__7438 (
            .O(N__34097),
            .I(N__34092));
    LocalMux I__7437 (
            .O(N__34092),
            .I(\b2v_inst11.dutycycle_0_6 ));
    CascadeMux I__7436 (
            .O(N__34089),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4_cascade_ ));
    InMux I__7435 (
            .O(N__34086),
            .I(N__34083));
    LocalMux I__7434 (
            .O(N__34083),
            .I(\b2v_inst11.dutycycle_eena_13 ));
    InMux I__7433 (
            .O(N__34080),
            .I(N__34077));
    LocalMux I__7432 (
            .O(N__34077),
            .I(N__34074));
    Span4Mux_s2_h I__7431 (
            .O(N__34074),
            .I(N__34071));
    Odrv4 I__7430 (
            .O(N__34071),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    CascadeMux I__7429 (
            .O(N__34068),
            .I(\b2v_inst11.dutycycleZ1Z_6_cascade_ ));
    InMux I__7428 (
            .O(N__34065),
            .I(N__34062));
    LocalMux I__7427 (
            .O(N__34062),
            .I(\b2v_inst11.dutycycle_RNILF063Z0Z_6 ));
    InMux I__7426 (
            .O(N__34059),
            .I(N__34055));
    InMux I__7425 (
            .O(N__34058),
            .I(N__34052));
    LocalMux I__7424 (
            .O(N__34055),
            .I(N__34042));
    LocalMux I__7423 (
            .O(N__34052),
            .I(N__34042));
    InMux I__7422 (
            .O(N__34051),
            .I(N__34037));
    InMux I__7421 (
            .O(N__34050),
            .I(N__34037));
    CascadeMux I__7420 (
            .O(N__34049),
            .I(N__34033));
    CascadeMux I__7419 (
            .O(N__34048),
            .I(N__34027));
    CascadeMux I__7418 (
            .O(N__34047),
            .I(N__34021));
    Span4Mux_v I__7417 (
            .O(N__34042),
            .I(N__34018));
    LocalMux I__7416 (
            .O(N__34037),
            .I(N__34015));
    InMux I__7415 (
            .O(N__34036),
            .I(N__34008));
    InMux I__7414 (
            .O(N__34033),
            .I(N__34008));
    InMux I__7413 (
            .O(N__34032),
            .I(N__34008));
    InMux I__7412 (
            .O(N__34031),
            .I(N__34005));
    InMux I__7411 (
            .O(N__34030),
            .I(N__34000));
    InMux I__7410 (
            .O(N__34027),
            .I(N__34000));
    InMux I__7409 (
            .O(N__34026),
            .I(N__33995));
    InMux I__7408 (
            .O(N__34025),
            .I(N__33995));
    InMux I__7407 (
            .O(N__34024),
            .I(N__33992));
    InMux I__7406 (
            .O(N__34021),
            .I(N__33989));
    IoSpan4Mux I__7405 (
            .O(N__34018),
            .I(N__33984));
    Span4Mux_h I__7404 (
            .O(N__34015),
            .I(N__33984));
    LocalMux I__7403 (
            .O(N__34008),
            .I(N__33981));
    LocalMux I__7402 (
            .O(N__34005),
            .I(N__33976));
    LocalMux I__7401 (
            .O(N__34000),
            .I(N__33976));
    LocalMux I__7400 (
            .O(N__33995),
            .I(N__33973));
    LocalMux I__7399 (
            .O(N__33992),
            .I(N__33970));
    LocalMux I__7398 (
            .O(N__33989),
            .I(N__33967));
    Span4Mux_s1_h I__7397 (
            .O(N__33984),
            .I(N__33964));
    Span4Mux_h I__7396 (
            .O(N__33981),
            .I(N__33961));
    Span4Mux_v I__7395 (
            .O(N__33976),
            .I(N__33958));
    Span12Mux_s1_h I__7394 (
            .O(N__33973),
            .I(N__33955));
    Odrv12 I__7393 (
            .O(N__33970),
            .I(\b2v_inst11.N_172 ));
    Odrv12 I__7392 (
            .O(N__33967),
            .I(\b2v_inst11.N_172 ));
    Odrv4 I__7391 (
            .O(N__33964),
            .I(\b2v_inst11.N_172 ));
    Odrv4 I__7390 (
            .O(N__33961),
            .I(\b2v_inst11.N_172 ));
    Odrv4 I__7389 (
            .O(N__33958),
            .I(\b2v_inst11.N_172 ));
    Odrv12 I__7388 (
            .O(N__33955),
            .I(\b2v_inst11.N_172 ));
    InMux I__7387 (
            .O(N__33942),
            .I(N__33935));
    InMux I__7386 (
            .O(N__33941),
            .I(N__33935));
    InMux I__7385 (
            .O(N__33940),
            .I(N__33932));
    LocalMux I__7384 (
            .O(N__33935),
            .I(N__33929));
    LocalMux I__7383 (
            .O(N__33932),
            .I(\b2v_inst11.N_185 ));
    Odrv12 I__7382 (
            .O(N__33929),
            .I(\b2v_inst11.N_185 ));
    CascadeMux I__7381 (
            .O(N__33924),
            .I(N__33921));
    InMux I__7380 (
            .O(N__33921),
            .I(N__33918));
    LocalMux I__7379 (
            .O(N__33918),
            .I(N__33915));
    Span4Mux_h I__7378 (
            .O(N__33915),
            .I(N__33912));
    Odrv4 I__7377 (
            .O(N__33912),
            .I(\b2v_inst11.dutycycle_set_1 ));
    InMux I__7376 (
            .O(N__33909),
            .I(N__33906));
    LocalMux I__7375 (
            .O(N__33906),
            .I(N__33902));
    InMux I__7374 (
            .O(N__33905),
            .I(N__33899));
    Odrv4 I__7373 (
            .O(N__33902),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    LocalMux I__7372 (
            .O(N__33899),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    InMux I__7371 (
            .O(N__33894),
            .I(N__33888));
    InMux I__7370 (
            .O(N__33893),
            .I(N__33888));
    LocalMux I__7369 (
            .O(N__33888),
            .I(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ));
    InMux I__7368 (
            .O(N__33885),
            .I(N__33882));
    LocalMux I__7367 (
            .O(N__33882),
            .I(\b2v_inst11.count_clk_0_15 ));
    InMux I__7366 (
            .O(N__33879),
            .I(N__33876));
    LocalMux I__7365 (
            .O(N__33876),
            .I(N__33873));
    Span4Mux_h I__7364 (
            .O(N__33873),
            .I(N__33870));
    Span4Mux_v I__7363 (
            .O(N__33870),
            .I(N__33866));
    InMux I__7362 (
            .O(N__33869),
            .I(N__33863));
    Span4Mux_v I__7361 (
            .O(N__33866),
            .I(N__33860));
    LocalMux I__7360 (
            .O(N__33863),
            .I(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ));
    Odrv4 I__7359 (
            .O(N__33860),
            .I(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ));
    InMux I__7358 (
            .O(N__33855),
            .I(N__33852));
    LocalMux I__7357 (
            .O(N__33852),
            .I(N__33849));
    Span4Mux_s1_h I__7356 (
            .O(N__33849),
            .I(N__33846));
    Span4Mux_v I__7355 (
            .O(N__33846),
            .I(N__33843));
    Span4Mux_h I__7354 (
            .O(N__33843),
            .I(N__33840));
    Odrv4 I__7353 (
            .O(N__33840),
            .I(\b2v_inst11.count_clk_0_6 ));
    CEMux I__7352 (
            .O(N__33837),
            .I(N__33832));
    CEMux I__7351 (
            .O(N__33836),
            .I(N__33827));
    CEMux I__7350 (
            .O(N__33835),
            .I(N__33819));
    LocalMux I__7349 (
            .O(N__33832),
            .I(N__33816));
    CascadeMux I__7348 (
            .O(N__33831),
            .I(N__33813));
    CascadeMux I__7347 (
            .O(N__33830),
            .I(N__33804));
    LocalMux I__7346 (
            .O(N__33827),
            .I(N__33798));
    CascadeMux I__7345 (
            .O(N__33826),
            .I(N__33793));
    CascadeMux I__7344 (
            .O(N__33825),
            .I(N__33790));
    CascadeMux I__7343 (
            .O(N__33824),
            .I(N__33787));
    CascadeMux I__7342 (
            .O(N__33823),
            .I(N__33783));
    CEMux I__7341 (
            .O(N__33822),
            .I(N__33780));
    LocalMux I__7340 (
            .O(N__33819),
            .I(N__33777));
    Span4Mux_h I__7339 (
            .O(N__33816),
            .I(N__33774));
    InMux I__7338 (
            .O(N__33813),
            .I(N__33769));
    InMux I__7337 (
            .O(N__33812),
            .I(N__33769));
    CascadeMux I__7336 (
            .O(N__33811),
            .I(N__33764));
    CascadeMux I__7335 (
            .O(N__33810),
            .I(N__33760));
    CascadeMux I__7334 (
            .O(N__33809),
            .I(N__33757));
    CEMux I__7333 (
            .O(N__33808),
            .I(N__33753));
    InMux I__7332 (
            .O(N__33807),
            .I(N__33744));
    InMux I__7331 (
            .O(N__33804),
            .I(N__33744));
    InMux I__7330 (
            .O(N__33803),
            .I(N__33744));
    InMux I__7329 (
            .O(N__33802),
            .I(N__33744));
    CEMux I__7328 (
            .O(N__33801),
            .I(N__33741));
    Span4Mux_v I__7327 (
            .O(N__33798),
            .I(N__33738));
    CEMux I__7326 (
            .O(N__33797),
            .I(N__33733));
    InMux I__7325 (
            .O(N__33796),
            .I(N__33733));
    InMux I__7324 (
            .O(N__33793),
            .I(N__33719));
    InMux I__7323 (
            .O(N__33790),
            .I(N__33719));
    InMux I__7322 (
            .O(N__33787),
            .I(N__33719));
    InMux I__7321 (
            .O(N__33786),
            .I(N__33719));
    InMux I__7320 (
            .O(N__33783),
            .I(N__33719));
    LocalMux I__7319 (
            .O(N__33780),
            .I(N__33716));
    Span4Mux_v I__7318 (
            .O(N__33777),
            .I(N__33711));
    Span4Mux_h I__7317 (
            .O(N__33774),
            .I(N__33711));
    LocalMux I__7316 (
            .O(N__33769),
            .I(N__33708));
    InMux I__7315 (
            .O(N__33768),
            .I(N__33695));
    CEMux I__7314 (
            .O(N__33767),
            .I(N__33695));
    InMux I__7313 (
            .O(N__33764),
            .I(N__33695));
    InMux I__7312 (
            .O(N__33763),
            .I(N__33695));
    InMux I__7311 (
            .O(N__33760),
            .I(N__33695));
    InMux I__7310 (
            .O(N__33757),
            .I(N__33695));
    CEMux I__7309 (
            .O(N__33756),
            .I(N__33692));
    LocalMux I__7308 (
            .O(N__33753),
            .I(N__33689));
    LocalMux I__7307 (
            .O(N__33744),
            .I(N__33686));
    LocalMux I__7306 (
            .O(N__33741),
            .I(N__33681));
    Span4Mux_h I__7305 (
            .O(N__33738),
            .I(N__33681));
    LocalMux I__7304 (
            .O(N__33733),
            .I(N__33678));
    InMux I__7303 (
            .O(N__33732),
            .I(N__33671));
    InMux I__7302 (
            .O(N__33731),
            .I(N__33671));
    InMux I__7301 (
            .O(N__33730),
            .I(N__33671));
    LocalMux I__7300 (
            .O(N__33719),
            .I(N__33668));
    Span4Mux_s0_h I__7299 (
            .O(N__33716),
            .I(N__33659));
    Span4Mux_v I__7298 (
            .O(N__33711),
            .I(N__33659));
    Span4Mux_h I__7297 (
            .O(N__33708),
            .I(N__33659));
    LocalMux I__7296 (
            .O(N__33695),
            .I(N__33659));
    LocalMux I__7295 (
            .O(N__33692),
            .I(N__33652));
    Span4Mux_h I__7294 (
            .O(N__33689),
            .I(N__33652));
    Span4Mux_h I__7293 (
            .O(N__33686),
            .I(N__33652));
    Odrv4 I__7292 (
            .O(N__33681),
            .I(\b2v_inst11.count_clk_en ));
    Odrv12 I__7291 (
            .O(N__33678),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__7290 (
            .O(N__33671),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__7289 (
            .O(N__33668),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__7288 (
            .O(N__33659),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__7287 (
            .O(N__33652),
            .I(\b2v_inst11.count_clk_en ));
    InMux I__7286 (
            .O(N__33639),
            .I(N__33635));
    InMux I__7285 (
            .O(N__33638),
            .I(N__33632));
    LocalMux I__7284 (
            .O(N__33635),
            .I(N__33626));
    LocalMux I__7283 (
            .O(N__33632),
            .I(N__33626));
    CascadeMux I__7282 (
            .O(N__33631),
            .I(N__33623));
    Span4Mux_h I__7281 (
            .O(N__33626),
            .I(N__33620));
    InMux I__7280 (
            .O(N__33623),
            .I(N__33617));
    Odrv4 I__7279 (
            .O(N__33620),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    LocalMux I__7278 (
            .O(N__33617),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    InMux I__7277 (
            .O(N__33612),
            .I(N__33608));
    InMux I__7276 (
            .O(N__33611),
            .I(N__33605));
    LocalMux I__7275 (
            .O(N__33608),
            .I(N__33602));
    LocalMux I__7274 (
            .O(N__33605),
            .I(N__33599));
    Span4Mux_s3_h I__7273 (
            .O(N__33602),
            .I(N__33596));
    Odrv4 I__7272 (
            .O(N__33599),
            .I(\b2v_inst6.N_241 ));
    Odrv4 I__7271 (
            .O(N__33596),
            .I(\b2v_inst6.N_241 ));
    InMux I__7270 (
            .O(N__33591),
            .I(N__33585));
    CascadeMux I__7269 (
            .O(N__33590),
            .I(N__33582));
    InMux I__7268 (
            .O(N__33589),
            .I(N__33577));
    InMux I__7267 (
            .O(N__33588),
            .I(N__33577));
    LocalMux I__7266 (
            .O(N__33585),
            .I(N__33574));
    InMux I__7265 (
            .O(N__33582),
            .I(N__33571));
    LocalMux I__7264 (
            .O(N__33577),
            .I(N__33568));
    Span4Mux_s2_h I__7263 (
            .O(N__33574),
            .I(N__33565));
    LocalMux I__7262 (
            .O(N__33571),
            .I(N__33560));
    Span4Mux_s1_v I__7261 (
            .O(N__33568),
            .I(N__33560));
    Span4Mux_v I__7260 (
            .O(N__33565),
            .I(N__33557));
    Odrv4 I__7259 (
            .O(N__33560),
            .I(\b2v_inst6.countZ0Z_0 ));
    Odrv4 I__7258 (
            .O(N__33557),
            .I(\b2v_inst6.countZ0Z_0 ));
    InMux I__7257 (
            .O(N__33552),
            .I(N__33546));
    InMux I__7256 (
            .O(N__33551),
            .I(N__33546));
    LocalMux I__7255 (
            .O(N__33546),
            .I(N__33543));
    Span4Mux_s2_v I__7254 (
            .O(N__33543),
            .I(N__33540));
    Span4Mux_v I__7253 (
            .O(N__33540),
            .I(N__33537));
    Odrv4 I__7252 (
            .O(N__33537),
            .I(\b2v_inst6.N_2994_i ));
    CascadeMux I__7251 (
            .O(N__33534),
            .I(\b2v_inst6.N_2994_i_cascade_ ));
    InMux I__7250 (
            .O(N__33531),
            .I(N__33526));
    InMux I__7249 (
            .O(N__33530),
            .I(N__33521));
    InMux I__7248 (
            .O(N__33529),
            .I(N__33521));
    LocalMux I__7247 (
            .O(N__33526),
            .I(N__33518));
    LocalMux I__7246 (
            .O(N__33521),
            .I(N__33515));
    Odrv12 I__7245 (
            .O(N__33518),
            .I(\b2v_inst6.N_389 ));
    Odrv4 I__7244 (
            .O(N__33515),
            .I(\b2v_inst6.N_389 ));
    InMux I__7243 (
            .O(N__33510),
            .I(N__33507));
    LocalMux I__7242 (
            .O(N__33507),
            .I(N__33504));
    Span4Mux_s2_v I__7241 (
            .O(N__33504),
            .I(N__33501));
    Span4Mux_v I__7240 (
            .O(N__33501),
            .I(N__33498));
    Span4Mux_h I__7239 (
            .O(N__33498),
            .I(N__33495));
    Odrv4 I__7238 (
            .O(N__33495),
            .I(\b2v_inst6.count_0_0 ));
    InMux I__7237 (
            .O(N__33492),
            .I(N__33489));
    LocalMux I__7236 (
            .O(N__33489),
            .I(N__33485));
    InMux I__7235 (
            .O(N__33488),
            .I(N__33482));
    Span4Mux_v I__7234 (
            .O(N__33485),
            .I(N__33479));
    LocalMux I__7233 (
            .O(N__33482),
            .I(\b2v_inst6.count_rst ));
    Odrv4 I__7232 (
            .O(N__33479),
            .I(\b2v_inst6.count_rst ));
    InMux I__7231 (
            .O(N__33474),
            .I(N__33471));
    LocalMux I__7230 (
            .O(N__33471),
            .I(N__33468));
    Odrv12 I__7229 (
            .O(N__33468),
            .I(\b2v_inst6.count_0_15 ));
    CascadeMux I__7228 (
            .O(N__33465),
            .I(N__33447));
    InMux I__7227 (
            .O(N__33464),
            .I(N__33438));
    CEMux I__7226 (
            .O(N__33463),
            .I(N__33438));
    InMux I__7225 (
            .O(N__33462),
            .I(N__33435));
    InMux I__7224 (
            .O(N__33461),
            .I(N__33430));
    InMux I__7223 (
            .O(N__33460),
            .I(N__33430));
    InMux I__7222 (
            .O(N__33459),
            .I(N__33427));
    InMux I__7221 (
            .O(N__33458),
            .I(N__33422));
    CEMux I__7220 (
            .O(N__33457),
            .I(N__33422));
    CEMux I__7219 (
            .O(N__33456),
            .I(N__33419));
    CascadeMux I__7218 (
            .O(N__33455),
            .I(N__33414));
    CascadeMux I__7217 (
            .O(N__33454),
            .I(N__33411));
    InMux I__7216 (
            .O(N__33453),
            .I(N__33398));
    InMux I__7215 (
            .O(N__33452),
            .I(N__33398));
    InMux I__7214 (
            .O(N__33451),
            .I(N__33398));
    InMux I__7213 (
            .O(N__33450),
            .I(N__33398));
    InMux I__7212 (
            .O(N__33447),
            .I(N__33389));
    InMux I__7211 (
            .O(N__33446),
            .I(N__33389));
    InMux I__7210 (
            .O(N__33445),
            .I(N__33389));
    CEMux I__7209 (
            .O(N__33444),
            .I(N__33389));
    CascadeMux I__7208 (
            .O(N__33443),
            .I(N__33380));
    LocalMux I__7207 (
            .O(N__33438),
            .I(N__33374));
    LocalMux I__7206 (
            .O(N__33435),
            .I(N__33367));
    LocalMux I__7205 (
            .O(N__33430),
            .I(N__33367));
    LocalMux I__7204 (
            .O(N__33427),
            .I(N__33367));
    LocalMux I__7203 (
            .O(N__33422),
            .I(N__33364));
    LocalMux I__7202 (
            .O(N__33419),
            .I(N__33361));
    CEMux I__7201 (
            .O(N__33418),
            .I(N__33358));
    CEMux I__7200 (
            .O(N__33417),
            .I(N__33355));
    InMux I__7199 (
            .O(N__33414),
            .I(N__33350));
    InMux I__7198 (
            .O(N__33411),
            .I(N__33350));
    InMux I__7197 (
            .O(N__33410),
            .I(N__33347));
    InMux I__7196 (
            .O(N__33409),
            .I(N__33342));
    InMux I__7195 (
            .O(N__33408),
            .I(N__33342));
    CEMux I__7194 (
            .O(N__33407),
            .I(N__33337));
    LocalMux I__7193 (
            .O(N__33398),
            .I(N__33334));
    LocalMux I__7192 (
            .O(N__33389),
            .I(N__33331));
    InMux I__7191 (
            .O(N__33388),
            .I(N__33326));
    InMux I__7190 (
            .O(N__33387),
            .I(N__33326));
    InMux I__7189 (
            .O(N__33386),
            .I(N__33319));
    CEMux I__7188 (
            .O(N__33385),
            .I(N__33319));
    InMux I__7187 (
            .O(N__33384),
            .I(N__33319));
    InMux I__7186 (
            .O(N__33383),
            .I(N__33308));
    InMux I__7185 (
            .O(N__33380),
            .I(N__33308));
    InMux I__7184 (
            .O(N__33379),
            .I(N__33308));
    InMux I__7183 (
            .O(N__33378),
            .I(N__33308));
    InMux I__7182 (
            .O(N__33377),
            .I(N__33308));
    Span4Mux_s2_v I__7181 (
            .O(N__33374),
            .I(N__33305));
    Span4Mux_s2_v I__7180 (
            .O(N__33367),
            .I(N__33302));
    Span4Mux_v I__7179 (
            .O(N__33364),
            .I(N__33297));
    Span4Mux_s2_v I__7178 (
            .O(N__33361),
            .I(N__33297));
    LocalMux I__7177 (
            .O(N__33358),
            .I(N__33288));
    LocalMux I__7176 (
            .O(N__33355),
            .I(N__33288));
    LocalMux I__7175 (
            .O(N__33350),
            .I(N__33288));
    LocalMux I__7174 (
            .O(N__33347),
            .I(N__33288));
    LocalMux I__7173 (
            .O(N__33342),
            .I(N__33285));
    InMux I__7172 (
            .O(N__33341),
            .I(N__33280));
    InMux I__7171 (
            .O(N__33340),
            .I(N__33280));
    LocalMux I__7170 (
            .O(N__33337),
            .I(N__33277));
    Span12Mux_s6_v I__7169 (
            .O(N__33334),
            .I(N__33274));
    Sp12to4 I__7168 (
            .O(N__33331),
            .I(N__33265));
    LocalMux I__7167 (
            .O(N__33326),
            .I(N__33265));
    LocalMux I__7166 (
            .O(N__33319),
            .I(N__33265));
    LocalMux I__7165 (
            .O(N__33308),
            .I(N__33265));
    Span4Mux_v I__7164 (
            .O(N__33305),
            .I(N__33260));
    Span4Mux_v I__7163 (
            .O(N__33302),
            .I(N__33260));
    Span4Mux_h I__7162 (
            .O(N__33297),
            .I(N__33251));
    Span4Mux_s2_v I__7161 (
            .O(N__33288),
            .I(N__33251));
    Span4Mux_s2_v I__7160 (
            .O(N__33285),
            .I(N__33251));
    LocalMux I__7159 (
            .O(N__33280),
            .I(N__33251));
    Odrv4 I__7158 (
            .O(N__33277),
            .I(\b2v_inst6.count_en ));
    Odrv12 I__7157 (
            .O(N__33274),
            .I(\b2v_inst6.count_en ));
    Odrv12 I__7156 (
            .O(N__33265),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7155 (
            .O(N__33260),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7154 (
            .O(N__33251),
            .I(\b2v_inst6.count_en ));
    SRMux I__7153 (
            .O(N__33240),
            .I(N__33232));
    InMux I__7152 (
            .O(N__33239),
            .I(N__33224));
    SRMux I__7151 (
            .O(N__33238),
            .I(N__33224));
    SRMux I__7150 (
            .O(N__33237),
            .I(N__33213));
    SRMux I__7149 (
            .O(N__33236),
            .I(N__33210));
    CascadeMux I__7148 (
            .O(N__33235),
            .I(N__33205));
    LocalMux I__7147 (
            .O(N__33232),
            .I(N__33199));
    CascadeMux I__7146 (
            .O(N__33231),
            .I(N__33192));
    CascadeMux I__7145 (
            .O(N__33230),
            .I(N__33189));
    InMux I__7144 (
            .O(N__33229),
            .I(N__33183));
    LocalMux I__7143 (
            .O(N__33224),
            .I(N__33180));
    InMux I__7142 (
            .O(N__33223),
            .I(N__33175));
    SRMux I__7141 (
            .O(N__33222),
            .I(N__33175));
    InMux I__7140 (
            .O(N__33221),
            .I(N__33164));
    InMux I__7139 (
            .O(N__33220),
            .I(N__33164));
    InMux I__7138 (
            .O(N__33219),
            .I(N__33164));
    InMux I__7137 (
            .O(N__33218),
            .I(N__33164));
    InMux I__7136 (
            .O(N__33217),
            .I(N__33164));
    SRMux I__7135 (
            .O(N__33216),
            .I(N__33152));
    LocalMux I__7134 (
            .O(N__33213),
            .I(N__33147));
    LocalMux I__7133 (
            .O(N__33210),
            .I(N__33147));
    CascadeMux I__7132 (
            .O(N__33209),
            .I(N__33144));
    InMux I__7131 (
            .O(N__33208),
            .I(N__33126));
    InMux I__7130 (
            .O(N__33205),
            .I(N__33126));
    InMux I__7129 (
            .O(N__33204),
            .I(N__33126));
    InMux I__7128 (
            .O(N__33203),
            .I(N__33126));
    InMux I__7127 (
            .O(N__33202),
            .I(N__33126));
    Span4Mux_s2_h I__7126 (
            .O(N__33199),
            .I(N__33123));
    InMux I__7125 (
            .O(N__33198),
            .I(N__33118));
    InMux I__7124 (
            .O(N__33197),
            .I(N__33118));
    SRMux I__7123 (
            .O(N__33196),
            .I(N__33107));
    InMux I__7122 (
            .O(N__33195),
            .I(N__33107));
    InMux I__7121 (
            .O(N__33192),
            .I(N__33107));
    InMux I__7120 (
            .O(N__33189),
            .I(N__33107));
    InMux I__7119 (
            .O(N__33188),
            .I(N__33107));
    InMux I__7118 (
            .O(N__33187),
            .I(N__33102));
    InMux I__7117 (
            .O(N__33186),
            .I(N__33102));
    LocalMux I__7116 (
            .O(N__33183),
            .I(N__33098));
    Span4Mux_v I__7115 (
            .O(N__33180),
            .I(N__33093));
    LocalMux I__7114 (
            .O(N__33175),
            .I(N__33093));
    LocalMux I__7113 (
            .O(N__33164),
            .I(N__33090));
    InMux I__7112 (
            .O(N__33163),
            .I(N__33085));
    InMux I__7111 (
            .O(N__33162),
            .I(N__33085));
    InMux I__7110 (
            .O(N__33161),
            .I(N__33076));
    SRMux I__7109 (
            .O(N__33160),
            .I(N__33076));
    InMux I__7108 (
            .O(N__33159),
            .I(N__33076));
    InMux I__7107 (
            .O(N__33158),
            .I(N__33076));
    InMux I__7106 (
            .O(N__33157),
            .I(N__33069));
    InMux I__7105 (
            .O(N__33156),
            .I(N__33069));
    InMux I__7104 (
            .O(N__33155),
            .I(N__33069));
    LocalMux I__7103 (
            .O(N__33152),
            .I(N__33066));
    Span4Mux_s3_v I__7102 (
            .O(N__33147),
            .I(N__33063));
    InMux I__7101 (
            .O(N__33144),
            .I(N__33054));
    InMux I__7100 (
            .O(N__33143),
            .I(N__33054));
    InMux I__7099 (
            .O(N__33142),
            .I(N__33054));
    InMux I__7098 (
            .O(N__33141),
            .I(N__33054));
    InMux I__7097 (
            .O(N__33140),
            .I(N__33045));
    InMux I__7096 (
            .O(N__33139),
            .I(N__33045));
    InMux I__7095 (
            .O(N__33138),
            .I(N__33045));
    InMux I__7094 (
            .O(N__33137),
            .I(N__33045));
    LocalMux I__7093 (
            .O(N__33126),
            .I(N__33042));
    Span4Mux_s0_v I__7092 (
            .O(N__33123),
            .I(N__33033));
    LocalMux I__7091 (
            .O(N__33118),
            .I(N__33033));
    LocalMux I__7090 (
            .O(N__33107),
            .I(N__33033));
    LocalMux I__7089 (
            .O(N__33102),
            .I(N__33033));
    InMux I__7088 (
            .O(N__33101),
            .I(N__33030));
    Span4Mux_v I__7087 (
            .O(N__33098),
            .I(N__33025));
    Span4Mux_s2_v I__7086 (
            .O(N__33093),
            .I(N__33025));
    Span4Mux_s2_h I__7085 (
            .O(N__33090),
            .I(N__33022));
    LocalMux I__7084 (
            .O(N__33085),
            .I(N__33015));
    LocalMux I__7083 (
            .O(N__33076),
            .I(N__33015));
    LocalMux I__7082 (
            .O(N__33069),
            .I(N__33015));
    Span4Mux_s3_h I__7081 (
            .O(N__33066),
            .I(N__33006));
    Span4Mux_s3_h I__7080 (
            .O(N__33063),
            .I(N__33006));
    LocalMux I__7079 (
            .O(N__33054),
            .I(N__33006));
    LocalMux I__7078 (
            .O(N__33045),
            .I(N__33006));
    Span4Mux_s2_h I__7077 (
            .O(N__33042),
            .I(N__33003));
    Span4Mux_s2_h I__7076 (
            .O(N__33033),
            .I(N__33000));
    LocalMux I__7075 (
            .O(N__33030),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    Odrv4 I__7074 (
            .O(N__33025),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    Odrv4 I__7073 (
            .O(N__33022),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    Odrv12 I__7072 (
            .O(N__33015),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    Odrv4 I__7071 (
            .O(N__33006),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    Odrv4 I__7070 (
            .O(N__33003),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    Odrv4 I__7069 (
            .O(N__33000),
            .I(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ));
    CascadeMux I__7068 (
            .O(N__32985),
            .I(N__32982));
    InMux I__7067 (
            .O(N__32982),
            .I(N__32979));
    LocalMux I__7066 (
            .O(N__32979),
            .I(N__32976));
    Odrv4 I__7065 (
            .O(N__32976),
            .I(\b2v_inst11.func_state_RNI_4Z0Z_1 ));
    InMux I__7064 (
            .O(N__32973),
            .I(N__32970));
    LocalMux I__7063 (
            .O(N__32970),
            .I(\b2v_inst11.un1_count_clk_2_axb_5 ));
    InMux I__7062 (
            .O(N__32967),
            .I(N__32961));
    InMux I__7061 (
            .O(N__32966),
            .I(N__32961));
    LocalMux I__7060 (
            .O(N__32961),
            .I(\b2v_inst11.count_clk_0_5 ));
    InMux I__7059 (
            .O(N__32958),
            .I(N__32949));
    InMux I__7058 (
            .O(N__32957),
            .I(N__32949));
    InMux I__7057 (
            .O(N__32956),
            .I(N__32949));
    LocalMux I__7056 (
            .O(N__32949),
            .I(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ));
    CascadeMux I__7055 (
            .O(N__32946),
            .I(N__32941));
    InMux I__7054 (
            .O(N__32945),
            .I(N__32934));
    InMux I__7053 (
            .O(N__32944),
            .I(N__32934));
    InMux I__7052 (
            .O(N__32941),
            .I(N__32934));
    LocalMux I__7051 (
            .O(N__32934),
            .I(N__32931));
    Odrv12 I__7050 (
            .O(N__32931),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    InMux I__7049 (
            .O(N__32928),
            .I(N__32925));
    LocalMux I__7048 (
            .O(N__32925),
            .I(N__32921));
    InMux I__7047 (
            .O(N__32924),
            .I(N__32918));
    Span4Mux_s1_h I__7046 (
            .O(N__32921),
            .I(N__32915));
    LocalMux I__7045 (
            .O(N__32918),
            .I(\b2v_inst11.count_clk_0_7 ));
    Odrv4 I__7044 (
            .O(N__32915),
            .I(\b2v_inst11.count_clk_0_7 ));
    InMux I__7043 (
            .O(N__32910),
            .I(N__32904));
    InMux I__7042 (
            .O(N__32909),
            .I(N__32904));
    LocalMux I__7041 (
            .O(N__32904),
            .I(N__32900));
    InMux I__7040 (
            .O(N__32903),
            .I(N__32897));
    Odrv4 I__7039 (
            .O(N__32900),
            .I(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ));
    LocalMux I__7038 (
            .O(N__32897),
            .I(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ));
    CascadeMux I__7037 (
            .O(N__32892),
            .I(N__32889));
    InMux I__7036 (
            .O(N__32889),
            .I(N__32886));
    LocalMux I__7035 (
            .O(N__32886),
            .I(\b2v_inst11.un1_count_clk_2_axb_7 ));
    CascadeMux I__7034 (
            .O(N__32883),
            .I(N__32880));
    InMux I__7033 (
            .O(N__32880),
            .I(N__32874));
    InMux I__7032 (
            .O(N__32879),
            .I(N__32874));
    LocalMux I__7031 (
            .O(N__32874),
            .I(N__32870));
    CascadeMux I__7030 (
            .O(N__32873),
            .I(N__32867));
    Span4Mux_v I__7029 (
            .O(N__32870),
            .I(N__32864));
    InMux I__7028 (
            .O(N__32867),
            .I(N__32861));
    Odrv4 I__7027 (
            .O(N__32864),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    LocalMux I__7026 (
            .O(N__32861),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    InMux I__7025 (
            .O(N__32856),
            .I(N__32850));
    InMux I__7024 (
            .O(N__32855),
            .I(N__32850));
    LocalMux I__7023 (
            .O(N__32850),
            .I(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ));
    InMux I__7022 (
            .O(N__32847),
            .I(N__32844));
    LocalMux I__7021 (
            .O(N__32844),
            .I(\b2v_inst11.count_clk_0_4 ));
    CascadeMux I__7020 (
            .O(N__32841),
            .I(N__32838));
    InMux I__7019 (
            .O(N__32838),
            .I(N__32835));
    LocalMux I__7018 (
            .O(N__32835),
            .I(\b2v_inst11.un1_count_clk_2_axb_2 ));
    InMux I__7017 (
            .O(N__32832),
            .I(N__32826));
    InMux I__7016 (
            .O(N__32831),
            .I(N__32826));
    LocalMux I__7015 (
            .O(N__32826),
            .I(\b2v_inst11.count_clk_0_2 ));
    InMux I__7014 (
            .O(N__32823),
            .I(N__32814));
    InMux I__7013 (
            .O(N__32822),
            .I(N__32814));
    InMux I__7012 (
            .O(N__32821),
            .I(N__32814));
    LocalMux I__7011 (
            .O(N__32814),
            .I(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ));
    InMux I__7010 (
            .O(N__32811),
            .I(N__32805));
    InMux I__7009 (
            .O(N__32810),
            .I(N__32805));
    LocalMux I__7008 (
            .O(N__32805),
            .I(N__32802));
    Span4Mux_v I__7007 (
            .O(N__32802),
            .I(N__32799));
    Odrv4 I__7006 (
            .O(N__32799),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    CascadeMux I__7005 (
            .O(N__32796),
            .I(N__32792));
    InMux I__7004 (
            .O(N__32795),
            .I(N__32784));
    InMux I__7003 (
            .O(N__32792),
            .I(N__32784));
    InMux I__7002 (
            .O(N__32791),
            .I(N__32784));
    LocalMux I__7001 (
            .O(N__32784),
            .I(\b2v_inst6.un2_count_1_cry_9_c_RNIVIZ0Z14 ));
    InMux I__7000 (
            .O(N__32781),
            .I(N__32778));
    LocalMux I__6999 (
            .O(N__32778),
            .I(\b2v_inst6.count_rst_4 ));
    CascadeMux I__6998 (
            .O(N__32775),
            .I(N__32772));
    InMux I__6997 (
            .O(N__32772),
            .I(N__32769));
    LocalMux I__6996 (
            .O(N__32769),
            .I(\b2v_inst6.countZ0Z_15 ));
    CascadeMux I__6995 (
            .O(N__32766),
            .I(N__32763));
    InMux I__6994 (
            .O(N__32763),
            .I(N__32759));
    InMux I__6993 (
            .O(N__32762),
            .I(N__32756));
    LocalMux I__6992 (
            .O(N__32759),
            .I(\b2v_inst6.count_0_13 ));
    LocalMux I__6991 (
            .O(N__32756),
            .I(\b2v_inst6.count_0_13 ));
    CascadeMux I__6990 (
            .O(N__32751),
            .I(\b2v_inst6.countZ0Z_15_cascade_ ));
    InMux I__6989 (
            .O(N__32748),
            .I(N__32745));
    LocalMux I__6988 (
            .O(N__32745),
            .I(N__32742));
    Odrv4 I__6987 (
            .O(N__32742),
            .I(\b2v_inst6.count_1_i_a3_2_0 ));
    CascadeMux I__6986 (
            .O(N__32739),
            .I(N__32735));
    InMux I__6985 (
            .O(N__32738),
            .I(N__32729));
    InMux I__6984 (
            .O(N__32735),
            .I(N__32729));
    InMux I__6983 (
            .O(N__32734),
            .I(N__32726));
    LocalMux I__6982 (
            .O(N__32729),
            .I(\b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0 ));
    LocalMux I__6981 (
            .O(N__32726),
            .I(\b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0 ));
    InMux I__6980 (
            .O(N__32721),
            .I(N__32718));
    LocalMux I__6979 (
            .O(N__32718),
            .I(\b2v_inst6.count_rst_1 ));
    InMux I__6978 (
            .O(N__32715),
            .I(N__32712));
    LocalMux I__6977 (
            .O(N__32712),
            .I(\b2v_inst11.un1_count_clk_2_axb_12 ));
    CascadeMux I__6976 (
            .O(N__32709),
            .I(N__32706));
    InMux I__6975 (
            .O(N__32706),
            .I(N__32703));
    LocalMux I__6974 (
            .O(N__32703),
            .I(N__32698));
    InMux I__6973 (
            .O(N__32702),
            .I(N__32693));
    InMux I__6972 (
            .O(N__32701),
            .I(N__32693));
    Odrv4 I__6971 (
            .O(N__32698),
            .I(\b2v_inst11.count_clk_1_12 ));
    LocalMux I__6970 (
            .O(N__32693),
            .I(\b2v_inst11.count_clk_1_12 ));
    InMux I__6969 (
            .O(N__32688),
            .I(N__32684));
    InMux I__6968 (
            .O(N__32687),
            .I(N__32681));
    LocalMux I__6967 (
            .O(N__32684),
            .I(\b2v_inst11.count_clk_0_12 ));
    LocalMux I__6966 (
            .O(N__32681),
            .I(\b2v_inst11.count_clk_0_12 ));
    InMux I__6965 (
            .O(N__32676),
            .I(N__32673));
    LocalMux I__6964 (
            .O(N__32673),
            .I(\b2v_inst11.un1_count_clk_2_axb_13 ));
    InMux I__6963 (
            .O(N__32670),
            .I(N__32667));
    LocalMux I__6962 (
            .O(N__32667),
            .I(N__32662));
    InMux I__6961 (
            .O(N__32666),
            .I(N__32657));
    InMux I__6960 (
            .O(N__32665),
            .I(N__32657));
    Odrv4 I__6959 (
            .O(N__32662),
            .I(\b2v_inst11.count_clk_1_13 ));
    LocalMux I__6958 (
            .O(N__32657),
            .I(\b2v_inst11.count_clk_1_13 ));
    InMux I__6957 (
            .O(N__32652),
            .I(N__32648));
    InMux I__6956 (
            .O(N__32651),
            .I(N__32645));
    LocalMux I__6955 (
            .O(N__32648),
            .I(\b2v_inst11.count_clk_0_13 ));
    LocalMux I__6954 (
            .O(N__32645),
            .I(\b2v_inst11.count_clk_0_13 ));
    CascadeMux I__6953 (
            .O(N__32640),
            .I(\b2v_inst6.countZ0Z_6_cascade_ ));
    CascadeMux I__6952 (
            .O(N__32637),
            .I(\b2v_inst6.count_1_i_a3_0_0_cascade_ ));
    InMux I__6951 (
            .O(N__32634),
            .I(N__32631));
    LocalMux I__6950 (
            .O(N__32631),
            .I(\b2v_inst6.count_1_i_a3_7_0 ));
    InMux I__6949 (
            .O(N__32628),
            .I(N__32622));
    InMux I__6948 (
            .O(N__32627),
            .I(N__32622));
    LocalMux I__6947 (
            .O(N__32622),
            .I(\b2v_inst6.count_0_6 ));
    InMux I__6946 (
            .O(N__32619),
            .I(N__32615));
    CascadeMux I__6945 (
            .O(N__32618),
            .I(N__32612));
    LocalMux I__6944 (
            .O(N__32615),
            .I(N__32608));
    InMux I__6943 (
            .O(N__32612),
            .I(N__32603));
    InMux I__6942 (
            .O(N__32611),
            .I(N__32603));
    Odrv4 I__6941 (
            .O(N__32608),
            .I(\b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ));
    LocalMux I__6940 (
            .O(N__32603),
            .I(\b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ));
    CascadeMux I__6939 (
            .O(N__32598),
            .I(N__32595));
    InMux I__6938 (
            .O(N__32595),
            .I(N__32592));
    LocalMux I__6937 (
            .O(N__32592),
            .I(\b2v_inst6.un2_count_1_axb_6 ));
    InMux I__6936 (
            .O(N__32589),
            .I(N__32586));
    LocalMux I__6935 (
            .O(N__32586),
            .I(\b2v_inst6.count_rst_2 ));
    CascadeMux I__6934 (
            .O(N__32583),
            .I(N__32579));
    InMux I__6933 (
            .O(N__32582),
            .I(N__32574));
    InMux I__6932 (
            .O(N__32579),
            .I(N__32574));
    LocalMux I__6931 (
            .O(N__32574),
            .I(\b2v_inst6.count_0_12 ));
    InMux I__6930 (
            .O(N__32571),
            .I(N__32562));
    InMux I__6929 (
            .O(N__32570),
            .I(N__32562));
    InMux I__6928 (
            .O(N__32569),
            .I(N__32562));
    LocalMux I__6927 (
            .O(N__32562),
            .I(\b2v_inst6.un2_count_1_cry_11_c_RNI8RABZ0 ));
    InMux I__6926 (
            .O(N__32559),
            .I(N__32556));
    LocalMux I__6925 (
            .O(N__32556),
            .I(\b2v_inst6.un2_count_1_axb_12 ));
    InMux I__6924 (
            .O(N__32553),
            .I(N__32550));
    LocalMux I__6923 (
            .O(N__32550),
            .I(\b2v_inst6.un2_count_1_axb_10 ));
    InMux I__6922 (
            .O(N__32547),
            .I(N__32543));
    InMux I__6921 (
            .O(N__32546),
            .I(N__32540));
    LocalMux I__6920 (
            .O(N__32543),
            .I(\b2v_inst6.count_0_10 ));
    LocalMux I__6919 (
            .O(N__32540),
            .I(\b2v_inst6.count_0_10 ));
    InMux I__6918 (
            .O(N__32535),
            .I(N__32529));
    InMux I__6917 (
            .O(N__32534),
            .I(N__32529));
    LocalMux I__6916 (
            .O(N__32529),
            .I(\b2v_inst6.count_0_14 ));
    InMux I__6915 (
            .O(N__32526),
            .I(N__32517));
    InMux I__6914 (
            .O(N__32525),
            .I(N__32517));
    InMux I__6913 (
            .O(N__32524),
            .I(N__32517));
    LocalMux I__6912 (
            .O(N__32517),
            .I(\b2v_inst6.un2_count_1_cry_13_c_RNIR6IOZ0Z5 ));
    CascadeMux I__6911 (
            .O(N__32514),
            .I(N__32511));
    InMux I__6910 (
            .O(N__32511),
            .I(N__32508));
    LocalMux I__6909 (
            .O(N__32508),
            .I(\b2v_inst6.un2_count_1_axb_14 ));
    InMux I__6908 (
            .O(N__32505),
            .I(N__32502));
    LocalMux I__6907 (
            .O(N__32502),
            .I(\b2v_inst6.countZ0Z_14 ));
    CascadeMux I__6906 (
            .O(N__32499),
            .I(\b2v_inst6.count_rst_12_cascade_ ));
    InMux I__6905 (
            .O(N__32496),
            .I(N__32493));
    LocalMux I__6904 (
            .O(N__32493),
            .I(N__32490));
    Odrv4 I__6903 (
            .O(N__32490),
            .I(\b2v_inst6.count_1_i_a3_12_0 ));
    CascadeMux I__6902 (
            .O(N__32487),
            .I(\b2v_inst6.count_1_i_a3_1_0_cascade_ ));
    InMux I__6901 (
            .O(N__32484),
            .I(N__32478));
    InMux I__6900 (
            .O(N__32483),
            .I(N__32478));
    LocalMux I__6899 (
            .O(N__32478),
            .I(\b2v_inst6.count_0_2 ));
    CascadeMux I__6898 (
            .O(N__32475),
            .I(N__32471));
    InMux I__6897 (
            .O(N__32474),
            .I(N__32463));
    InMux I__6896 (
            .O(N__32471),
            .I(N__32463));
    InMux I__6895 (
            .O(N__32470),
            .I(N__32463));
    LocalMux I__6894 (
            .O(N__32463),
            .I(\b2v_inst6.un2_count_1_cry_1_c_RNIN2PZ0Z3 ));
    InMux I__6893 (
            .O(N__32460),
            .I(N__32457));
    LocalMux I__6892 (
            .O(N__32457),
            .I(\b2v_inst6.un2_count_1_axb_2 ));
    InMux I__6891 (
            .O(N__32454),
            .I(N__32451));
    LocalMux I__6890 (
            .O(N__32451),
            .I(\b2v_inst6.count_rst_7 ));
    InMux I__6889 (
            .O(N__32448),
            .I(N__32444));
    InMux I__6888 (
            .O(N__32447),
            .I(N__32441));
    LocalMux I__6887 (
            .O(N__32444),
            .I(\b2v_inst6.count_0_7 ));
    LocalMux I__6886 (
            .O(N__32441),
            .I(\b2v_inst6.count_0_7 ));
    CascadeMux I__6885 (
            .O(N__32436),
            .I(\b2v_inst6.countZ0Z_5_cascade_ ));
    CascadeMux I__6884 (
            .O(N__32433),
            .I(\b2v_inst6.count_RNICV5H1Z0Z_1_cascade_ ));
    InMux I__6883 (
            .O(N__32430),
            .I(N__32426));
    InMux I__6882 (
            .O(N__32429),
            .I(N__32423));
    LocalMux I__6881 (
            .O(N__32426),
            .I(\b2v_inst6.un2_count_1_axb_1 ));
    LocalMux I__6880 (
            .O(N__32423),
            .I(\b2v_inst6.un2_count_1_axb_1 ));
    CascadeMux I__6879 (
            .O(N__32418),
            .I(\b2v_inst6.un2_count_1_axb_1_cascade_ ));
    InMux I__6878 (
            .O(N__32415),
            .I(N__32412));
    LocalMux I__6877 (
            .O(N__32412),
            .I(\b2v_inst6.count_RNICV5H1Z0Z_1 ));
    CascadeMux I__6876 (
            .O(N__32409),
            .I(N__32405));
    InMux I__6875 (
            .O(N__32408),
            .I(N__32401));
    InMux I__6874 (
            .O(N__32405),
            .I(N__32398));
    InMux I__6873 (
            .O(N__32404),
            .I(N__32395));
    LocalMux I__6872 (
            .O(N__32401),
            .I(N__32392));
    LocalMux I__6871 (
            .O(N__32398),
            .I(\b2v_inst6.countZ0Z_11 ));
    LocalMux I__6870 (
            .O(N__32395),
            .I(\b2v_inst6.countZ0Z_11 ));
    Odrv4 I__6869 (
            .O(N__32392),
            .I(\b2v_inst6.countZ0Z_11 ));
    InMux I__6868 (
            .O(N__32385),
            .I(N__32379));
    InMux I__6867 (
            .O(N__32384),
            .I(N__32379));
    LocalMux I__6866 (
            .O(N__32379),
            .I(\b2v_inst6.count_0_1 ));
    InMux I__6865 (
            .O(N__32376),
            .I(N__32373));
    LocalMux I__6864 (
            .O(N__32373),
            .I(N__32370));
    Odrv12 I__6863 (
            .O(N__32370),
            .I(\b2v_inst6.count_1_i_a3_4_0 ));
    InMux I__6862 (
            .O(N__32367),
            .I(N__32364));
    LocalMux I__6861 (
            .O(N__32364),
            .I(N__32361));
    Odrv12 I__6860 (
            .O(N__32361),
            .I(\b2v_inst6.count_1_i_a3_6_0 ));
    CascadeMux I__6859 (
            .O(N__32358),
            .I(\b2v_inst6.count_1_i_a3_3_0_cascade_ ));
    InMux I__6858 (
            .O(N__32355),
            .I(N__32352));
    LocalMux I__6857 (
            .O(N__32352),
            .I(\b2v_inst6.count_1_i_a3_5_0 ));
    InMux I__6856 (
            .O(N__32349),
            .I(N__32343));
    InMux I__6855 (
            .O(N__32348),
            .I(N__32343));
    LocalMux I__6854 (
            .O(N__32343),
            .I(\b2v_inst6.count_0_5 ));
    InMux I__6853 (
            .O(N__32340),
            .I(N__32334));
    InMux I__6852 (
            .O(N__32339),
            .I(N__32334));
    LocalMux I__6851 (
            .O(N__32334),
            .I(\b2v_inst6.count_rst_9 ));
    CascadeMux I__6850 (
            .O(N__32331),
            .I(N__32327));
    CascadeMux I__6849 (
            .O(N__32330),
            .I(N__32324));
    InMux I__6848 (
            .O(N__32327),
            .I(N__32318));
    InMux I__6847 (
            .O(N__32324),
            .I(N__32318));
    InMux I__6846 (
            .O(N__32323),
            .I(N__32315));
    LocalMux I__6845 (
            .O(N__32318),
            .I(\b2v_inst6.un2_count_1_axb_5 ));
    LocalMux I__6844 (
            .O(N__32315),
            .I(\b2v_inst6.un2_count_1_axb_5 ));
    InMux I__6843 (
            .O(N__32310),
            .I(N__32298));
    InMux I__6842 (
            .O(N__32309),
            .I(N__32289));
    InMux I__6841 (
            .O(N__32308),
            .I(N__32286));
    CascadeMux I__6840 (
            .O(N__32307),
            .I(N__32279));
    InMux I__6839 (
            .O(N__32306),
            .I(N__32270));
    InMux I__6838 (
            .O(N__32305),
            .I(N__32263));
    InMux I__6837 (
            .O(N__32304),
            .I(N__32260));
    InMux I__6836 (
            .O(N__32303),
            .I(N__32253));
    InMux I__6835 (
            .O(N__32302),
            .I(N__32253));
    InMux I__6834 (
            .O(N__32301),
            .I(N__32253));
    LocalMux I__6833 (
            .O(N__32298),
            .I(N__32250));
    InMux I__6832 (
            .O(N__32297),
            .I(N__32243));
    InMux I__6831 (
            .O(N__32296),
            .I(N__32243));
    InMux I__6830 (
            .O(N__32295),
            .I(N__32234));
    InMux I__6829 (
            .O(N__32294),
            .I(N__32234));
    InMux I__6828 (
            .O(N__32293),
            .I(N__32234));
    InMux I__6827 (
            .O(N__32292),
            .I(N__32234));
    LocalMux I__6826 (
            .O(N__32289),
            .I(N__32229));
    LocalMux I__6825 (
            .O(N__32286),
            .I(N__32229));
    InMux I__6824 (
            .O(N__32285),
            .I(N__32226));
    InMux I__6823 (
            .O(N__32284),
            .I(N__32217));
    InMux I__6822 (
            .O(N__32283),
            .I(N__32217));
    InMux I__6821 (
            .O(N__32282),
            .I(N__32217));
    InMux I__6820 (
            .O(N__32279),
            .I(N__32217));
    CascadeMux I__6819 (
            .O(N__32278),
            .I(N__32214));
    InMux I__6818 (
            .O(N__32277),
            .I(N__32205));
    InMux I__6817 (
            .O(N__32276),
            .I(N__32205));
    InMux I__6816 (
            .O(N__32275),
            .I(N__32205));
    InMux I__6815 (
            .O(N__32274),
            .I(N__32205));
    CascadeMux I__6814 (
            .O(N__32273),
            .I(N__32200));
    LocalMux I__6813 (
            .O(N__32270),
            .I(N__32193));
    InMux I__6812 (
            .O(N__32269),
            .I(N__32186));
    InMux I__6811 (
            .O(N__32268),
            .I(N__32186));
    InMux I__6810 (
            .O(N__32267),
            .I(N__32186));
    InMux I__6809 (
            .O(N__32266),
            .I(N__32177));
    LocalMux I__6808 (
            .O(N__32263),
            .I(N__32174));
    LocalMux I__6807 (
            .O(N__32260),
            .I(N__32167));
    LocalMux I__6806 (
            .O(N__32253),
            .I(N__32167));
    Span4Mux_v I__6805 (
            .O(N__32250),
            .I(N__32167));
    InMux I__6804 (
            .O(N__32249),
            .I(N__32164));
    InMux I__6803 (
            .O(N__32248),
            .I(N__32160));
    LocalMux I__6802 (
            .O(N__32243),
            .I(N__32157));
    LocalMux I__6801 (
            .O(N__32234),
            .I(N__32148));
    Span4Mux_v I__6800 (
            .O(N__32229),
            .I(N__32148));
    LocalMux I__6799 (
            .O(N__32226),
            .I(N__32148));
    LocalMux I__6798 (
            .O(N__32217),
            .I(N__32148));
    InMux I__6797 (
            .O(N__32214),
            .I(N__32143));
    LocalMux I__6796 (
            .O(N__32205),
            .I(N__32140));
    InMux I__6795 (
            .O(N__32204),
            .I(N__32125));
    InMux I__6794 (
            .O(N__32203),
            .I(N__32125));
    InMux I__6793 (
            .O(N__32200),
            .I(N__32125));
    InMux I__6792 (
            .O(N__32199),
            .I(N__32125));
    InMux I__6791 (
            .O(N__32198),
            .I(N__32125));
    InMux I__6790 (
            .O(N__32197),
            .I(N__32125));
    InMux I__6789 (
            .O(N__32196),
            .I(N__32125));
    Span4Mux_v I__6788 (
            .O(N__32193),
            .I(N__32120));
    LocalMux I__6787 (
            .O(N__32186),
            .I(N__32120));
    InMux I__6786 (
            .O(N__32185),
            .I(N__32107));
    InMux I__6785 (
            .O(N__32184),
            .I(N__32107));
    InMux I__6784 (
            .O(N__32183),
            .I(N__32107));
    InMux I__6783 (
            .O(N__32182),
            .I(N__32107));
    InMux I__6782 (
            .O(N__32181),
            .I(N__32107));
    InMux I__6781 (
            .O(N__32180),
            .I(N__32107));
    LocalMux I__6780 (
            .O(N__32177),
            .I(N__32104));
    Span4Mux_v I__6779 (
            .O(N__32174),
            .I(N__32097));
    Span4Mux_v I__6778 (
            .O(N__32167),
            .I(N__32097));
    LocalMux I__6777 (
            .O(N__32164),
            .I(N__32097));
    InMux I__6776 (
            .O(N__32163),
            .I(N__32094));
    LocalMux I__6775 (
            .O(N__32160),
            .I(N__32087));
    Span4Mux_v I__6774 (
            .O(N__32157),
            .I(N__32087));
    Span4Mux_v I__6773 (
            .O(N__32148),
            .I(N__32087));
    InMux I__6772 (
            .O(N__32147),
            .I(N__32082));
    InMux I__6771 (
            .O(N__32146),
            .I(N__32082));
    LocalMux I__6770 (
            .O(N__32143),
            .I(N__32073));
    Span4Mux_h I__6769 (
            .O(N__32140),
            .I(N__32073));
    LocalMux I__6768 (
            .O(N__32125),
            .I(N__32073));
    Span4Mux_h I__6767 (
            .O(N__32120),
            .I(N__32073));
    LocalMux I__6766 (
            .O(N__32107),
            .I(N__32070));
    Odrv12 I__6765 (
            .O(N__32104),
            .I(\b2v_inst11.N_2904_i ));
    Odrv4 I__6764 (
            .O(N__32097),
            .I(\b2v_inst11.N_2904_i ));
    LocalMux I__6763 (
            .O(N__32094),
            .I(\b2v_inst11.N_2904_i ));
    Odrv4 I__6762 (
            .O(N__32087),
            .I(\b2v_inst11.N_2904_i ));
    LocalMux I__6761 (
            .O(N__32082),
            .I(\b2v_inst11.N_2904_i ));
    Odrv4 I__6760 (
            .O(N__32073),
            .I(\b2v_inst11.N_2904_i ));
    Odrv12 I__6759 (
            .O(N__32070),
            .I(\b2v_inst11.N_2904_i ));
    CascadeMux I__6758 (
            .O(N__32055),
            .I(N__32052));
    InMux I__6757 (
            .O(N__32052),
            .I(N__32049));
    LocalMux I__6756 (
            .O(N__32049),
            .I(N__32046));
    Span12Mux_s1_h I__6755 (
            .O(N__32046),
            .I(N__32043));
    Odrv12 I__6754 (
            .O(N__32043),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_12 ));
    InMux I__6753 (
            .O(N__32040),
            .I(N__32037));
    LocalMux I__6752 (
            .O(N__32037),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_7 ));
    CascadeMux I__6751 (
            .O(N__32034),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ));
    CascadeMux I__6750 (
            .O(N__32031),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_9_cascade_ ));
    CascadeMux I__6749 (
            .O(N__32028),
            .I(N__32025));
    InMux I__6748 (
            .O(N__32025),
            .I(N__32022));
    LocalMux I__6747 (
            .O(N__32022),
            .I(N__32019));
    Span4Mux_v I__6746 (
            .O(N__32019),
            .I(N__32016));
    Odrv4 I__6745 (
            .O(N__32016),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_10 ));
    InMux I__6744 (
            .O(N__32013),
            .I(N__32010));
    LocalMux I__6743 (
            .O(N__32010),
            .I(N__32007));
    Span4Mux_v I__6742 (
            .O(N__32007),
            .I(N__32004));
    Odrv4 I__6741 (
            .O(N__32004),
            .I(\b2v_inst11.un1_dutycycle_94_s1_9 ));
    InMux I__6740 (
            .O(N__32001),
            .I(N__31998));
    LocalMux I__6739 (
            .O(N__31998),
            .I(N__31995));
    Odrv4 I__6738 (
            .O(N__31995),
            .I(\b2v_inst11.un1_dutycycle_94_s0_9 ));
    CascadeMux I__6737 (
            .O(N__31992),
            .I(\b2v_inst11.i2_mux_cascade_ ));
    CascadeMux I__6736 (
            .O(N__31989),
            .I(N__31980));
    InMux I__6735 (
            .O(N__31988),
            .I(N__31977));
    InMux I__6734 (
            .O(N__31987),
            .I(N__31974));
    InMux I__6733 (
            .O(N__31986),
            .I(N__31971));
    InMux I__6732 (
            .O(N__31985),
            .I(N__31966));
    CascadeMux I__6731 (
            .O(N__31984),
            .I(N__31962));
    InMux I__6730 (
            .O(N__31983),
            .I(N__31958));
    InMux I__6729 (
            .O(N__31980),
            .I(N__31955));
    LocalMux I__6728 (
            .O(N__31977),
            .I(N__31952));
    LocalMux I__6727 (
            .O(N__31974),
            .I(N__31949));
    LocalMux I__6726 (
            .O(N__31971),
            .I(N__31945));
    InMux I__6725 (
            .O(N__31970),
            .I(N__31942));
    InMux I__6724 (
            .O(N__31969),
            .I(N__31939));
    LocalMux I__6723 (
            .O(N__31966),
            .I(N__31936));
    InMux I__6722 (
            .O(N__31965),
            .I(N__31929));
    InMux I__6721 (
            .O(N__31962),
            .I(N__31929));
    InMux I__6720 (
            .O(N__31961),
            .I(N__31929));
    LocalMux I__6719 (
            .O(N__31958),
            .I(N__31926));
    LocalMux I__6718 (
            .O(N__31955),
            .I(N__31923));
    Span4Mux_v I__6717 (
            .O(N__31952),
            .I(N__31920));
    Span4Mux_h I__6716 (
            .O(N__31949),
            .I(N__31917));
    InMux I__6715 (
            .O(N__31948),
            .I(N__31914));
    Span4Mux_s3_h I__6714 (
            .O(N__31945),
            .I(N__31903));
    LocalMux I__6713 (
            .O(N__31942),
            .I(N__31903));
    LocalMux I__6712 (
            .O(N__31939),
            .I(N__31903));
    Span4Mux_s1_v I__6711 (
            .O(N__31936),
            .I(N__31903));
    LocalMux I__6710 (
            .O(N__31929),
            .I(N__31903));
    Span4Mux_s2_h I__6709 (
            .O(N__31926),
            .I(N__31898));
    Span4Mux_s2_h I__6708 (
            .O(N__31923),
            .I(N__31898));
    Odrv4 I__6707 (
            .O(N__31920),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__6706 (
            .O(N__31917),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__6705 (
            .O(N__31914),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__6704 (
            .O(N__31903),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__6703 (
            .O(N__31898),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    CascadeMux I__6702 (
            .O(N__31887),
            .I(\b2v_inst11.un1_N_5_cascade_ ));
    InMux I__6701 (
            .O(N__31884),
            .I(N__31880));
    InMux I__6700 (
            .O(N__31883),
            .I(N__31877));
    LocalMux I__6699 (
            .O(N__31880),
            .I(\b2v_inst11.un1_i2_mux_0_0 ));
    LocalMux I__6698 (
            .O(N__31877),
            .I(\b2v_inst11.un1_i2_mux_0_0 ));
    CascadeMux I__6697 (
            .O(N__31872),
            .I(N__31869));
    InMux I__6696 (
            .O(N__31869),
            .I(N__31866));
    LocalMux I__6695 (
            .O(N__31866),
            .I(N__31863));
    Span4Mux_h I__6694 (
            .O(N__31863),
            .I(N__31860));
    Odrv4 I__6693 (
            .O(N__31860),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_11 ));
    CascadeMux I__6692 (
            .O(N__31857),
            .I(N__31854));
    InMux I__6691 (
            .O(N__31854),
            .I(N__31851));
    LocalMux I__6690 (
            .O(N__31851),
            .I(N__31848));
    Odrv4 I__6689 (
            .O(N__31848),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_14 ));
    InMux I__6688 (
            .O(N__31845),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_s0 ));
    InMux I__6687 (
            .O(N__31842),
            .I(N__31839));
    LocalMux I__6686 (
            .O(N__31839),
            .I(N__31836));
    Span4Mux_s3_v I__6685 (
            .O(N__31836),
            .I(N__31833));
    Odrv4 I__6684 (
            .O(N__31833),
            .I(\b2v_inst11.un1_dutycycle_94_axb_15_s0 ));
    InMux I__6683 (
            .O(N__31830),
            .I(N__31827));
    LocalMux I__6682 (
            .O(N__31827),
            .I(N__31824));
    Odrv12 I__6681 (
            .O(N__31824),
            .I(\b2v_inst11.un1_dutycycle_94_s1_15 ));
    InMux I__6680 (
            .O(N__31821),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14_s0 ));
    InMux I__6679 (
            .O(N__31818),
            .I(N__31815));
    LocalMux I__6678 (
            .O(N__31815),
            .I(N__31812));
    Odrv4 I__6677 (
            .O(N__31812),
            .I(\b2v_inst11.un1_dutycycle_53_axb_12_1 ));
    CascadeMux I__6676 (
            .O(N__31809),
            .I(N__31806));
    InMux I__6675 (
            .O(N__31806),
            .I(N__31803));
    LocalMux I__6674 (
            .O(N__31803),
            .I(N__31800));
    Odrv4 I__6673 (
            .O(N__31800),
            .I(\b2v_inst11.un1_dutycycle_53_3_1 ));
    CascadeMux I__6672 (
            .O(N__31797),
            .I(\b2v_inst11.un1_dutycycle_53_31_cascade_ ));
    InMux I__6671 (
            .O(N__31794),
            .I(N__31791));
    LocalMux I__6670 (
            .O(N__31791),
            .I(N__31788));
    Odrv4 I__6669 (
            .O(N__31788),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_13 ));
    InMux I__6668 (
            .O(N__31785),
            .I(N__31782));
    LocalMux I__6667 (
            .O(N__31782),
            .I(\b2v_inst11.un1_dutycycle_53_31 ));
    InMux I__6666 (
            .O(N__31779),
            .I(N__31773));
    InMux I__6665 (
            .O(N__31778),
            .I(N__31773));
    LocalMux I__6664 (
            .O(N__31773),
            .I(N__31770));
    Span12Mux_s3_h I__6663 (
            .O(N__31770),
            .I(N__31767));
    Odrv12 I__6662 (
            .O(N__31767),
            .I(\b2v_inst11.un1_dutycycle_53_55_0_tz ));
    CascadeMux I__6661 (
            .O(N__31764),
            .I(\b2v_inst11.un1_dutycycle_53_axb_14_1_cascade_ ));
    CascadeMux I__6660 (
            .O(N__31761),
            .I(\b2v_inst11.un1_dutycycle_53_axb_14_cascade_ ));
    CascadeMux I__6659 (
            .O(N__31758),
            .I(N__31755));
    InMux I__6658 (
            .O(N__31755),
            .I(N__31752));
    LocalMux I__6657 (
            .O(N__31752),
            .I(N__31749));
    Odrv4 I__6656 (
            .O(N__31749),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_14 ));
    InMux I__6655 (
            .O(N__31746),
            .I(N__31743));
    LocalMux I__6654 (
            .O(N__31743),
            .I(N__31740));
    Span4Mux_h I__6653 (
            .O(N__31740),
            .I(N__31737));
    Odrv4 I__6652 (
            .O(N__31737),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_9 ));
    CascadeMux I__6651 (
            .O(N__31734),
            .I(N__31731));
    InMux I__6650 (
            .O(N__31731),
            .I(N__31728));
    LocalMux I__6649 (
            .O(N__31728),
            .I(N__31725));
    Odrv4 I__6648 (
            .O(N__31725),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_6 ));
    InMux I__6647 (
            .O(N__31722),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_s0 ));
    InMux I__6646 (
            .O(N__31719),
            .I(N__31716));
    LocalMux I__6645 (
            .O(N__31716),
            .I(\b2v_inst11.dutycycle_RNI_10Z0Z_7 ));
    InMux I__6644 (
            .O(N__31713),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_s0 ));
    InMux I__6643 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__6642 (
            .O(N__31707),
            .I(N__31704));
    Span4Mux_h I__6641 (
            .O(N__31704),
            .I(N__31701));
    Odrv4 I__6640 (
            .O(N__31701),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_8 ));
    InMux I__6639 (
            .O(N__31698),
            .I(bfn_11_14_0_));
    InMux I__6638 (
            .O(N__31695),
            .I(N__31692));
    LocalMux I__6637 (
            .O(N__31692),
            .I(N__31689));
    Odrv4 I__6636 (
            .O(N__31689),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_9 ));
    InMux I__6635 (
            .O(N__31686),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_s0 ));
    InMux I__6634 (
            .O(N__31683),
            .I(N__31680));
    LocalMux I__6633 (
            .O(N__31680),
            .I(N__31677));
    Odrv12 I__6632 (
            .O(N__31677),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_10 ));
    InMux I__6631 (
            .O(N__31674),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_s0 ));
    InMux I__6630 (
            .O(N__31671),
            .I(N__31668));
    LocalMux I__6629 (
            .O(N__31668),
            .I(N__31665));
    Span4Mux_s1_h I__6628 (
            .O(N__31665),
            .I(N__31662));
    Odrv4 I__6627 (
            .O(N__31662),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_11 ));
    InMux I__6626 (
            .O(N__31659),
            .I(N__31656));
    LocalMux I__6625 (
            .O(N__31656),
            .I(N__31653));
    Odrv4 I__6624 (
            .O(N__31653),
            .I(\b2v_inst11.un1_dutycycle_94_s0_11 ));
    InMux I__6623 (
            .O(N__31650),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10_s0 ));
    InMux I__6622 (
            .O(N__31647),
            .I(N__31644));
    LocalMux I__6621 (
            .O(N__31644),
            .I(N__31641));
    Odrv4 I__6620 (
            .O(N__31641),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_12 ));
    InMux I__6619 (
            .O(N__31638),
            .I(N__31635));
    LocalMux I__6618 (
            .O(N__31635),
            .I(N__31632));
    Odrv4 I__6617 (
            .O(N__31632),
            .I(\b2v_inst11.un1_dutycycle_94_s0_12 ));
    InMux I__6616 (
            .O(N__31629),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11_s0 ));
    CascadeMux I__6615 (
            .O(N__31626),
            .I(N__31623));
    InMux I__6614 (
            .O(N__31623),
            .I(N__31620));
    LocalMux I__6613 (
            .O(N__31620),
            .I(N__31617));
    Span4Mux_s1_h I__6612 (
            .O(N__31617),
            .I(N__31614));
    Odrv4 I__6611 (
            .O(N__31614),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_13 ));
    InMux I__6610 (
            .O(N__31611),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_s0 ));
    InMux I__6609 (
            .O(N__31608),
            .I(N__31605));
    LocalMux I__6608 (
            .O(N__31605),
            .I(N__31602));
    Odrv4 I__6607 (
            .O(N__31602),
            .I(\b2v_inst11.un1_dutycycle_94_s1_11 ));
    InMux I__6606 (
            .O(N__31599),
            .I(N__31593));
    InMux I__6605 (
            .O(N__31598),
            .I(N__31593));
    LocalMux I__6604 (
            .O(N__31593),
            .I(N__31590));
    Span4Mux_h I__6603 (
            .O(N__31590),
            .I(N__31587));
    Odrv4 I__6602 (
            .O(N__31587),
            .I(\b2v_inst11.dutycycle_rst_6 ));
    InMux I__6601 (
            .O(N__31584),
            .I(N__31578));
    CascadeMux I__6600 (
            .O(N__31583),
            .I(N__31574));
    InMux I__6599 (
            .O(N__31582),
            .I(N__31571));
    CascadeMux I__6598 (
            .O(N__31581),
            .I(N__31567));
    LocalMux I__6597 (
            .O(N__31578),
            .I(N__31564));
    InMux I__6596 (
            .O(N__31577),
            .I(N__31559));
    InMux I__6595 (
            .O(N__31574),
            .I(N__31559));
    LocalMux I__6594 (
            .O(N__31571),
            .I(N__31549));
    InMux I__6593 (
            .O(N__31570),
            .I(N__31544));
    InMux I__6592 (
            .O(N__31567),
            .I(N__31544));
    Span4Mux_s2_h I__6591 (
            .O(N__31564),
            .I(N__31541));
    LocalMux I__6590 (
            .O(N__31559),
            .I(N__31538));
    InMux I__6589 (
            .O(N__31558),
            .I(N__31535));
    CascadeMux I__6588 (
            .O(N__31557),
            .I(N__31529));
    CascadeMux I__6587 (
            .O(N__31556),
            .I(N__31524));
    InMux I__6586 (
            .O(N__31555),
            .I(N__31515));
    InMux I__6585 (
            .O(N__31554),
            .I(N__31515));
    InMux I__6584 (
            .O(N__31553),
            .I(N__31515));
    InMux I__6583 (
            .O(N__31552),
            .I(N__31515));
    Span4Mux_v I__6582 (
            .O(N__31549),
            .I(N__31512));
    LocalMux I__6581 (
            .O(N__31544),
            .I(N__31509));
    Span4Mux_v I__6580 (
            .O(N__31541),
            .I(N__31506));
    Span12Mux_s7_v I__6579 (
            .O(N__31538),
            .I(N__31501));
    LocalMux I__6578 (
            .O(N__31535),
            .I(N__31501));
    InMux I__6577 (
            .O(N__31534),
            .I(N__31494));
    InMux I__6576 (
            .O(N__31533),
            .I(N__31494));
    InMux I__6575 (
            .O(N__31532),
            .I(N__31494));
    InMux I__6574 (
            .O(N__31529),
            .I(N__31489));
    InMux I__6573 (
            .O(N__31528),
            .I(N__31489));
    InMux I__6572 (
            .O(N__31527),
            .I(N__31484));
    InMux I__6571 (
            .O(N__31524),
            .I(N__31484));
    LocalMux I__6570 (
            .O(N__31515),
            .I(N__31477));
    Span4Mux_h I__6569 (
            .O(N__31512),
            .I(N__31477));
    Span4Mux_v I__6568 (
            .O(N__31509),
            .I(N__31477));
    Odrv4 I__6567 (
            .O(N__31506),
            .I(\b2v_inst11.dutycycle ));
    Odrv12 I__6566 (
            .O(N__31501),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__6565 (
            .O(N__31494),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__6564 (
            .O(N__31489),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__6563 (
            .O(N__31484),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__6562 (
            .O(N__31477),
            .I(\b2v_inst11.dutycycle ));
    InMux I__6561 (
            .O(N__31464),
            .I(N__31457));
    InMux I__6560 (
            .O(N__31463),
            .I(N__31450));
    CascadeMux I__6559 (
            .O(N__31462),
            .I(N__31445));
    InMux I__6558 (
            .O(N__31461),
            .I(N__31435));
    InMux I__6557 (
            .O(N__31460),
            .I(N__31435));
    LocalMux I__6556 (
            .O(N__31457),
            .I(N__31432));
    InMux I__6555 (
            .O(N__31456),
            .I(N__31429));
    CascadeMux I__6554 (
            .O(N__31455),
            .I(N__31426));
    InMux I__6553 (
            .O(N__31454),
            .I(N__31418));
    InMux I__6552 (
            .O(N__31453),
            .I(N__31418));
    LocalMux I__6551 (
            .O(N__31450),
            .I(N__31415));
    InMux I__6550 (
            .O(N__31449),
            .I(N__31406));
    InMux I__6549 (
            .O(N__31448),
            .I(N__31406));
    InMux I__6548 (
            .O(N__31445),
            .I(N__31406));
    InMux I__6547 (
            .O(N__31444),
            .I(N__31406));
    InMux I__6546 (
            .O(N__31443),
            .I(N__31399));
    InMux I__6545 (
            .O(N__31442),
            .I(N__31399));
    InMux I__6544 (
            .O(N__31441),
            .I(N__31399));
    CascadeMux I__6543 (
            .O(N__31440),
            .I(N__31396));
    LocalMux I__6542 (
            .O(N__31435),
            .I(N__31390));
    Span4Mux_v I__6541 (
            .O(N__31432),
            .I(N__31385));
    LocalMux I__6540 (
            .O(N__31429),
            .I(N__31385));
    InMux I__6539 (
            .O(N__31426),
            .I(N__31382));
    InMux I__6538 (
            .O(N__31425),
            .I(N__31375));
    InMux I__6537 (
            .O(N__31424),
            .I(N__31375));
    InMux I__6536 (
            .O(N__31423),
            .I(N__31375));
    LocalMux I__6535 (
            .O(N__31418),
            .I(N__31366));
    Span4Mux_v I__6534 (
            .O(N__31415),
            .I(N__31366));
    LocalMux I__6533 (
            .O(N__31406),
            .I(N__31366));
    LocalMux I__6532 (
            .O(N__31399),
            .I(N__31366));
    InMux I__6531 (
            .O(N__31396),
            .I(N__31363));
    InMux I__6530 (
            .O(N__31395),
            .I(N__31360));
    InMux I__6529 (
            .O(N__31394),
            .I(N__31355));
    InMux I__6528 (
            .O(N__31393),
            .I(N__31355));
    Span4Mux_h I__6527 (
            .O(N__31390),
            .I(N__31352));
    Span4Mux_v I__6526 (
            .O(N__31385),
            .I(N__31341));
    LocalMux I__6525 (
            .O(N__31382),
            .I(N__31341));
    LocalMux I__6524 (
            .O(N__31375),
            .I(N__31341));
    Span4Mux_v I__6523 (
            .O(N__31366),
            .I(N__31341));
    LocalMux I__6522 (
            .O(N__31363),
            .I(N__31341));
    LocalMux I__6521 (
            .O(N__31360),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    LocalMux I__6520 (
            .O(N__31355),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv4 I__6519 (
            .O(N__31352),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv4 I__6518 (
            .O(N__31341),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    CascadeMux I__6517 (
            .O(N__31332),
            .I(N__31329));
    InMux I__6516 (
            .O(N__31329),
            .I(N__31326));
    LocalMux I__6515 (
            .O(N__31326),
            .I(N__31323));
    Odrv12 I__6514 (
            .O(N__31323),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_1 ));
    InMux I__6513 (
            .O(N__31320),
            .I(N__31317));
    LocalMux I__6512 (
            .O(N__31317),
            .I(N__31314));
    Span4Mux_h I__6511 (
            .O(N__31314),
            .I(N__31311));
    Span4Mux_v I__6510 (
            .O(N__31311),
            .I(N__31308));
    Odrv4 I__6509 (
            .O(N__31308),
            .I(\b2v_inst11.un1_dutycycle_94_s0_1 ));
    InMux I__6508 (
            .O(N__31305),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_s0 ));
    CascadeMux I__6507 (
            .O(N__31302),
            .I(N__31292));
    CascadeMux I__6506 (
            .O(N__31301),
            .I(N__31286));
    InMux I__6505 (
            .O(N__31300),
            .I(N__31283));
    InMux I__6504 (
            .O(N__31299),
            .I(N__31280));
    InMux I__6503 (
            .O(N__31298),
            .I(N__31277));
    InMux I__6502 (
            .O(N__31297),
            .I(N__31274));
    InMux I__6501 (
            .O(N__31296),
            .I(N__31271));
    InMux I__6500 (
            .O(N__31295),
            .I(N__31268));
    InMux I__6499 (
            .O(N__31292),
            .I(N__31265));
    CascadeMux I__6498 (
            .O(N__31291),
            .I(N__31262));
    CascadeMux I__6497 (
            .O(N__31290),
            .I(N__31259));
    InMux I__6496 (
            .O(N__31289),
            .I(N__31252));
    InMux I__6495 (
            .O(N__31286),
            .I(N__31252));
    LocalMux I__6494 (
            .O(N__31283),
            .I(N__31249));
    LocalMux I__6493 (
            .O(N__31280),
            .I(N__31246));
    LocalMux I__6492 (
            .O(N__31277),
            .I(N__31243));
    LocalMux I__6491 (
            .O(N__31274),
            .I(N__31236));
    LocalMux I__6490 (
            .O(N__31271),
            .I(N__31236));
    LocalMux I__6489 (
            .O(N__31268),
            .I(N__31236));
    LocalMux I__6488 (
            .O(N__31265),
            .I(N__31233));
    InMux I__6487 (
            .O(N__31262),
            .I(N__31230));
    InMux I__6486 (
            .O(N__31259),
            .I(N__31227));
    InMux I__6485 (
            .O(N__31258),
            .I(N__31222));
    InMux I__6484 (
            .O(N__31257),
            .I(N__31222));
    LocalMux I__6483 (
            .O(N__31252),
            .I(N__31219));
    Span4Mux_v I__6482 (
            .O(N__31249),
            .I(N__31210));
    Span4Mux_v I__6481 (
            .O(N__31246),
            .I(N__31210));
    Span4Mux_v I__6480 (
            .O(N__31243),
            .I(N__31210));
    Span4Mux_v I__6479 (
            .O(N__31236),
            .I(N__31210));
    Span4Mux_h I__6478 (
            .O(N__31233),
            .I(N__31207));
    LocalMux I__6477 (
            .O(N__31230),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__6476 (
            .O(N__31227),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__6475 (
            .O(N__31222),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__6474 (
            .O(N__31219),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__6473 (
            .O(N__31210),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__6472 (
            .O(N__31207),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    CascadeMux I__6471 (
            .O(N__31194),
            .I(N__31191));
    InMux I__6470 (
            .O(N__31191),
            .I(N__31188));
    LocalMux I__6469 (
            .O(N__31188),
            .I(N__31185));
    Span4Mux_s2_h I__6468 (
            .O(N__31185),
            .I(N__31182));
    Odrv4 I__6467 (
            .O(N__31182),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_2 ));
    InMux I__6466 (
            .O(N__31179),
            .I(N__31176));
    LocalMux I__6465 (
            .O(N__31176),
            .I(N__31173));
    Span4Mux_v I__6464 (
            .O(N__31173),
            .I(N__31170));
    Span4Mux_h I__6463 (
            .O(N__31170),
            .I(N__31167));
    Odrv4 I__6462 (
            .O(N__31167),
            .I(\b2v_inst11.un1_dutycycle_94_s0_2 ));
    InMux I__6461 (
            .O(N__31164),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_s0 ));
    CascadeMux I__6460 (
            .O(N__31161),
            .I(N__31158));
    InMux I__6459 (
            .O(N__31158),
            .I(N__31155));
    LocalMux I__6458 (
            .O(N__31155),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_3 ));
    InMux I__6457 (
            .O(N__31152),
            .I(N__31149));
    LocalMux I__6456 (
            .O(N__31149),
            .I(N__31146));
    Odrv4 I__6455 (
            .O(N__31146),
            .I(\b2v_inst11.un1_dutycycle_94_s0_3 ));
    InMux I__6454 (
            .O(N__31143),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2_s0 ));
    CascadeMux I__6453 (
            .O(N__31140),
            .I(N__31137));
    InMux I__6452 (
            .O(N__31137),
            .I(N__31134));
    LocalMux I__6451 (
            .O(N__31134),
            .I(N__31131));
    Odrv12 I__6450 (
            .O(N__31131),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_4 ));
    InMux I__6449 (
            .O(N__31128),
            .I(N__31125));
    LocalMux I__6448 (
            .O(N__31125),
            .I(N__31122));
    Span4Mux_h I__6447 (
            .O(N__31122),
            .I(N__31119));
    Odrv4 I__6446 (
            .O(N__31119),
            .I(\b2v_inst11.un1_dutycycle_94_s0_4 ));
    InMux I__6445 (
            .O(N__31116),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3_s0 ));
    InMux I__6444 (
            .O(N__31113),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4_s0 ));
    InMux I__6443 (
            .O(N__31110),
            .I(N__31107));
    LocalMux I__6442 (
            .O(N__31107),
            .I(N__31104));
    Odrv4 I__6441 (
            .O(N__31104),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_3 ));
    CascadeMux I__6440 (
            .O(N__31101),
            .I(N__31098));
    InMux I__6439 (
            .O(N__31098),
            .I(N__31095));
    LocalMux I__6438 (
            .O(N__31095),
            .I(N__31092));
    Odrv4 I__6437 (
            .O(N__31092),
            .I(\b2v_inst11.un1_dutycycle_94_s1_12 ));
    InMux I__6436 (
            .O(N__31089),
            .I(N__31085));
    InMux I__6435 (
            .O(N__31088),
            .I(N__31082));
    LocalMux I__6434 (
            .O(N__31085),
            .I(N__31077));
    LocalMux I__6433 (
            .O(N__31082),
            .I(N__31077));
    Odrv4 I__6432 (
            .O(N__31077),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EGZ0Z1 ));
    InMux I__6431 (
            .O(N__31074),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10_s1 ));
    InMux I__6430 (
            .O(N__31071),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11_s1 ));
    CascadeMux I__6429 (
            .O(N__31068),
            .I(N__31065));
    InMux I__6428 (
            .O(N__31065),
            .I(N__31062));
    LocalMux I__6427 (
            .O(N__31062),
            .I(N__31059));
    Span4Mux_s3_h I__6426 (
            .O(N__31059),
            .I(N__31056));
    Odrv4 I__6425 (
            .O(N__31056),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ));
    InMux I__6424 (
            .O(N__31053),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_s1 ));
    CascadeMux I__6423 (
            .O(N__31050),
            .I(N__31047));
    InMux I__6422 (
            .O(N__31047),
            .I(N__31044));
    LocalMux I__6421 (
            .O(N__31044),
            .I(N__31041));
    Span4Mux_s2_h I__6420 (
            .O(N__31041),
            .I(N__31038));
    Odrv4 I__6419 (
            .O(N__31038),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_14 ));
    InMux I__6418 (
            .O(N__31035),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_s1 ));
    InMux I__6417 (
            .O(N__31032),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14_s1 ));
    CascadeMux I__6416 (
            .O(N__31029),
            .I(N__31026));
    InMux I__6415 (
            .O(N__31026),
            .I(N__31023));
    LocalMux I__6414 (
            .O(N__31023),
            .I(N__31020));
    Odrv4 I__6413 (
            .O(N__31020),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_6 ));
    CascadeMux I__6412 (
            .O(N__31017),
            .I(N__31014));
    InMux I__6411 (
            .O(N__31014),
            .I(N__31011));
    LocalMux I__6410 (
            .O(N__31011),
            .I(N__31008));
    Odrv4 I__6409 (
            .O(N__31008),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_11 ));
    InMux I__6408 (
            .O(N__31005),
            .I(N__31002));
    LocalMux I__6407 (
            .O(N__31002),
            .I(N__30999));
    Odrv12 I__6406 (
            .O(N__30999),
            .I(\b2v_inst11.un1_dutycycle_94_s1_3 ));
    CascadeMux I__6405 (
            .O(N__30996),
            .I(N__30993));
    InMux I__6404 (
            .O(N__30993),
            .I(N__30990));
    LocalMux I__6403 (
            .O(N__30990),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_8 ));
    InMux I__6402 (
            .O(N__30987),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_s1 ));
    InMux I__6401 (
            .O(N__30984),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2_s1 ));
    CascadeMux I__6400 (
            .O(N__30981),
            .I(N__30978));
    InMux I__6399 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__6398 (
            .O(N__30975),
            .I(N__30972));
    Odrv4 I__6397 (
            .O(N__30972),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_4 ));
    InMux I__6396 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__6395 (
            .O(N__30966),
            .I(N__30963));
    Span4Mux_h I__6394 (
            .O(N__30963),
            .I(N__30960));
    Span4Mux_v I__6393 (
            .O(N__30960),
            .I(N__30957));
    Odrv4 I__6392 (
            .O(N__30957),
            .I(\b2v_inst11.un1_dutycycle_94_s1_4 ));
    InMux I__6391 (
            .O(N__30954),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3_s1 ));
    InMux I__6390 (
            .O(N__30951),
            .I(N__30948));
    LocalMux I__6389 (
            .O(N__30948),
            .I(N__30942));
    InMux I__6388 (
            .O(N__30947),
            .I(N__30939));
    InMux I__6387 (
            .O(N__30946),
            .I(N__30936));
    IoInMux I__6386 (
            .O(N__30945),
            .I(N__30933));
    Span4Mux_v I__6385 (
            .O(N__30942),
            .I(N__30930));
    LocalMux I__6384 (
            .O(N__30939),
            .I(N__30925));
    LocalMux I__6383 (
            .O(N__30936),
            .I(N__30925));
    LocalMux I__6382 (
            .O(N__30933),
            .I(N__30922));
    Span4Mux_h I__6381 (
            .O(N__30930),
            .I(N__30917));
    Span4Mux_v I__6380 (
            .O(N__30925),
            .I(N__30917));
    Span4Mux_s1_h I__6379 (
            .O(N__30922),
            .I(N__30914));
    Sp12to4 I__6378 (
            .O(N__30917),
            .I(N__30911));
    Span4Mux_v I__6377 (
            .O(N__30914),
            .I(N__30908));
    Odrv12 I__6376 (
            .O(N__30911),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6375 (
            .O(N__30908),
            .I(CONSTANT_ONE_NET));
    InMux I__6374 (
            .O(N__30903),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4_s1 ));
    InMux I__6373 (
            .O(N__30900),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_s1 ));
    CascadeMux I__6372 (
            .O(N__30897),
            .I(N__30894));
    InMux I__6371 (
            .O(N__30894),
            .I(N__30891));
    LocalMux I__6370 (
            .O(N__30891),
            .I(N__30888));
    Span4Mux_s2_h I__6369 (
            .O(N__30888),
            .I(N__30885));
    Odrv4 I__6368 (
            .O(N__30885),
            .I(\b2v_inst11.dutycycle_RNI_9Z0Z_7 ));
    InMux I__6367 (
            .O(N__30882),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_s1 ));
    InMux I__6366 (
            .O(N__30879),
            .I(bfn_11_10_0_));
    CascadeMux I__6365 (
            .O(N__30876),
            .I(N__30873));
    InMux I__6364 (
            .O(N__30873),
            .I(N__30870));
    LocalMux I__6363 (
            .O(N__30870),
            .I(N__30867));
    Odrv12 I__6362 (
            .O(N__30867),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_9 ));
    InMux I__6361 (
            .O(N__30864),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_s1 ));
    InMux I__6360 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__6359 (
            .O(N__30858),
            .I(N__30855));
    Odrv12 I__6358 (
            .O(N__30855),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_10 ));
    InMux I__6357 (
            .O(N__30852),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_s1 ));
    CascadeMux I__6356 (
            .O(N__30849),
            .I(\b2v_inst11.count_clk_en_cascade_ ));
    InMux I__6355 (
            .O(N__30846),
            .I(N__30842));
    InMux I__6354 (
            .O(N__30845),
            .I(N__30839));
    LocalMux I__6353 (
            .O(N__30842),
            .I(N__30836));
    LocalMux I__6352 (
            .O(N__30839),
            .I(N__30833));
    Odrv12 I__6351 (
            .O(N__30836),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    Odrv4 I__6350 (
            .O(N__30833),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    CascadeMux I__6349 (
            .O(N__30828),
            .I(N__30825));
    InMux I__6348 (
            .O(N__30825),
            .I(N__30821));
    InMux I__6347 (
            .O(N__30824),
            .I(N__30818));
    LocalMux I__6346 (
            .O(N__30821),
            .I(N__30815));
    LocalMux I__6345 (
            .O(N__30818),
            .I(N__30812));
    Span4Mux_s3_h I__6344 (
            .O(N__30815),
            .I(N__30809));
    Span4Mux_v I__6343 (
            .O(N__30812),
            .I(N__30806));
    Odrv4 I__6342 (
            .O(N__30809),
            .I(\b2v_inst11.N_417 ));
    Odrv4 I__6341 (
            .O(N__30806),
            .I(\b2v_inst11.N_417 ));
    CascadeMux I__6340 (
            .O(N__30801),
            .I(N__30796));
    CascadeMux I__6339 (
            .O(N__30800),
            .I(N__30793));
    InMux I__6338 (
            .O(N__30799),
            .I(N__30783));
    InMux I__6337 (
            .O(N__30796),
            .I(N__30783));
    InMux I__6336 (
            .O(N__30793),
            .I(N__30783));
    InMux I__6335 (
            .O(N__30792),
            .I(N__30783));
    LocalMux I__6334 (
            .O(N__30783),
            .I(N__30779));
    InMux I__6333 (
            .O(N__30782),
            .I(N__30776));
    Odrv12 I__6332 (
            .O(N__30779),
            .I(\b2v_inst11.func_state_RNID7Q51Z0Z_0 ));
    LocalMux I__6331 (
            .O(N__30776),
            .I(\b2v_inst11.func_state_RNID7Q51Z0Z_0 ));
    InMux I__6330 (
            .O(N__30771),
            .I(N__30762));
    InMux I__6329 (
            .O(N__30770),
            .I(N__30762));
    CascadeMux I__6328 (
            .O(N__30769),
            .I(N__30758));
    CascadeMux I__6327 (
            .O(N__30768),
            .I(N__30755));
    InMux I__6326 (
            .O(N__30767),
            .I(N__30750));
    LocalMux I__6325 (
            .O(N__30762),
            .I(N__30744));
    InMux I__6324 (
            .O(N__30761),
            .I(N__30741));
    InMux I__6323 (
            .O(N__30758),
            .I(N__30732));
    InMux I__6322 (
            .O(N__30755),
            .I(N__30732));
    InMux I__6321 (
            .O(N__30754),
            .I(N__30732));
    InMux I__6320 (
            .O(N__30753),
            .I(N__30732));
    LocalMux I__6319 (
            .O(N__30750),
            .I(N__30729));
    InMux I__6318 (
            .O(N__30749),
            .I(N__30722));
    InMux I__6317 (
            .O(N__30748),
            .I(N__30722));
    InMux I__6316 (
            .O(N__30747),
            .I(N__30722));
    Span4Mux_v I__6315 (
            .O(N__30744),
            .I(N__30719));
    LocalMux I__6314 (
            .O(N__30741),
            .I(N__30714));
    LocalMux I__6313 (
            .O(N__30732),
            .I(N__30714));
    Odrv12 I__6312 (
            .O(N__30729),
            .I(\b2v_inst11.count_off_RNI_1Z0Z_1 ));
    LocalMux I__6311 (
            .O(N__30722),
            .I(\b2v_inst11.count_off_RNI_1Z0Z_1 ));
    Odrv4 I__6310 (
            .O(N__30719),
            .I(\b2v_inst11.count_off_RNI_1Z0Z_1 ));
    Odrv4 I__6309 (
            .O(N__30714),
            .I(\b2v_inst11.count_off_RNI_1Z0Z_1 ));
    InMux I__6308 (
            .O(N__30705),
            .I(N__30702));
    LocalMux I__6307 (
            .O(N__30702),
            .I(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0 ));
    InMux I__6306 (
            .O(N__30699),
            .I(N__30693));
    InMux I__6305 (
            .O(N__30698),
            .I(N__30693));
    LocalMux I__6304 (
            .O(N__30693),
            .I(N__30690));
    Odrv12 I__6303 (
            .O(N__30690),
            .I(\b2v_inst11.func_state_RNI6M5R2Z0Z_1 ));
    CascadeMux I__6302 (
            .O(N__30687),
            .I(N__30684));
    InMux I__6301 (
            .O(N__30684),
            .I(N__30672));
    InMux I__6300 (
            .O(N__30683),
            .I(N__30672));
    InMux I__6299 (
            .O(N__30682),
            .I(N__30672));
    InMux I__6298 (
            .O(N__30681),
            .I(N__30672));
    LocalMux I__6297 (
            .O(N__30672),
            .I(N__30669));
    Span4Mux_s1_h I__6296 (
            .O(N__30669),
            .I(N__30666));
    Odrv4 I__6295 (
            .O(N__30666),
            .I(\b2v_inst11.func_state_RNIJGA54Z0Z_1 ));
    InMux I__6294 (
            .O(N__30663),
            .I(N__30657));
    InMux I__6293 (
            .O(N__30662),
            .I(N__30657));
    LocalMux I__6292 (
            .O(N__30657),
            .I(N__30654));
    Odrv4 I__6291 (
            .O(N__30654),
            .I(\b2v_inst11.count_clk_1_14 ));
    InMux I__6290 (
            .O(N__30651),
            .I(N__30648));
    LocalMux I__6289 (
            .O(N__30648),
            .I(\b2v_inst11.count_clk_0_14 ));
    InMux I__6288 (
            .O(N__30645),
            .I(N__30638));
    InMux I__6287 (
            .O(N__30644),
            .I(N__30638));
    CascadeMux I__6286 (
            .O(N__30643),
            .I(N__30630));
    LocalMux I__6285 (
            .O(N__30638),
            .I(N__30624));
    InMux I__6284 (
            .O(N__30637),
            .I(N__30621));
    InMux I__6283 (
            .O(N__30636),
            .I(N__30616));
    InMux I__6282 (
            .O(N__30635),
            .I(N__30616));
    InMux I__6281 (
            .O(N__30634),
            .I(N__30613));
    InMux I__6280 (
            .O(N__30633),
            .I(N__30610));
    InMux I__6279 (
            .O(N__30630),
            .I(N__30605));
    InMux I__6278 (
            .O(N__30629),
            .I(N__30605));
    InMux I__6277 (
            .O(N__30628),
            .I(N__30600));
    InMux I__6276 (
            .O(N__30627),
            .I(N__30600));
    Span4Mux_h I__6275 (
            .O(N__30624),
            .I(N__30595));
    LocalMux I__6274 (
            .O(N__30621),
            .I(N__30595));
    LocalMux I__6273 (
            .O(N__30616),
            .I(N__30592));
    LocalMux I__6272 (
            .O(N__30613),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__6271 (
            .O(N__30610),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__6270 (
            .O(N__30605),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__6269 (
            .O(N__30600),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    Odrv4 I__6268 (
            .O(N__30595),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    Odrv4 I__6267 (
            .O(N__30592),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    CascadeMux I__6266 (
            .O(N__30579),
            .I(\b2v_inst11.N_2904_i_cascade_ ));
    InMux I__6265 (
            .O(N__30576),
            .I(N__30573));
    LocalMux I__6264 (
            .O(N__30573),
            .I(N__30570));
    Span4Mux_v I__6263 (
            .O(N__30570),
            .I(N__30567));
    Span4Mux_h I__6262 (
            .O(N__30567),
            .I(N__30564));
    Odrv4 I__6261 (
            .O(N__30564),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_1 ));
    InMux I__6260 (
            .O(N__30561),
            .I(N__30558));
    LocalMux I__6259 (
            .O(N__30558),
            .I(N__30555));
    Odrv4 I__6258 (
            .O(N__30555),
            .I(\b2v_inst11.un1_dutycycle_94_s1_1 ));
    InMux I__6257 (
            .O(N__30552),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_s1 ));
    CascadeMux I__6256 (
            .O(N__30549),
            .I(N__30546));
    InMux I__6255 (
            .O(N__30546),
            .I(N__30543));
    LocalMux I__6254 (
            .O(N__30543),
            .I(N__30540));
    Span4Mux_s2_h I__6253 (
            .O(N__30540),
            .I(N__30537));
    Odrv4 I__6252 (
            .O(N__30537),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_2 ));
    InMux I__6251 (
            .O(N__30534),
            .I(N__30531));
    LocalMux I__6250 (
            .O(N__30531),
            .I(N__30528));
    Span4Mux_h I__6249 (
            .O(N__30528),
            .I(N__30525));
    Odrv4 I__6248 (
            .O(N__30525),
            .I(\b2v_inst11.un1_dutycycle_94_s1_2 ));
    InMux I__6247 (
            .O(N__30522),
            .I(N__30515));
    InMux I__6246 (
            .O(N__30521),
            .I(N__30515));
    InMux I__6245 (
            .O(N__30520),
            .I(N__30512));
    LocalMux I__6244 (
            .O(N__30515),
            .I(N__30509));
    LocalMux I__6243 (
            .O(N__30512),
            .I(N__30506));
    Span4Mux_v I__6242 (
            .O(N__30509),
            .I(N__30503));
    Odrv4 I__6241 (
            .O(N__30506),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    Odrv4 I__6240 (
            .O(N__30503),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    InMux I__6239 (
            .O(N__30498),
            .I(N__30492));
    InMux I__6238 (
            .O(N__30497),
            .I(N__30492));
    LocalMux I__6237 (
            .O(N__30492),
            .I(N__30489));
    Odrv4 I__6236 (
            .O(N__30489),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ));
    InMux I__6235 (
            .O(N__30486),
            .I(N__30483));
    LocalMux I__6234 (
            .O(N__30483),
            .I(\b2v_inst11.count_clk_0_8 ));
    InMux I__6233 (
            .O(N__30480),
            .I(N__30471));
    InMux I__6232 (
            .O(N__30479),
            .I(N__30471));
    InMux I__6231 (
            .O(N__30478),
            .I(N__30471));
    LocalMux I__6230 (
            .O(N__30471),
            .I(N__30467));
    InMux I__6229 (
            .O(N__30470),
            .I(N__30464));
    Span4Mux_h I__6228 (
            .O(N__30467),
            .I(N__30461));
    LocalMux I__6227 (
            .O(N__30464),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    Odrv4 I__6226 (
            .O(N__30461),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    InMux I__6225 (
            .O(N__30456),
            .I(N__30450));
    InMux I__6224 (
            .O(N__30455),
            .I(N__30450));
    LocalMux I__6223 (
            .O(N__30450),
            .I(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ));
    InMux I__6222 (
            .O(N__30447),
            .I(N__30444));
    LocalMux I__6221 (
            .O(N__30444),
            .I(\b2v_inst11.count_clk_0_9 ));
    InMux I__6220 (
            .O(N__30441),
            .I(N__30431));
    InMux I__6219 (
            .O(N__30440),
            .I(N__30431));
    InMux I__6218 (
            .O(N__30439),
            .I(N__30425));
    InMux I__6217 (
            .O(N__30438),
            .I(N__30422));
    InMux I__6216 (
            .O(N__30437),
            .I(N__30417));
    InMux I__6215 (
            .O(N__30436),
            .I(N__30417));
    LocalMux I__6214 (
            .O(N__30431),
            .I(N__30414));
    InMux I__6213 (
            .O(N__30430),
            .I(N__30411));
    InMux I__6212 (
            .O(N__30429),
            .I(N__30406));
    InMux I__6211 (
            .O(N__30428),
            .I(N__30406));
    LocalMux I__6210 (
            .O(N__30425),
            .I(N__30403));
    LocalMux I__6209 (
            .O(N__30422),
            .I(N__30392));
    LocalMux I__6208 (
            .O(N__30417),
            .I(N__30392));
    Span4Mux_v I__6207 (
            .O(N__30414),
            .I(N__30392));
    LocalMux I__6206 (
            .O(N__30411),
            .I(N__30392));
    LocalMux I__6205 (
            .O(N__30406),
            .I(N__30392));
    Span4Mux_v I__6204 (
            .O(N__30403),
            .I(N__30389));
    Span4Mux_v I__6203 (
            .O(N__30392),
            .I(N__30386));
    Odrv4 I__6202 (
            .O(N__30389),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__6201 (
            .O(N__30386),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    CascadeMux I__6200 (
            .O(N__30381),
            .I(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0_cascade_ ));
    InMux I__6199 (
            .O(N__30378),
            .I(N__30374));
    CascadeMux I__6198 (
            .O(N__30377),
            .I(N__30371));
    LocalMux I__6197 (
            .O(N__30374),
            .I(N__30367));
    InMux I__6196 (
            .O(N__30371),
            .I(N__30364));
    InMux I__6195 (
            .O(N__30370),
            .I(N__30361));
    Span4Mux_s2_h I__6194 (
            .O(N__30367),
            .I(N__30358));
    LocalMux I__6193 (
            .O(N__30364),
            .I(\b2v_inst11.N_369 ));
    LocalMux I__6192 (
            .O(N__30361),
            .I(\b2v_inst11.N_369 ));
    Odrv4 I__6191 (
            .O(N__30358),
            .I(\b2v_inst11.N_369 ));
    InMux I__6190 (
            .O(N__30351),
            .I(bfn_11_6_0_));
    InMux I__6189 (
            .O(N__30348),
            .I(N__30345));
    LocalMux I__6188 (
            .O(N__30345),
            .I(N__30342));
    Odrv4 I__6187 (
            .O(N__30342),
            .I(\b2v_inst11.un1_count_clk_2_axb_10 ));
    InMux I__6186 (
            .O(N__30339),
            .I(N__30330));
    InMux I__6185 (
            .O(N__30338),
            .I(N__30330));
    InMux I__6184 (
            .O(N__30337),
            .I(N__30330));
    LocalMux I__6183 (
            .O(N__30330),
            .I(N__30327));
    Odrv4 I__6182 (
            .O(N__30327),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ));
    InMux I__6181 (
            .O(N__30324),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__6180 (
            .O(N__30321),
            .I(N__30318));
    LocalMux I__6179 (
            .O(N__30318),
            .I(N__30315));
    Span4Mux_s3_h I__6178 (
            .O(N__30315),
            .I(N__30312));
    Odrv4 I__6177 (
            .O(N__30312),
            .I(\b2v_inst11.un1_count_clk_2_axb_11 ));
    InMux I__6176 (
            .O(N__30309),
            .I(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ));
    InMux I__6175 (
            .O(N__30306),
            .I(\b2v_inst11.un1_count_clk_2_cry_11 ));
    InMux I__6174 (
            .O(N__30303),
            .I(\b2v_inst11.un1_count_clk_2_cry_12 ));
    InMux I__6173 (
            .O(N__30300),
            .I(\b2v_inst11.un1_count_clk_2_cry_13 ));
    InMux I__6172 (
            .O(N__30297),
            .I(N__30291));
    InMux I__6171 (
            .O(N__30296),
            .I(N__30291));
    LocalMux I__6170 (
            .O(N__30291),
            .I(N__30276));
    InMux I__6169 (
            .O(N__30290),
            .I(N__30267));
    InMux I__6168 (
            .O(N__30289),
            .I(N__30267));
    InMux I__6167 (
            .O(N__30288),
            .I(N__30267));
    InMux I__6166 (
            .O(N__30287),
            .I(N__30267));
    InMux I__6165 (
            .O(N__30286),
            .I(N__30255));
    InMux I__6164 (
            .O(N__30285),
            .I(N__30255));
    InMux I__6163 (
            .O(N__30284),
            .I(N__30255));
    InMux I__6162 (
            .O(N__30283),
            .I(N__30255));
    InMux I__6161 (
            .O(N__30282),
            .I(N__30243));
    InMux I__6160 (
            .O(N__30281),
            .I(N__30243));
    InMux I__6159 (
            .O(N__30280),
            .I(N__30243));
    InMux I__6158 (
            .O(N__30279),
            .I(N__30243));
    Span4Mux_v I__6157 (
            .O(N__30276),
            .I(N__30240));
    LocalMux I__6156 (
            .O(N__30267),
            .I(N__30237));
    InMux I__6155 (
            .O(N__30266),
            .I(N__30230));
    InMux I__6154 (
            .O(N__30265),
            .I(N__30230));
    InMux I__6153 (
            .O(N__30264),
            .I(N__30230));
    LocalMux I__6152 (
            .O(N__30255),
            .I(N__30227));
    InMux I__6151 (
            .O(N__30254),
            .I(N__30220));
    InMux I__6150 (
            .O(N__30253),
            .I(N__30220));
    InMux I__6149 (
            .O(N__30252),
            .I(N__30220));
    LocalMux I__6148 (
            .O(N__30243),
            .I(N__30211));
    Span4Mux_s0_h I__6147 (
            .O(N__30240),
            .I(N__30211));
    Span4Mux_v I__6146 (
            .O(N__30237),
            .I(N__30211));
    LocalMux I__6145 (
            .O(N__30230),
            .I(N__30211));
    Odrv4 I__6144 (
            .O(N__30227),
            .I(\b2v_inst11.func_state_RNIIGCET1_0_1 ));
    LocalMux I__6143 (
            .O(N__30220),
            .I(\b2v_inst11.func_state_RNIIGCET1_0_1 ));
    Odrv4 I__6142 (
            .O(N__30211),
            .I(\b2v_inst11.func_state_RNIIGCET1_0_1 ));
    InMux I__6141 (
            .O(N__30204),
            .I(\b2v_inst11.un1_count_clk_2_cry_14 ));
    InMux I__6140 (
            .O(N__30201),
            .I(N__30196));
    InMux I__6139 (
            .O(N__30200),
            .I(N__30193));
    InMux I__6138 (
            .O(N__30199),
            .I(N__30190));
    LocalMux I__6137 (
            .O(N__30196),
            .I(N__30187));
    LocalMux I__6136 (
            .O(N__30193),
            .I(N__30184));
    LocalMux I__6135 (
            .O(N__30190),
            .I(N__30179));
    Span4Mux_v I__6134 (
            .O(N__30187),
            .I(N__30179));
    Odrv4 I__6133 (
            .O(N__30184),
            .I(\b2v_inst11.count_clk_1_11 ));
    Odrv4 I__6132 (
            .O(N__30179),
            .I(\b2v_inst11.count_clk_1_11 ));
    InMux I__6131 (
            .O(N__30174),
            .I(N__30170));
    InMux I__6130 (
            .O(N__30173),
            .I(N__30167));
    LocalMux I__6129 (
            .O(N__30170),
            .I(N__30164));
    LocalMux I__6128 (
            .O(N__30167),
            .I(N__30161));
    Span4Mux_h I__6127 (
            .O(N__30164),
            .I(N__30158));
    Odrv4 I__6126 (
            .O(N__30161),
            .I(\b2v_inst11.count_clk_0_11 ));
    Odrv4 I__6125 (
            .O(N__30158),
            .I(\b2v_inst11.count_clk_0_11 ));
    InMux I__6124 (
            .O(N__30153),
            .I(N__30143));
    InMux I__6123 (
            .O(N__30152),
            .I(N__30143));
    InMux I__6122 (
            .O(N__30151),
            .I(N__30143));
    InMux I__6121 (
            .O(N__30150),
            .I(N__30140));
    LocalMux I__6120 (
            .O(N__30143),
            .I(N__30137));
    LocalMux I__6119 (
            .O(N__30140),
            .I(N__30134));
    Span4Mux_h I__6118 (
            .O(N__30137),
            .I(N__30129));
    Span4Mux_h I__6117 (
            .O(N__30134),
            .I(N__30129));
    Odrv4 I__6116 (
            .O(N__30129),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    InMux I__6115 (
            .O(N__30126),
            .I(N__30120));
    InMux I__6114 (
            .O(N__30125),
            .I(N__30120));
    LocalMux I__6113 (
            .O(N__30120),
            .I(\b2v_inst11.count_clk_0_10 ));
    InMux I__6112 (
            .O(N__30117),
            .I(N__30114));
    LocalMux I__6111 (
            .O(N__30114),
            .I(N__30110));
    InMux I__6110 (
            .O(N__30113),
            .I(N__30107));
    Span4Mux_s2_h I__6109 (
            .O(N__30110),
            .I(N__30104));
    LocalMux I__6108 (
            .O(N__30107),
            .I(\b2v_inst11.un1_count_clk_2_axb_1 ));
    Odrv4 I__6107 (
            .O(N__30104),
            .I(\b2v_inst11.un1_count_clk_2_axb_1 ));
    CascadeMux I__6106 (
            .O(N__30099),
            .I(N__30096));
    InMux I__6105 (
            .O(N__30096),
            .I(N__30091));
    InMux I__6104 (
            .O(N__30095),
            .I(N__30088));
    CascadeMux I__6103 (
            .O(N__30094),
            .I(N__30085));
    LocalMux I__6102 (
            .O(N__30091),
            .I(N__30080));
    LocalMux I__6101 (
            .O(N__30088),
            .I(N__30077));
    InMux I__6100 (
            .O(N__30085),
            .I(N__30070));
    InMux I__6099 (
            .O(N__30084),
            .I(N__30070));
    InMux I__6098 (
            .O(N__30083),
            .I(N__30070));
    Span4Mux_s2_h I__6097 (
            .O(N__30080),
            .I(N__30067));
    Odrv12 I__6096 (
            .O(N__30077),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    LocalMux I__6095 (
            .O(N__30070),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    Odrv4 I__6094 (
            .O(N__30067),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    InMux I__6093 (
            .O(N__30060),
            .I(\b2v_inst11.un1_count_clk_2_cry_1 ));
    CascadeMux I__6092 (
            .O(N__30057),
            .I(N__30054));
    InMux I__6091 (
            .O(N__30054),
            .I(N__30051));
    LocalMux I__6090 (
            .O(N__30051),
            .I(N__30048));
    Odrv12 I__6089 (
            .O(N__30048),
            .I(\b2v_inst11.un1_count_clk_2_axb_3 ));
    InMux I__6088 (
            .O(N__30045),
            .I(N__30036));
    InMux I__6087 (
            .O(N__30044),
            .I(N__30036));
    InMux I__6086 (
            .O(N__30043),
            .I(N__30036));
    LocalMux I__6085 (
            .O(N__30036),
            .I(N__30033));
    Odrv4 I__6084 (
            .O(N__30033),
            .I(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ));
    InMux I__6083 (
            .O(N__30030),
            .I(\b2v_inst11.un1_count_clk_2_cry_2 ));
    InMux I__6082 (
            .O(N__30027),
            .I(\b2v_inst11.un1_count_clk_2_cry_3 ));
    InMux I__6081 (
            .O(N__30024),
            .I(\b2v_inst11.un1_count_clk_2_cry_4 ));
    InMux I__6080 (
            .O(N__30021),
            .I(\b2v_inst11.un1_count_clk_2_cry_5 ));
    InMux I__6079 (
            .O(N__30018),
            .I(\b2v_inst11.un1_count_clk_2_cry_6 ));
    InMux I__6078 (
            .O(N__30015),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__6077 (
            .O(N__30012),
            .I(\b2v_inst6.un2_count_1_cry_14 ));
    InMux I__6076 (
            .O(N__30009),
            .I(N__30006));
    LocalMux I__6075 (
            .O(N__30006),
            .I(\b2v_inst6.un2_count_1_axb_13 ));
    InMux I__6074 (
            .O(N__30003),
            .I(N__30000));
    LocalMux I__6073 (
            .O(N__30000),
            .I(\b2v_inst11.count_clkZ0Z_10 ));
    InMux I__6072 (
            .O(N__29997),
            .I(N__29994));
    LocalMux I__6071 (
            .O(N__29994),
            .I(\b2v_inst11.count_clkZ0Z_12 ));
    CascadeMux I__6070 (
            .O(N__29991),
            .I(\b2v_inst11.count_clkZ0Z_13_cascade_ ));
    InMux I__6069 (
            .O(N__29988),
            .I(N__29985));
    LocalMux I__6068 (
            .O(N__29985),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    CascadeMux I__6067 (
            .O(N__29982),
            .I(\b2v_inst11.un2_count_clk_17_0_o2_4_cascade_ ));
    InMux I__6066 (
            .O(N__29979),
            .I(N__29967));
    InMux I__6065 (
            .O(N__29978),
            .I(N__29967));
    InMux I__6064 (
            .O(N__29977),
            .I(N__29967));
    InMux I__6063 (
            .O(N__29976),
            .I(N__29967));
    LocalMux I__6062 (
            .O(N__29967),
            .I(N__29964));
    Span4Mux_v I__6061 (
            .O(N__29964),
            .I(N__29961));
    Odrv4 I__6060 (
            .O(N__29961),
            .I(\b2v_inst11.N_175 ));
    InMux I__6059 (
            .O(N__29958),
            .I(N__29954));
    InMux I__6058 (
            .O(N__29957),
            .I(N__29951));
    LocalMux I__6057 (
            .O(N__29954),
            .I(\b2v_inst6.un2_count_1_axb_7 ));
    LocalMux I__6056 (
            .O(N__29951),
            .I(\b2v_inst6.un2_count_1_axb_7 ));
    InMux I__6055 (
            .O(N__29946),
            .I(N__29940));
    InMux I__6054 (
            .O(N__29945),
            .I(N__29940));
    LocalMux I__6053 (
            .O(N__29940),
            .I(\b2v_inst6.un2_count_1_cry_6_THRU_CO ));
    InMux I__6052 (
            .O(N__29937),
            .I(\b2v_inst6.un2_count_1_cry_6 ));
    InMux I__6051 (
            .O(N__29934),
            .I(N__29931));
    LocalMux I__6050 (
            .O(N__29931),
            .I(N__29927));
    InMux I__6049 (
            .O(N__29930),
            .I(N__29924));
    Span4Mux_s2_h I__6048 (
            .O(N__29927),
            .I(N__29921));
    LocalMux I__6047 (
            .O(N__29924),
            .I(\b2v_inst6.un2_count_1_axb_8 ));
    Odrv4 I__6046 (
            .O(N__29921),
            .I(\b2v_inst6.un2_count_1_axb_8 ));
    CascadeMux I__6045 (
            .O(N__29916),
            .I(N__29913));
    InMux I__6044 (
            .O(N__29913),
            .I(N__29907));
    InMux I__6043 (
            .O(N__29912),
            .I(N__29907));
    LocalMux I__6042 (
            .O(N__29907),
            .I(N__29904));
    Span4Mux_s1_v I__6041 (
            .O(N__29904),
            .I(N__29901));
    Odrv4 I__6040 (
            .O(N__29901),
            .I(\b2v_inst6.un2_count_1_cry_7_THRU_CO ));
    InMux I__6039 (
            .O(N__29898),
            .I(\b2v_inst6.un2_count_1_cry_7 ));
    InMux I__6038 (
            .O(N__29895),
            .I(N__29891));
    InMux I__6037 (
            .O(N__29894),
            .I(N__29888));
    LocalMux I__6036 (
            .O(N__29891),
            .I(N__29885));
    LocalMux I__6035 (
            .O(N__29888),
            .I(N__29880));
    Span4Mux_v I__6034 (
            .O(N__29885),
            .I(N__29880));
    Odrv4 I__6033 (
            .O(N__29880),
            .I(\b2v_inst6.un2_count_1_axb_9 ));
    InMux I__6032 (
            .O(N__29877),
            .I(N__29871));
    InMux I__6031 (
            .O(N__29876),
            .I(N__29871));
    LocalMux I__6030 (
            .O(N__29871),
            .I(N__29868));
    Span4Mux_s2_v I__6029 (
            .O(N__29868),
            .I(N__29865));
    Odrv4 I__6028 (
            .O(N__29865),
            .I(\b2v_inst6.un2_count_1_cry_8_THRU_CO ));
    InMux I__6027 (
            .O(N__29862),
            .I(bfn_11_3_0_));
    InMux I__6026 (
            .O(N__29859),
            .I(\b2v_inst6.un2_count_1_cry_9 ));
    InMux I__6025 (
            .O(N__29856),
            .I(N__29850));
    InMux I__6024 (
            .O(N__29855),
            .I(N__29850));
    LocalMux I__6023 (
            .O(N__29850),
            .I(N__29847));
    Odrv4 I__6022 (
            .O(N__29847),
            .I(\b2v_inst6.un2_count_1_cry_10_THRU_CO ));
    InMux I__6021 (
            .O(N__29844),
            .I(\b2v_inst6.un2_count_1_cry_10 ));
    InMux I__6020 (
            .O(N__29841),
            .I(\b2v_inst6.un2_count_1_cry_11 ));
    InMux I__6019 (
            .O(N__29838),
            .I(\b2v_inst6.un2_count_1_cry_12 ));
    InMux I__6018 (
            .O(N__29835),
            .I(\b2v_inst6.un2_count_1_cry_13 ));
    CascadeMux I__6017 (
            .O(N__29832),
            .I(\b2v_inst6.count_rst_3_cascade_ ));
    CascadeMux I__6016 (
            .O(N__29829),
            .I(\b2v_inst6.countZ0Z_11_cascade_ ));
    InMux I__6015 (
            .O(N__29826),
            .I(N__29823));
    LocalMux I__6014 (
            .O(N__29823),
            .I(\b2v_inst6.count_0_11 ));
    InMux I__6013 (
            .O(N__29820),
            .I(N__29810));
    InMux I__6012 (
            .O(N__29819),
            .I(N__29797));
    InMux I__6011 (
            .O(N__29818),
            .I(N__29797));
    InMux I__6010 (
            .O(N__29817),
            .I(N__29797));
    InMux I__6009 (
            .O(N__29816),
            .I(N__29797));
    InMux I__6008 (
            .O(N__29815),
            .I(N__29797));
    InMux I__6007 (
            .O(N__29814),
            .I(N__29797));
    InMux I__6006 (
            .O(N__29813),
            .I(N__29790));
    LocalMux I__6005 (
            .O(N__29810),
            .I(N__29787));
    LocalMux I__6004 (
            .O(N__29797),
            .I(N__29784));
    InMux I__6003 (
            .O(N__29796),
            .I(N__29770));
    InMux I__6002 (
            .O(N__29795),
            .I(N__29770));
    InMux I__6001 (
            .O(N__29794),
            .I(N__29770));
    InMux I__6000 (
            .O(N__29793),
            .I(N__29770));
    LocalMux I__5999 (
            .O(N__29790),
            .I(N__29763));
    Span4Mux_v I__5998 (
            .O(N__29787),
            .I(N__29763));
    Span4Mux_s1_v I__5997 (
            .O(N__29784),
            .I(N__29763));
    InMux I__5996 (
            .O(N__29783),
            .I(N__29754));
    InMux I__5995 (
            .O(N__29782),
            .I(N__29754));
    InMux I__5994 (
            .O(N__29781),
            .I(N__29754));
    InMux I__5993 (
            .O(N__29780),
            .I(N__29754));
    InMux I__5992 (
            .O(N__29779),
            .I(N__29751));
    LocalMux I__5991 (
            .O(N__29770),
            .I(\b2v_inst6.N_394 ));
    Odrv4 I__5990 (
            .O(N__29763),
            .I(\b2v_inst6.N_394 ));
    LocalMux I__5989 (
            .O(N__29754),
            .I(\b2v_inst6.N_394 ));
    LocalMux I__5988 (
            .O(N__29751),
            .I(\b2v_inst6.N_394 ));
    InMux I__5987 (
            .O(N__29742),
            .I(\b2v_inst6.un2_count_1_cry_1 ));
    InMux I__5986 (
            .O(N__29739),
            .I(N__29735));
    CascadeMux I__5985 (
            .O(N__29738),
            .I(N__29732));
    LocalMux I__5984 (
            .O(N__29735),
            .I(N__29729));
    InMux I__5983 (
            .O(N__29732),
            .I(N__29726));
    Span4Mux_s3_h I__5982 (
            .O(N__29729),
            .I(N__29723));
    LocalMux I__5981 (
            .O(N__29726),
            .I(\b2v_inst6.un2_count_1_axb_3 ));
    Odrv4 I__5980 (
            .O(N__29723),
            .I(\b2v_inst6.un2_count_1_axb_3 ));
    InMux I__5979 (
            .O(N__29718),
            .I(N__29712));
    InMux I__5978 (
            .O(N__29717),
            .I(N__29712));
    LocalMux I__5977 (
            .O(N__29712),
            .I(N__29709));
    Span4Mux_s1_v I__5976 (
            .O(N__29709),
            .I(N__29706));
    Odrv4 I__5975 (
            .O(N__29706),
            .I(\b2v_inst6.un2_count_1_cry_2_THRU_CO ));
    InMux I__5974 (
            .O(N__29703),
            .I(\b2v_inst6.un2_count_1_cry_2 ));
    InMux I__5973 (
            .O(N__29700),
            .I(N__29695));
    CascadeMux I__5972 (
            .O(N__29699),
            .I(N__29692));
    CascadeMux I__5971 (
            .O(N__29698),
            .I(N__29689));
    LocalMux I__5970 (
            .O(N__29695),
            .I(N__29686));
    InMux I__5969 (
            .O(N__29692),
            .I(N__29681));
    InMux I__5968 (
            .O(N__29689),
            .I(N__29681));
    Span4Mux_v I__5967 (
            .O(N__29686),
            .I(N__29678));
    LocalMux I__5966 (
            .O(N__29681),
            .I(\b2v_inst6.un2_count_1_axb_4 ));
    Odrv4 I__5965 (
            .O(N__29678),
            .I(\b2v_inst6.un2_count_1_axb_4 ));
    InMux I__5964 (
            .O(N__29673),
            .I(N__29667));
    InMux I__5963 (
            .O(N__29672),
            .I(N__29667));
    LocalMux I__5962 (
            .O(N__29667),
            .I(N__29664));
    Span4Mux_h I__5961 (
            .O(N__29664),
            .I(N__29661));
    Odrv4 I__5960 (
            .O(N__29661),
            .I(\b2v_inst6.un2_count_1_cry_3_THRU_CO ));
    InMux I__5959 (
            .O(N__29658),
            .I(\b2v_inst6.un2_count_1_cry_3 ));
    InMux I__5958 (
            .O(N__29655),
            .I(N__29649));
    InMux I__5957 (
            .O(N__29654),
            .I(N__29649));
    LocalMux I__5956 (
            .O(N__29649),
            .I(\b2v_inst6.un2_count_1_cry_4_THRU_CO ));
    InMux I__5955 (
            .O(N__29646),
            .I(\b2v_inst6.un2_count_1_cry_4 ));
    InMux I__5954 (
            .O(N__29643),
            .I(\b2v_inst6.un2_count_1_cry_5 ));
    CascadeMux I__5953 (
            .O(N__29640),
            .I(\b2v_inst11.N_11_cascade_ ));
    InMux I__5952 (
            .O(N__29637),
            .I(N__29634));
    LocalMux I__5951 (
            .O(N__29634),
            .I(\b2v_inst11.N_35_0 ));
    CascadeMux I__5950 (
            .O(N__29631),
            .I(\b2v_inst11.N_13_cascade_ ));
    CascadeMux I__5949 (
            .O(N__29628),
            .I(N__29624));
    InMux I__5948 (
            .O(N__29627),
            .I(N__29619));
    InMux I__5947 (
            .O(N__29624),
            .I(N__29619));
    LocalMux I__5946 (
            .O(N__29619),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_11 ));
    CascadeMux I__5945 (
            .O(N__29616),
            .I(N__29613));
    InMux I__5944 (
            .O(N__29613),
            .I(N__29610));
    LocalMux I__5943 (
            .O(N__29610),
            .I(\b2v_inst11.g0_6_a5_1_0 ));
    CascadeMux I__5942 (
            .O(N__29607),
            .I(\b2v_inst6.count_rst_7_cascade_ ));
    CascadeMux I__5941 (
            .O(N__29604),
            .I(\b2v_inst6.un2_count_1_axb_7_cascade_ ));
    InMux I__5940 (
            .O(N__29601),
            .I(N__29598));
    LocalMux I__5939 (
            .O(N__29598),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_6 ));
    CascadeMux I__5938 (
            .O(N__29595),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_6_cascade_ ));
    InMux I__5937 (
            .O(N__29592),
            .I(N__29589));
    LocalMux I__5936 (
            .O(N__29589),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ));
    CascadeMux I__5935 (
            .O(N__29586),
            .I(N__29583));
    InMux I__5934 (
            .O(N__29583),
            .I(N__29580));
    LocalMux I__5933 (
            .O(N__29580),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_15 ));
    CascadeMux I__5932 (
            .O(N__29577),
            .I(N__29574));
    InMux I__5931 (
            .O(N__29574),
            .I(N__29571));
    LocalMux I__5930 (
            .O(N__29571),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_14 ));
    InMux I__5929 (
            .O(N__29568),
            .I(N__29562));
    InMux I__5928 (
            .O(N__29567),
            .I(N__29562));
    LocalMux I__5927 (
            .O(N__29562),
            .I(\b2v_inst11.un1_dutycycle_53_44_0_0 ));
    InMux I__5926 (
            .O(N__29559),
            .I(N__29556));
    LocalMux I__5925 (
            .O(N__29556),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_8 ));
    CascadeMux I__5924 (
            .O(N__29553),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_ ));
    InMux I__5923 (
            .O(N__29550),
            .I(N__29547));
    LocalMux I__5922 (
            .O(N__29547),
            .I(N__29544));
    Span4Mux_s1_v I__5921 (
            .O(N__29544),
            .I(N__29541));
    Odrv4 I__5920 (
            .O(N__29541),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_7 ));
    CascadeMux I__5919 (
            .O(N__29538),
            .I(N__29535));
    InMux I__5918 (
            .O(N__29535),
            .I(N__29532));
    LocalMux I__5917 (
            .O(N__29532),
            .I(\b2v_inst11.un1_dutycycle_53_axb_10 ));
    InMux I__5916 (
            .O(N__29529),
            .I(N__29526));
    LocalMux I__5915 (
            .O(N__29526),
            .I(N__29522));
    InMux I__5914 (
            .O(N__29525),
            .I(N__29519));
    Odrv4 I__5913 (
            .O(N__29522),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_7 ));
    LocalMux I__5912 (
            .O(N__29519),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_7 ));
    InMux I__5911 (
            .O(N__29514),
            .I(N__29511));
    LocalMux I__5910 (
            .O(N__29511),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_7 ));
    InMux I__5909 (
            .O(N__29508),
            .I(N__29504));
    InMux I__5908 (
            .O(N__29507),
            .I(N__29501));
    LocalMux I__5907 (
            .O(N__29504),
            .I(N__29498));
    LocalMux I__5906 (
            .O(N__29501),
            .I(\b2v_inst11.CO2_THRU_CO ));
    Odrv4 I__5905 (
            .O(N__29498),
            .I(\b2v_inst11.CO2_THRU_CO ));
    CascadeMux I__5904 (
            .O(N__29493),
            .I(N__29490));
    InMux I__5903 (
            .O(N__29490),
            .I(N__29487));
    LocalMux I__5902 (
            .O(N__29487),
            .I(N__29484));
    Odrv4 I__5901 (
            .O(N__29484),
            .I(\b2v_inst11.mult1_un54_sum_axb_6_i_l_fx ));
    CascadeMux I__5900 (
            .O(N__29481),
            .I(N__29478));
    InMux I__5899 (
            .O(N__29478),
            .I(N__29471));
    InMux I__5898 (
            .O(N__29477),
            .I(N__29471));
    InMux I__5897 (
            .O(N__29476),
            .I(N__29468));
    LocalMux I__5896 (
            .O(N__29471),
            .I(N__29465));
    LocalMux I__5895 (
            .O(N__29468),
            .I(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ));
    Odrv4 I__5894 (
            .O(N__29465),
            .I(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ));
    CascadeMux I__5893 (
            .O(N__29460),
            .I(N__29457));
    InMux I__5892 (
            .O(N__29457),
            .I(N__29454));
    LocalMux I__5891 (
            .O(N__29454),
            .I(N__29451));
    Odrv4 I__5890 (
            .O(N__29451),
            .I(\b2v_inst11.mult1_un54_sum_axb_5_i_l_ofx ));
    CascadeMux I__5889 (
            .O(N__29448),
            .I(N__29443));
    CascadeMux I__5888 (
            .O(N__29447),
            .I(N__29438));
    InMux I__5887 (
            .O(N__29446),
            .I(N__29435));
    InMux I__5886 (
            .O(N__29443),
            .I(N__29432));
    InMux I__5885 (
            .O(N__29442),
            .I(N__29425));
    InMux I__5884 (
            .O(N__29441),
            .I(N__29425));
    InMux I__5883 (
            .O(N__29438),
            .I(N__29425));
    LocalMux I__5882 (
            .O(N__29435),
            .I(N__29422));
    LocalMux I__5881 (
            .O(N__29432),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0 ));
    LocalMux I__5880 (
            .O(N__29425),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0 ));
    Odrv4 I__5879 (
            .O(N__29422),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0 ));
    CascadeMux I__5878 (
            .O(N__29415),
            .I(N__29410));
    InMux I__5877 (
            .O(N__29414),
            .I(N__29406));
    InMux I__5876 (
            .O(N__29413),
            .I(N__29399));
    InMux I__5875 (
            .O(N__29410),
            .I(N__29399));
    InMux I__5874 (
            .O(N__29409),
            .I(N__29399));
    LocalMux I__5873 (
            .O(N__29406),
            .I(\b2v_inst11.mult1_un40_sum_i_2 ));
    LocalMux I__5872 (
            .O(N__29399),
            .I(\b2v_inst11.mult1_un40_sum_i_2 ));
    CascadeMux I__5871 (
            .O(N__29394),
            .I(N__29391));
    InMux I__5870 (
            .O(N__29391),
            .I(N__29388));
    LocalMux I__5869 (
            .O(N__29388),
            .I(N__29385));
    Odrv4 I__5868 (
            .O(N__29385),
            .I(\b2v_inst11.mult1_un47_sum1_3 ));
    CascadeMux I__5867 (
            .O(N__29382),
            .I(\b2v_inst11.un1_dutycycle_53_axb_12_cascade_ ));
    InMux I__5866 (
            .O(N__29379),
            .I(N__29376));
    LocalMux I__5865 (
            .O(N__29376),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_15 ));
    CascadeMux I__5864 (
            .O(N__29373),
            .I(N__29370));
    InMux I__5863 (
            .O(N__29370),
            .I(N__29367));
    LocalMux I__5862 (
            .O(N__29367),
            .I(\b2v_inst11.dutycycle_eena_9 ));
    InMux I__5861 (
            .O(N__29364),
            .I(N__29358));
    InMux I__5860 (
            .O(N__29363),
            .I(N__29358));
    LocalMux I__5859 (
            .O(N__29358),
            .I(\b2v_inst11.dutycycleZ1Z_12 ));
    InMux I__5858 (
            .O(N__29355),
            .I(N__29349));
    InMux I__5857 (
            .O(N__29354),
            .I(N__29349));
    LocalMux I__5856 (
            .O(N__29349),
            .I(\b2v_inst11.dutycycleZ1Z_11 ));
    InMux I__5855 (
            .O(N__29346),
            .I(N__29343));
    LocalMux I__5854 (
            .O(N__29343),
            .I(\b2v_inst11.dutycycle_eena_7 ));
    InMux I__5853 (
            .O(N__29340),
            .I(N__29337));
    LocalMux I__5852 (
            .O(N__29337),
            .I(\b2v_inst11.N_6_0 ));
    CascadeMux I__5851 (
            .O(N__29334),
            .I(\b2v_inst11.N_8_cascade_ ));
    InMux I__5850 (
            .O(N__29331),
            .I(N__29328));
    LocalMux I__5849 (
            .O(N__29328),
            .I(N__29324));
    InMux I__5848 (
            .O(N__29327),
            .I(N__29321));
    Span4Mux_h I__5847 (
            .O(N__29324),
            .I(N__29318));
    LocalMux I__5846 (
            .O(N__29321),
            .I(\b2v_inst11.N_355 ));
    Odrv4 I__5845 (
            .O(N__29318),
            .I(\b2v_inst11.N_355 ));
    CascadeMux I__5844 (
            .O(N__29313),
            .I(\b2v_inst11.g0_6_a5_0_0_cascade_ ));
    InMux I__5843 (
            .O(N__29310),
            .I(N__29307));
    LocalMux I__5842 (
            .O(N__29307),
            .I(\b2v_inst11.g0_6_a5_2_1 ));
    InMux I__5841 (
            .O(N__29304),
            .I(N__29301));
    LocalMux I__5840 (
            .O(N__29301),
            .I(N__29298));
    Span4Mux_v I__5839 (
            .O(N__29298),
            .I(N__29294));
    InMux I__5838 (
            .O(N__29297),
            .I(N__29291));
    Odrv4 I__5837 (
            .O(N__29294),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    LocalMux I__5836 (
            .O(N__29291),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    CascadeMux I__5835 (
            .O(N__29286),
            .I(\b2v_inst11.dutycycle_eena_9_cascade_ ));
    CascadeMux I__5834 (
            .O(N__29283),
            .I(\b2v_inst11.dutycycle_eena_7_cascade_ ));
    CascadeMux I__5833 (
            .O(N__29280),
            .I(N__29272));
    InMux I__5832 (
            .O(N__29279),
            .I(N__29263));
    InMux I__5831 (
            .O(N__29278),
            .I(N__29263));
    InMux I__5830 (
            .O(N__29277),
            .I(N__29263));
    InMux I__5829 (
            .O(N__29276),
            .I(N__29263));
    InMux I__5828 (
            .O(N__29275),
            .I(N__29258));
    InMux I__5827 (
            .O(N__29272),
            .I(N__29258));
    LocalMux I__5826 (
            .O(N__29263),
            .I(N__29253));
    LocalMux I__5825 (
            .O(N__29258),
            .I(N__29253));
    Span4Mux_h I__5824 (
            .O(N__29253),
            .I(N__29250));
    Odrv4 I__5823 (
            .O(N__29250),
            .I(\b2v_inst11.N_2943_i ));
    CascadeMux I__5822 (
            .O(N__29247),
            .I(N__29244));
    InMux I__5821 (
            .O(N__29244),
            .I(N__29236));
    InMux I__5820 (
            .O(N__29243),
            .I(N__29236));
    InMux I__5819 (
            .O(N__29242),
            .I(N__29233));
    InMux I__5818 (
            .O(N__29241),
            .I(N__29230));
    LocalMux I__5817 (
            .O(N__29236),
            .I(N__29225));
    LocalMux I__5816 (
            .O(N__29233),
            .I(N__29225));
    LocalMux I__5815 (
            .O(N__29230),
            .I(N__29221));
    Span4Mux_h I__5814 (
            .O(N__29225),
            .I(N__29218));
    InMux I__5813 (
            .O(N__29224),
            .I(N__29215));
    Odrv4 I__5812 (
            .O(N__29221),
            .I(\b2v_inst11.func_state_RNIDQ4A1Z0Z_1 ));
    Odrv4 I__5811 (
            .O(N__29218),
            .I(\b2v_inst11.func_state_RNIDQ4A1Z0Z_1 ));
    LocalMux I__5810 (
            .O(N__29215),
            .I(\b2v_inst11.func_state_RNIDQ4A1Z0Z_1 ));
    CascadeMux I__5809 (
            .O(N__29208),
            .I(\b2v_inst11.N_360_cascade_ ));
    InMux I__5808 (
            .O(N__29205),
            .I(N__29202));
    LocalMux I__5807 (
            .O(N__29202),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ));
    InMux I__5806 (
            .O(N__29199),
            .I(N__29193));
    InMux I__5805 (
            .O(N__29198),
            .I(N__29193));
    LocalMux I__5804 (
            .O(N__29193),
            .I(\b2v_inst11.N_234_N ));
    InMux I__5803 (
            .O(N__29190),
            .I(N__29187));
    LocalMux I__5802 (
            .O(N__29187),
            .I(N__29184));
    Span4Mux_h I__5801 (
            .O(N__29184),
            .I(N__29181));
    Odrv4 I__5800 (
            .O(N__29181),
            .I(\b2v_inst11.N_309 ));
    InMux I__5799 (
            .O(N__29178),
            .I(N__29175));
    LocalMux I__5798 (
            .O(N__29175),
            .I(N__29172));
    Odrv4 I__5797 (
            .O(N__29172),
            .I(\b2v_inst11.un1_dutycycle_96_0_a3_1 ));
    CascadeMux I__5796 (
            .O(N__29169),
            .I(N__29166));
    InMux I__5795 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__5794 (
            .O(N__29163),
            .I(N__29159));
    InMux I__5793 (
            .O(N__29162),
            .I(N__29156));
    Odrv4 I__5792 (
            .O(N__29159),
            .I(\b2v_inst11.dutycycle_eena_0 ));
    LocalMux I__5791 (
            .O(N__29156),
            .I(\b2v_inst11.dutycycle_eena_0 ));
    InMux I__5790 (
            .O(N__29151),
            .I(N__29146));
    InMux I__5789 (
            .O(N__29150),
            .I(N__29141));
    InMux I__5788 (
            .O(N__29149),
            .I(N__29141));
    LocalMux I__5787 (
            .O(N__29146),
            .I(N__29138));
    LocalMux I__5786 (
            .O(N__29141),
            .I(N__29135));
    Odrv4 I__5785 (
            .O(N__29138),
            .I(\b2v_inst11.un1_clk_100khz_25_and_i_0_1_0 ));
    Odrv4 I__5784 (
            .O(N__29135),
            .I(\b2v_inst11.un1_clk_100khz_25_and_i_0_1_0 ));
    InMux I__5783 (
            .O(N__29130),
            .I(N__29127));
    LocalMux I__5782 (
            .O(N__29127),
            .I(\b2v_inst11.N_186_i ));
    InMux I__5781 (
            .O(N__29124),
            .I(N__29121));
    LocalMux I__5780 (
            .O(N__29121),
            .I(\b2v_inst11.N_117_f0_1 ));
    CascadeMux I__5779 (
            .O(N__29118),
            .I(N__29113));
    IoInMux I__5778 (
            .O(N__29117),
            .I(N__29109));
    IoInMux I__5777 (
            .O(N__29116),
            .I(N__29104));
    InMux I__5776 (
            .O(N__29113),
            .I(N__29099));
    InMux I__5775 (
            .O(N__29112),
            .I(N__29099));
    LocalMux I__5774 (
            .O(N__29109),
            .I(N__29096));
    CascadeMux I__5773 (
            .O(N__29108),
            .I(N__29093));
    CascadeMux I__5772 (
            .O(N__29107),
            .I(N__29090));
    LocalMux I__5771 (
            .O(N__29104),
            .I(N__29084));
    LocalMux I__5770 (
            .O(N__29099),
            .I(N__29081));
    IoSpan4Mux I__5769 (
            .O(N__29096),
            .I(N__29078));
    InMux I__5768 (
            .O(N__29093),
            .I(N__29075));
    InMux I__5767 (
            .O(N__29090),
            .I(N__29068));
    InMux I__5766 (
            .O(N__29089),
            .I(N__29068));
    InMux I__5765 (
            .O(N__29088),
            .I(N__29068));
    CascadeMux I__5764 (
            .O(N__29087),
            .I(N__29065));
    Span4Mux_s2_h I__5763 (
            .O(N__29084),
            .I(N__29062));
    Span4Mux_h I__5762 (
            .O(N__29081),
            .I(N__29059));
    Span4Mux_s2_h I__5761 (
            .O(N__29078),
            .I(N__29056));
    LocalMux I__5760 (
            .O(N__29075),
            .I(N__29051));
    LocalMux I__5759 (
            .O(N__29068),
            .I(N__29051));
    InMux I__5758 (
            .O(N__29065),
            .I(N__29048));
    Span4Mux_h I__5757 (
            .O(N__29062),
            .I(N__29043));
    Span4Mux_v I__5756 (
            .O(N__29059),
            .I(N__29043));
    Span4Mux_h I__5755 (
            .O(N__29056),
            .I(N__29038));
    Span4Mux_h I__5754 (
            .O(N__29051),
            .I(N__29038));
    LocalMux I__5753 (
            .O(N__29048),
            .I(v5s_enn));
    Odrv4 I__5752 (
            .O(N__29043),
            .I(v5s_enn));
    Odrv4 I__5751 (
            .O(N__29038),
            .I(v5s_enn));
    CascadeMux I__5750 (
            .O(N__29031),
            .I(\b2v_inst11.N_117_f0_1_cascade_ ));
    InMux I__5749 (
            .O(N__29028),
            .I(N__29022));
    InMux I__5748 (
            .O(N__29027),
            .I(N__29022));
    LocalMux I__5747 (
            .O(N__29022),
            .I(\b2v_inst11.dutycycle_eena ));
    InMux I__5746 (
            .O(N__29019),
            .I(N__29013));
    InMux I__5745 (
            .O(N__29018),
            .I(N__29013));
    LocalMux I__5744 (
            .O(N__29013),
            .I(\b2v_inst11.dutycycleZ1Z_2 ));
    CascadeMux I__5743 (
            .O(N__29010),
            .I(N__29006));
    InMux I__5742 (
            .O(N__29009),
            .I(N__29003));
    InMux I__5741 (
            .O(N__29006),
            .I(N__29000));
    LocalMux I__5740 (
            .O(N__29003),
            .I(N__28995));
    LocalMux I__5739 (
            .O(N__29000),
            .I(N__28995));
    Span4Mux_v I__5738 (
            .O(N__28995),
            .I(N__28992));
    Odrv4 I__5737 (
            .O(N__28992),
            .I(\b2v_inst11.N_73 ));
    InMux I__5736 (
            .O(N__28989),
            .I(N__28983));
    InMux I__5735 (
            .O(N__28988),
            .I(N__28983));
    LocalMux I__5734 (
            .O(N__28983),
            .I(\b2v_inst11.dutycycle_eena_1 ));
    InMux I__5733 (
            .O(N__28980),
            .I(N__28977));
    LocalMux I__5732 (
            .O(N__28977),
            .I(N__28974));
    Span4Mux_h I__5731 (
            .O(N__28974),
            .I(N__28971));
    Odrv4 I__5730 (
            .O(N__28971),
            .I(\b2v_inst11.N_159 ));
    CascadeMux I__5729 (
            .O(N__28968),
            .I(\b2v_inst11.dutycycleZ0Z_1_cascade_ ));
    InMux I__5728 (
            .O(N__28965),
            .I(N__28961));
    CascadeMux I__5727 (
            .O(N__28964),
            .I(N__28957));
    LocalMux I__5726 (
            .O(N__28961),
            .I(N__28953));
    InMux I__5725 (
            .O(N__28960),
            .I(N__28946));
    InMux I__5724 (
            .O(N__28957),
            .I(N__28946));
    InMux I__5723 (
            .O(N__28956),
            .I(N__28946));
    Span4Mux_h I__5722 (
            .O(N__28953),
            .I(N__28943));
    LocalMux I__5721 (
            .O(N__28946),
            .I(\b2v_inst11.N_363 ));
    Odrv4 I__5720 (
            .O(N__28943),
            .I(\b2v_inst11.N_363 ));
    CascadeMux I__5719 (
            .O(N__28938),
            .I(\b2v_inst11.dutycycle_1_0_1_cascade_ ));
    InMux I__5718 (
            .O(N__28935),
            .I(N__28929));
    InMux I__5717 (
            .O(N__28934),
            .I(N__28929));
    LocalMux I__5716 (
            .O(N__28929),
            .I(N__28926));
    Odrv4 I__5715 (
            .O(N__28926),
            .I(\b2v_inst11.dutycycleZ1Z_1 ));
    InMux I__5714 (
            .O(N__28923),
            .I(N__28920));
    LocalMux I__5713 (
            .O(N__28920),
            .I(\b2v_inst11.dutycycle_1_0_0 ));
    CascadeMux I__5712 (
            .O(N__28917),
            .I(N__28914));
    InMux I__5711 (
            .O(N__28914),
            .I(N__28908));
    InMux I__5710 (
            .O(N__28913),
            .I(N__28908));
    LocalMux I__5709 (
            .O(N__28908),
            .I(\b2v_inst11.dutycycleZ1Z_0 ));
    CascadeMux I__5708 (
            .O(N__28905),
            .I(\b2v_inst11.dutycycle_1_0_0_cascade_ ));
    InMux I__5707 (
            .O(N__28902),
            .I(N__28896));
    InMux I__5706 (
            .O(N__28901),
            .I(N__28896));
    LocalMux I__5705 (
            .O(N__28896),
            .I(\b2v_inst11.dutycycle_RNI_8Z0Z_0 ));
    InMux I__5704 (
            .O(N__28893),
            .I(N__28889));
    InMux I__5703 (
            .O(N__28892),
            .I(N__28886));
    LocalMux I__5702 (
            .O(N__28889),
            .I(N__28880));
    LocalMux I__5701 (
            .O(N__28886),
            .I(N__28880));
    InMux I__5700 (
            .O(N__28885),
            .I(N__28877));
    Odrv4 I__5699 (
            .O(N__28880),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_2 ));
    LocalMux I__5698 (
            .O(N__28877),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_2 ));
    CascadeMux I__5697 (
            .O(N__28872),
            .I(N__28868));
    InMux I__5696 (
            .O(N__28871),
            .I(N__28863));
    InMux I__5695 (
            .O(N__28868),
            .I(N__28863));
    LocalMux I__5694 (
            .O(N__28863),
            .I(N__28855));
    InMux I__5693 (
            .O(N__28862),
            .I(N__28852));
    InMux I__5692 (
            .O(N__28861),
            .I(N__28849));
    InMux I__5691 (
            .O(N__28860),
            .I(N__28842));
    InMux I__5690 (
            .O(N__28859),
            .I(N__28842));
    InMux I__5689 (
            .O(N__28858),
            .I(N__28842));
    Span4Mux_h I__5688 (
            .O(N__28855),
            .I(N__28839));
    LocalMux I__5687 (
            .O(N__28852),
            .I(\b2v_inst11.N_19_i ));
    LocalMux I__5686 (
            .O(N__28849),
            .I(\b2v_inst11.N_19_i ));
    LocalMux I__5685 (
            .O(N__28842),
            .I(\b2v_inst11.N_19_i ));
    Odrv4 I__5684 (
            .O(N__28839),
            .I(\b2v_inst11.N_19_i ));
    CascadeMux I__5683 (
            .O(N__28830),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_0_cascade_ ));
    InMux I__5682 (
            .O(N__28827),
            .I(N__28824));
    LocalMux I__5681 (
            .O(N__28824),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1 ));
    CascadeMux I__5680 (
            .O(N__28821),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    CascadeMux I__5679 (
            .O(N__28818),
            .I(\b2v_inst11.N_186_i_cascade_ ));
    CascadeMux I__5678 (
            .O(N__28815),
            .I(N__28811));
    InMux I__5677 (
            .O(N__28814),
            .I(N__28801));
    InMux I__5676 (
            .O(N__28811),
            .I(N__28801));
    InMux I__5675 (
            .O(N__28810),
            .I(N__28801));
    InMux I__5674 (
            .O(N__28809),
            .I(N__28797));
    InMux I__5673 (
            .O(N__28808),
            .I(N__28791));
    LocalMux I__5672 (
            .O(N__28801),
            .I(N__28787));
    InMux I__5671 (
            .O(N__28800),
            .I(N__28784));
    LocalMux I__5670 (
            .O(N__28797),
            .I(N__28781));
    InMux I__5669 (
            .O(N__28796),
            .I(N__28774));
    InMux I__5668 (
            .O(N__28795),
            .I(N__28774));
    InMux I__5667 (
            .O(N__28794),
            .I(N__28774));
    LocalMux I__5666 (
            .O(N__28791),
            .I(N__28771));
    InMux I__5665 (
            .O(N__28790),
            .I(N__28766));
    Span4Mux_h I__5664 (
            .O(N__28787),
            .I(N__28763));
    LocalMux I__5663 (
            .O(N__28784),
            .I(N__28754));
    Span4Mux_v I__5662 (
            .O(N__28781),
            .I(N__28754));
    LocalMux I__5661 (
            .O(N__28774),
            .I(N__28754));
    Span4Mux_h I__5660 (
            .O(N__28771),
            .I(N__28754));
    InMux I__5659 (
            .O(N__28770),
            .I(N__28749));
    InMux I__5658 (
            .O(N__28769),
            .I(N__28749));
    LocalMux I__5657 (
            .O(N__28766),
            .I(curr_state_RNID8DP1_0_0));
    Odrv4 I__5656 (
            .O(N__28763),
            .I(curr_state_RNID8DP1_0_0));
    Odrv4 I__5655 (
            .O(N__28754),
            .I(curr_state_RNID8DP1_0_0));
    LocalMux I__5654 (
            .O(N__28749),
            .I(curr_state_RNID8DP1_0_0));
    InMux I__5653 (
            .O(N__28740),
            .I(N__28737));
    LocalMux I__5652 (
            .O(N__28737),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0_0 ));
    CascadeMux I__5651 (
            .O(N__28734),
            .I(N__28730));
    InMux I__5650 (
            .O(N__28733),
            .I(N__28725));
    InMux I__5649 (
            .O(N__28730),
            .I(N__28725));
    LocalMux I__5648 (
            .O(N__28725),
            .I(\b2v_inst11.N_160_i ));
    CascadeMux I__5647 (
            .O(N__28722),
            .I(\b2v_inst11.N_160_i_cascade_ ));
    CascadeMux I__5646 (
            .O(N__28719),
            .I(N__28715));
    InMux I__5645 (
            .O(N__28718),
            .I(N__28711));
    InMux I__5644 (
            .O(N__28715),
            .I(N__28706));
    InMux I__5643 (
            .O(N__28714),
            .I(N__28706));
    LocalMux I__5642 (
            .O(N__28711),
            .I(N__28702));
    LocalMux I__5641 (
            .O(N__28706),
            .I(N__28699));
    InMux I__5640 (
            .O(N__28705),
            .I(N__28696));
    Span4Mux_v I__5639 (
            .O(N__28702),
            .I(N__28693));
    Span4Mux_h I__5638 (
            .O(N__28699),
            .I(N__28690));
    LocalMux I__5637 (
            .O(N__28696),
            .I(N__28687));
    Odrv4 I__5636 (
            .O(N__28693),
            .I(\b2v_inst11.func_state_RNI5DLRZ0Z_0 ));
    Odrv4 I__5635 (
            .O(N__28690),
            .I(\b2v_inst11.func_state_RNI5DLRZ0Z_0 ));
    Odrv4 I__5634 (
            .O(N__28687),
            .I(\b2v_inst11.func_state_RNI5DLRZ0Z_0 ));
    CascadeMux I__5633 (
            .O(N__28680),
            .I(N__28675));
    CascadeMux I__5632 (
            .O(N__28679),
            .I(N__28672));
    CascadeMux I__5631 (
            .O(N__28678),
            .I(N__28667));
    InMux I__5630 (
            .O(N__28675),
            .I(N__28663));
    InMux I__5629 (
            .O(N__28672),
            .I(N__28658));
    InMux I__5628 (
            .O(N__28671),
            .I(N__28658));
    InMux I__5627 (
            .O(N__28670),
            .I(N__28651));
    InMux I__5626 (
            .O(N__28667),
            .I(N__28651));
    InMux I__5625 (
            .O(N__28666),
            .I(N__28651));
    LocalMux I__5624 (
            .O(N__28663),
            .I(N__28646));
    LocalMux I__5623 (
            .O(N__28658),
            .I(N__28646));
    LocalMux I__5622 (
            .O(N__28651),
            .I(N__28643));
    Span4Mux_h I__5621 (
            .O(N__28646),
            .I(N__28640));
    Span4Mux_h I__5620 (
            .O(N__28643),
            .I(N__28637));
    Odrv4 I__5619 (
            .O(N__28640),
            .I(\b2v_inst11.N_366 ));
    Odrv4 I__5618 (
            .O(N__28637),
            .I(\b2v_inst11.N_366 ));
    InMux I__5617 (
            .O(N__28632),
            .I(N__28623));
    InMux I__5616 (
            .O(N__28631),
            .I(N__28623));
    InMux I__5615 (
            .O(N__28630),
            .I(N__28618));
    InMux I__5614 (
            .O(N__28629),
            .I(N__28618));
    InMux I__5613 (
            .O(N__28628),
            .I(N__28615));
    LocalMux I__5612 (
            .O(N__28623),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ));
    LocalMux I__5611 (
            .O(N__28618),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ));
    LocalMux I__5610 (
            .O(N__28615),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ));
    InMux I__5609 (
            .O(N__28608),
            .I(N__28605));
    LocalMux I__5608 (
            .O(N__28605),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_313_N ));
    CascadeMux I__5607 (
            .O(N__28602),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2BZ0_cascade_ ));
    InMux I__5606 (
            .O(N__28599),
            .I(N__28596));
    LocalMux I__5605 (
            .O(N__28596),
            .I(\b2v_inst11.dutycycle_1_0_1 ));
    InMux I__5604 (
            .O(N__28593),
            .I(N__28590));
    LocalMux I__5603 (
            .O(N__28590),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    InMux I__5602 (
            .O(N__28587),
            .I(N__28584));
    LocalMux I__5601 (
            .O(N__28584),
            .I(N__28581));
    Span4Mux_v I__5600 (
            .O(N__28581),
            .I(N__28576));
    InMux I__5599 (
            .O(N__28580),
            .I(N__28573));
    InMux I__5598 (
            .O(N__28579),
            .I(N__28570));
    Odrv4 I__5597 (
            .O(N__28576),
            .I(\b2v_inst11.count_clk_RNIG510TZ0Z_5 ));
    LocalMux I__5596 (
            .O(N__28573),
            .I(\b2v_inst11.count_clk_RNIG510TZ0Z_5 ));
    LocalMux I__5595 (
            .O(N__28570),
            .I(\b2v_inst11.count_clk_RNIG510TZ0Z_5 ));
    CascadeMux I__5594 (
            .O(N__28563),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ));
    InMux I__5593 (
            .O(N__28560),
            .I(N__28557));
    LocalMux I__5592 (
            .O(N__28557),
            .I(\b2v_inst11.un1_func_state25_6_0_1 ));
    CascadeMux I__5591 (
            .O(N__28554),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_ ));
    CascadeMux I__5590 (
            .O(N__28551),
            .I(N__28540));
    CascadeMux I__5589 (
            .O(N__28550),
            .I(N__28537));
    CascadeMux I__5588 (
            .O(N__28549),
            .I(N__28534));
    CEMux I__5587 (
            .O(N__28548),
            .I(N__28528));
    CEMux I__5586 (
            .O(N__28547),
            .I(N__28521));
    InMux I__5585 (
            .O(N__28546),
            .I(N__28512));
    InMux I__5584 (
            .O(N__28545),
            .I(N__28512));
    InMux I__5583 (
            .O(N__28544),
            .I(N__28512));
    InMux I__5582 (
            .O(N__28543),
            .I(N__28512));
    InMux I__5581 (
            .O(N__28540),
            .I(N__28503));
    InMux I__5580 (
            .O(N__28537),
            .I(N__28503));
    InMux I__5579 (
            .O(N__28534),
            .I(N__28503));
    InMux I__5578 (
            .O(N__28533),
            .I(N__28503));
    CEMux I__5577 (
            .O(N__28532),
            .I(N__28495));
    CEMux I__5576 (
            .O(N__28531),
            .I(N__28492));
    LocalMux I__5575 (
            .O(N__28528),
            .I(N__28489));
    InMux I__5574 (
            .O(N__28527),
            .I(N__28482));
    InMux I__5573 (
            .O(N__28526),
            .I(N__28482));
    InMux I__5572 (
            .O(N__28525),
            .I(N__28482));
    CEMux I__5571 (
            .O(N__28524),
            .I(N__28479));
    LocalMux I__5570 (
            .O(N__28521),
            .I(N__28472));
    LocalMux I__5569 (
            .O(N__28512),
            .I(N__28472));
    LocalMux I__5568 (
            .O(N__28503),
            .I(N__28472));
    InMux I__5567 (
            .O(N__28502),
            .I(N__28469));
    InMux I__5566 (
            .O(N__28501),
            .I(N__28464));
    InMux I__5565 (
            .O(N__28500),
            .I(N__28464));
    InMux I__5564 (
            .O(N__28499),
            .I(N__28459));
    InMux I__5563 (
            .O(N__28498),
            .I(N__28459));
    LocalMux I__5562 (
            .O(N__28495),
            .I(N__28456));
    LocalMux I__5561 (
            .O(N__28492),
            .I(N__28453));
    Span4Mux_v I__5560 (
            .O(N__28489),
            .I(N__28450));
    LocalMux I__5559 (
            .O(N__28482),
            .I(N__28447));
    LocalMux I__5558 (
            .O(N__28479),
            .I(N__28436));
    Span4Mux_v I__5557 (
            .O(N__28472),
            .I(N__28436));
    LocalMux I__5556 (
            .O(N__28469),
            .I(N__28436));
    LocalMux I__5555 (
            .O(N__28464),
            .I(N__28436));
    LocalMux I__5554 (
            .O(N__28459),
            .I(N__28436));
    Span4Mux_h I__5553 (
            .O(N__28456),
            .I(N__28433));
    Span4Mux_h I__5552 (
            .O(N__28453),
            .I(N__28428));
    Span4Mux_h I__5551 (
            .O(N__28450),
            .I(N__28428));
    Span4Mux_h I__5550 (
            .O(N__28447),
            .I(N__28425));
    Span4Mux_h I__5549 (
            .O(N__28436),
            .I(N__28422));
    Odrv4 I__5548 (
            .O(N__28433),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__5547 (
            .O(N__28428),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__5546 (
            .O(N__28425),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__5545 (
            .O(N__28422),
            .I(\b2v_inst11.count_off_enZ0 ));
    CascadeMux I__5544 (
            .O(N__28413),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_ ));
    CascadeMux I__5543 (
            .O(N__28410),
            .I(N__28384));
    InMux I__5542 (
            .O(N__28409),
            .I(N__28379));
    InMux I__5541 (
            .O(N__28408),
            .I(N__28372));
    InMux I__5540 (
            .O(N__28407),
            .I(N__28372));
    InMux I__5539 (
            .O(N__28406),
            .I(N__28372));
    InMux I__5538 (
            .O(N__28405),
            .I(N__28365));
    InMux I__5537 (
            .O(N__28404),
            .I(N__28365));
    InMux I__5536 (
            .O(N__28403),
            .I(N__28365));
    InMux I__5535 (
            .O(N__28402),
            .I(N__28362));
    InMux I__5534 (
            .O(N__28401),
            .I(N__28353));
    InMux I__5533 (
            .O(N__28400),
            .I(N__28353));
    InMux I__5532 (
            .O(N__28399),
            .I(N__28353));
    InMux I__5531 (
            .O(N__28398),
            .I(N__28353));
    InMux I__5530 (
            .O(N__28397),
            .I(N__28344));
    InMux I__5529 (
            .O(N__28396),
            .I(N__28344));
    InMux I__5528 (
            .O(N__28395),
            .I(N__28344));
    InMux I__5527 (
            .O(N__28394),
            .I(N__28340));
    InMux I__5526 (
            .O(N__28393),
            .I(N__28331));
    InMux I__5525 (
            .O(N__28392),
            .I(N__28331));
    InMux I__5524 (
            .O(N__28391),
            .I(N__28331));
    InMux I__5523 (
            .O(N__28390),
            .I(N__28331));
    InMux I__5522 (
            .O(N__28389),
            .I(N__28321));
    InMux I__5521 (
            .O(N__28388),
            .I(N__28314));
    InMux I__5520 (
            .O(N__28387),
            .I(N__28314));
    InMux I__5519 (
            .O(N__28384),
            .I(N__28311));
    InMux I__5518 (
            .O(N__28383),
            .I(N__28306));
    InMux I__5517 (
            .O(N__28382),
            .I(N__28306));
    LocalMux I__5516 (
            .O(N__28379),
            .I(N__28295));
    LocalMux I__5515 (
            .O(N__28372),
            .I(N__28295));
    LocalMux I__5514 (
            .O(N__28365),
            .I(N__28295));
    LocalMux I__5513 (
            .O(N__28362),
            .I(N__28295));
    LocalMux I__5512 (
            .O(N__28353),
            .I(N__28295));
    InMux I__5511 (
            .O(N__28352),
            .I(N__28290));
    InMux I__5510 (
            .O(N__28351),
            .I(N__28290));
    LocalMux I__5509 (
            .O(N__28344),
            .I(N__28287));
    InMux I__5508 (
            .O(N__28343),
            .I(N__28284));
    LocalMux I__5507 (
            .O(N__28340),
            .I(N__28279));
    LocalMux I__5506 (
            .O(N__28331),
            .I(N__28279));
    InMux I__5505 (
            .O(N__28330),
            .I(N__28274));
    InMux I__5504 (
            .O(N__28329),
            .I(N__28274));
    InMux I__5503 (
            .O(N__28328),
            .I(N__28267));
    InMux I__5502 (
            .O(N__28327),
            .I(N__28267));
    InMux I__5501 (
            .O(N__28326),
            .I(N__28267));
    CascadeMux I__5500 (
            .O(N__28325),
            .I(N__28264));
    CascadeMux I__5499 (
            .O(N__28324),
            .I(N__28261));
    LocalMux I__5498 (
            .O(N__28321),
            .I(N__28254));
    InMux I__5497 (
            .O(N__28320),
            .I(N__28249));
    InMux I__5496 (
            .O(N__28319),
            .I(N__28249));
    LocalMux I__5495 (
            .O(N__28314),
            .I(N__28242));
    LocalMux I__5494 (
            .O(N__28311),
            .I(N__28242));
    LocalMux I__5493 (
            .O(N__28306),
            .I(N__28242));
    Span4Mux_v I__5492 (
            .O(N__28295),
            .I(N__28235));
    LocalMux I__5491 (
            .O(N__28290),
            .I(N__28235));
    Span4Mux_v I__5490 (
            .O(N__28287),
            .I(N__28226));
    LocalMux I__5489 (
            .O(N__28284),
            .I(N__28226));
    Span4Mux_v I__5488 (
            .O(N__28279),
            .I(N__28226));
    LocalMux I__5487 (
            .O(N__28274),
            .I(N__28226));
    LocalMux I__5486 (
            .O(N__28267),
            .I(N__28223));
    InMux I__5485 (
            .O(N__28264),
            .I(N__28220));
    InMux I__5484 (
            .O(N__28261),
            .I(N__28215));
    InMux I__5483 (
            .O(N__28260),
            .I(N__28215));
    InMux I__5482 (
            .O(N__28259),
            .I(N__28212));
    InMux I__5481 (
            .O(N__28258),
            .I(N__28209));
    InMux I__5480 (
            .O(N__28257),
            .I(N__28206));
    Span4Mux_h I__5479 (
            .O(N__28254),
            .I(N__28203));
    LocalMux I__5478 (
            .O(N__28249),
            .I(N__28200));
    Span12Mux_s6_v I__5477 (
            .O(N__28242),
            .I(N__28197));
    InMux I__5476 (
            .O(N__28241),
            .I(N__28192));
    InMux I__5475 (
            .O(N__28240),
            .I(N__28192));
    Span4Mux_h I__5474 (
            .O(N__28235),
            .I(N__28185));
    Span4Mux_h I__5473 (
            .O(N__28226),
            .I(N__28185));
    Span4Mux_h I__5472 (
            .O(N__28223),
            .I(N__28185));
    LocalMux I__5471 (
            .O(N__28220),
            .I(N__28180));
    LocalMux I__5470 (
            .O(N__28215),
            .I(N__28180));
    LocalMux I__5469 (
            .O(N__28212),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__5468 (
            .O(N__28209),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__5467 (
            .O(N__28206),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__5466 (
            .O(N__28203),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__5465 (
            .O(N__28200),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv12 I__5464 (
            .O(N__28197),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__5463 (
            .O(N__28192),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__5462 (
            .O(N__28185),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__5461 (
            .O(N__28180),
            .I(SYNTHESIZED_WIRE_1keep_3));
    CascadeMux I__5460 (
            .O(N__28161),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6_cascade_ ));
    InMux I__5459 (
            .O(N__28158),
            .I(N__28154));
    InMux I__5458 (
            .O(N__28157),
            .I(N__28151));
    LocalMux I__5457 (
            .O(N__28154),
            .I(\b2v_inst11.N_382_N ));
    LocalMux I__5456 (
            .O(N__28151),
            .I(\b2v_inst11.N_382_N ));
    CascadeMux I__5455 (
            .O(N__28146),
            .I(N__28139));
    InMux I__5454 (
            .O(N__28145),
            .I(N__28136));
    InMux I__5453 (
            .O(N__28144),
            .I(N__28133));
    InMux I__5452 (
            .O(N__28143),
            .I(N__28130));
    InMux I__5451 (
            .O(N__28142),
            .I(N__28125));
    InMux I__5450 (
            .O(N__28139),
            .I(N__28125));
    LocalMux I__5449 (
            .O(N__28136),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    LocalMux I__5448 (
            .O(N__28133),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    LocalMux I__5447 (
            .O(N__28130),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    LocalMux I__5446 (
            .O(N__28125),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    InMux I__5445 (
            .O(N__28116),
            .I(N__28108));
    CascadeMux I__5444 (
            .O(N__28115),
            .I(N__28104));
    InMux I__5443 (
            .O(N__28114),
            .I(N__28097));
    InMux I__5442 (
            .O(N__28113),
            .I(N__28097));
    InMux I__5441 (
            .O(N__28112),
            .I(N__28097));
    InMux I__5440 (
            .O(N__28111),
            .I(N__28094));
    LocalMux I__5439 (
            .O(N__28108),
            .I(N__28091));
    InMux I__5438 (
            .O(N__28107),
            .I(N__28086));
    InMux I__5437 (
            .O(N__28104),
            .I(N__28086));
    LocalMux I__5436 (
            .O(N__28097),
            .I(N__28082));
    LocalMux I__5435 (
            .O(N__28094),
            .I(N__28079));
    Span4Mux_v I__5434 (
            .O(N__28091),
            .I(N__28073));
    LocalMux I__5433 (
            .O(N__28086),
            .I(N__28073));
    InMux I__5432 (
            .O(N__28085),
            .I(N__28070));
    Span4Mux_v I__5431 (
            .O(N__28082),
            .I(N__28067));
    Span4Mux_h I__5430 (
            .O(N__28079),
            .I(N__28064));
    InMux I__5429 (
            .O(N__28078),
            .I(N__28061));
    Odrv4 I__5428 (
            .O(N__28073),
            .I(RSMRSTn_0));
    LocalMux I__5427 (
            .O(N__28070),
            .I(RSMRSTn_0));
    Odrv4 I__5426 (
            .O(N__28067),
            .I(RSMRSTn_0));
    Odrv4 I__5425 (
            .O(N__28064),
            .I(RSMRSTn_0));
    LocalMux I__5424 (
            .O(N__28061),
            .I(RSMRSTn_0));
    CascadeMux I__5423 (
            .O(N__28050),
            .I(\b2v_inst11.g0_4_sx_cascade_ ));
    InMux I__5422 (
            .O(N__28047),
            .I(N__28044));
    LocalMux I__5421 (
            .O(N__28044),
            .I(\b2v_inst11.N_428 ));
    CascadeMux I__5420 (
            .O(N__28041),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ));
    CascadeMux I__5419 (
            .O(N__28038),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_ ));
    InMux I__5418 (
            .O(N__28035),
            .I(N__28032));
    LocalMux I__5417 (
            .O(N__28032),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0 ));
    InMux I__5416 (
            .O(N__28029),
            .I(N__28023));
    InMux I__5415 (
            .O(N__28028),
            .I(N__28023));
    LocalMux I__5414 (
            .O(N__28023),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ));
    CascadeMux I__5413 (
            .O(N__28020),
            .I(\b2v_inst11.func_state_1_m2_am_1_0_cascade_ ));
    InMux I__5412 (
            .O(N__28017),
            .I(N__28014));
    LocalMux I__5411 (
            .O(N__28014),
            .I(N__28011));
    Span4Mux_h I__5410 (
            .O(N__28011),
            .I(N__28008));
    Odrv4 I__5409 (
            .O(N__28008),
            .I(\b2v_inst11.func_state_RNINCPR4Z0Z_0 ));
    InMux I__5408 (
            .O(N__28005),
            .I(N__27998));
    InMux I__5407 (
            .O(N__28004),
            .I(N__27998));
    InMux I__5406 (
            .O(N__28003),
            .I(N__27995));
    LocalMux I__5405 (
            .O(N__27998),
            .I(\b2v_inst11.N_382 ));
    LocalMux I__5404 (
            .O(N__27995),
            .I(\b2v_inst11.N_382 ));
    InMux I__5403 (
            .O(N__27990),
            .I(N__27987));
    LocalMux I__5402 (
            .O(N__27987),
            .I(\b2v_inst11.N_315 ));
    IoInMux I__5401 (
            .O(N__27984),
            .I(N__27981));
    LocalMux I__5400 (
            .O(N__27981),
            .I(N__27978));
    Span4Mux_s3_h I__5399 (
            .O(N__27978),
            .I(N__27975));
    Span4Mux_h I__5398 (
            .O(N__27975),
            .I(N__27972));
    Span4Mux_v I__5397 (
            .O(N__27972),
            .I(N__27969));
    Odrv4 I__5396 (
            .O(N__27969),
            .I(vccst_en));
    InMux I__5395 (
            .O(N__27966),
            .I(N__27963));
    LocalMux I__5394 (
            .O(N__27963),
            .I(\b2v_inst11.count_clk_RNIZ0Z_1 ));
    InMux I__5393 (
            .O(N__27960),
            .I(N__27951));
    InMux I__5392 (
            .O(N__27959),
            .I(N__27951));
    InMux I__5391 (
            .O(N__27958),
            .I(N__27951));
    LocalMux I__5390 (
            .O(N__27951),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    InMux I__5389 (
            .O(N__27948),
            .I(N__27939));
    InMux I__5388 (
            .O(N__27947),
            .I(N__27939));
    InMux I__5387 (
            .O(N__27946),
            .I(N__27939));
    LocalMux I__5386 (
            .O(N__27939),
            .I(\b2v_inst11.N_379 ));
    CascadeMux I__5385 (
            .O(N__27936),
            .I(\b2v_inst11.count_clkZ0Z_3_cascade_ ));
    InMux I__5384 (
            .O(N__27933),
            .I(N__27930));
    LocalMux I__5383 (
            .O(N__27930),
            .I(\b2v_inst11.N_190 ));
    CascadeMux I__5382 (
            .O(N__27927),
            .I(\b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ));
    InMux I__5381 (
            .O(N__27924),
            .I(N__27921));
    LocalMux I__5380 (
            .O(N__27921),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    InMux I__5379 (
            .O(N__27918),
            .I(N__27915));
    LocalMux I__5378 (
            .O(N__27915),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0 ));
    CascadeMux I__5377 (
            .O(N__27912),
            .I(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5Z0Z_0_cascade_ ));
    InMux I__5376 (
            .O(N__27909),
            .I(N__27903));
    InMux I__5375 (
            .O(N__27908),
            .I(N__27903));
    LocalMux I__5374 (
            .O(N__27903),
            .I(\b2v_inst11.count_clk_0_3 ));
    InMux I__5373 (
            .O(N__27900),
            .I(N__27894));
    InMux I__5372 (
            .O(N__27899),
            .I(N__27894));
    LocalMux I__5371 (
            .O(N__27894),
            .I(\b2v_inst6.N_276_0 ));
    CascadeMux I__5370 (
            .O(N__27891),
            .I(\b2v_inst6.curr_state_RNIKIRD1Z0Z_0_cascade_ ));
    CascadeMux I__5369 (
            .O(N__27888),
            .I(N__27884));
    InMux I__5368 (
            .O(N__27887),
            .I(N__27879));
    InMux I__5367 (
            .O(N__27884),
            .I(N__27879));
    LocalMux I__5366 (
            .O(N__27879),
            .I(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ));
    InMux I__5365 (
            .O(N__27876),
            .I(N__27869));
    InMux I__5364 (
            .O(N__27875),
            .I(N__27869));
    InMux I__5363 (
            .O(N__27874),
            .I(N__27866));
    LocalMux I__5362 (
            .O(N__27869),
            .I(\b2v_inst6.N_2992_i ));
    LocalMux I__5361 (
            .O(N__27866),
            .I(\b2v_inst6.N_2992_i ));
    InMux I__5360 (
            .O(N__27861),
            .I(N__27855));
    InMux I__5359 (
            .O(N__27860),
            .I(N__27848));
    InMux I__5358 (
            .O(N__27859),
            .I(N__27848));
    InMux I__5357 (
            .O(N__27858),
            .I(N__27848));
    LocalMux I__5356 (
            .O(N__27855),
            .I(\b2v_inst6.N_3011_i ));
    LocalMux I__5355 (
            .O(N__27848),
            .I(\b2v_inst6.N_3011_i ));
    InMux I__5354 (
            .O(N__27843),
            .I(N__27834));
    InMux I__5353 (
            .O(N__27842),
            .I(N__27834));
    InMux I__5352 (
            .O(N__27841),
            .I(N__27834));
    LocalMux I__5351 (
            .O(N__27834),
            .I(N__27831));
    Odrv4 I__5350 (
            .O(N__27831),
            .I(\b2v_inst6.N_192 ));
    CascadeMux I__5349 (
            .O(N__27828),
            .I(\b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ));
    CascadeMux I__5348 (
            .O(N__27825),
            .I(\b2v_inst11.count_clkZ0Z_0_cascade_ ));
    CascadeMux I__5347 (
            .O(N__27822),
            .I(\b2v_inst11.count_clk_RNIZ0Z_1_cascade_ ));
    CascadeMux I__5346 (
            .O(N__27819),
            .I(\b2v_inst11.un1_count_clk_2_axb_1_cascade_ ));
    InMux I__5345 (
            .O(N__27816),
            .I(N__27813));
    LocalMux I__5344 (
            .O(N__27813),
            .I(\b2v_inst11.count_clk_0_0 ));
    InMux I__5343 (
            .O(N__27810),
            .I(N__27804));
    InMux I__5342 (
            .O(N__27809),
            .I(N__27804));
    LocalMux I__5341 (
            .O(N__27804),
            .I(\b2v_inst11.count_clk_0_1 ));
    InMux I__5340 (
            .O(N__27801),
            .I(N__27798));
    LocalMux I__5339 (
            .O(N__27798),
            .I(\b2v_inst6.curr_state_1_0 ));
    CascadeMux I__5338 (
            .O(N__27795),
            .I(\b2v_inst6.curr_state_7_0_cascade_ ));
    CascadeMux I__5337 (
            .O(N__27792),
            .I(\b2v_inst6.count_RNICV5H1Z0Z_0_cascade_ ));
    CascadeMux I__5336 (
            .O(N__27789),
            .I(\b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ));
    InMux I__5335 (
            .O(N__27786),
            .I(N__27783));
    LocalMux I__5334 (
            .O(N__27783),
            .I(N__27779));
    CascadeMux I__5333 (
            .O(N__27782),
            .I(N__27774));
    Span4Mux_h I__5332 (
            .O(N__27779),
            .I(N__27771));
    InMux I__5331 (
            .O(N__27778),
            .I(N__27766));
    InMux I__5330 (
            .O(N__27777),
            .I(N__27766));
    InMux I__5329 (
            .O(N__27774),
            .I(N__27763));
    Span4Mux_v I__5328 (
            .O(N__27771),
            .I(N__27754));
    LocalMux I__5327 (
            .O(N__27766),
            .I(N__27754));
    LocalMux I__5326 (
            .O(N__27763),
            .I(N__27754));
    InMux I__5325 (
            .O(N__27762),
            .I(N__27749));
    InMux I__5324 (
            .O(N__27761),
            .I(N__27749));
    Span4Mux_v I__5323 (
            .O(N__27754),
            .I(N__27744));
    LocalMux I__5322 (
            .O(N__27749),
            .I(N__27744));
    Span4Mux_h I__5321 (
            .O(N__27744),
            .I(N__27741));
    Odrv4 I__5320 (
            .O(N__27741),
            .I(N_222));
    CascadeMux I__5319 (
            .O(N__27738),
            .I(\b2v_inst6.N_2992_i_cascade_ ));
    CascadeMux I__5318 (
            .O(N__27735),
            .I(N__27727));
    InMux I__5317 (
            .O(N__27734),
            .I(N__27718));
    InMux I__5316 (
            .O(N__27733),
            .I(N__27718));
    InMux I__5315 (
            .O(N__27732),
            .I(N__27718));
    InMux I__5314 (
            .O(N__27731),
            .I(N__27718));
    InMux I__5313 (
            .O(N__27730),
            .I(N__27715));
    InMux I__5312 (
            .O(N__27727),
            .I(N__27712));
    LocalMux I__5311 (
            .O(N__27718),
            .I(SYNTHESIZED_WIRE_8));
    LocalMux I__5310 (
            .O(N__27715),
            .I(SYNTHESIZED_WIRE_8));
    LocalMux I__5309 (
            .O(N__27712),
            .I(SYNTHESIZED_WIRE_8));
    InMux I__5308 (
            .O(N__27705),
            .I(N__27702));
    LocalMux I__5307 (
            .O(N__27702),
            .I(N__27699));
    IoSpan4Mux I__5306 (
            .O(N__27699),
            .I(N__27696));
    Odrv4 I__5305 (
            .O(N__27696),
            .I(v5s_ok));
    InMux I__5304 (
            .O(N__27693),
            .I(N__27690));
    LocalMux I__5303 (
            .O(N__27690),
            .I(N__27687));
    Span4Mux_v I__5302 (
            .O(N__27687),
            .I(N__27684));
    Span4Mux_v I__5301 (
            .O(N__27684),
            .I(N__27681));
    Span4Mux_v I__5300 (
            .O(N__27681),
            .I(N__27678));
    Odrv4 I__5299 (
            .O(N__27678),
            .I(v33s_ok));
    IoInMux I__5298 (
            .O(N__27675),
            .I(N__27672));
    LocalMux I__5297 (
            .O(N__27672),
            .I(N__27669));
    Span4Mux_s2_v I__5296 (
            .O(N__27669),
            .I(N__27665));
    IoInMux I__5295 (
            .O(N__27668),
            .I(N__27662));
    Span4Mux_v I__5294 (
            .O(N__27665),
            .I(N__27659));
    LocalMux I__5293 (
            .O(N__27662),
            .I(N__27656));
    Span4Mux_v I__5292 (
            .O(N__27659),
            .I(N__27653));
    Span4Mux_s3_h I__5291 (
            .O(N__27656),
            .I(N__27650));
    Odrv4 I__5290 (
            .O(N__27653),
            .I(vccinaux_en));
    Odrv4 I__5289 (
            .O(N__27650),
            .I(vccinaux_en));
    InMux I__5288 (
            .O(N__27645),
            .I(N__27642));
    LocalMux I__5287 (
            .O(N__27642),
            .I(N__27637));
    InMux I__5286 (
            .O(N__27641),
            .I(N__27632));
    InMux I__5285 (
            .O(N__27640),
            .I(N__27632));
    Odrv4 I__5284 (
            .O(N__27637),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    LocalMux I__5283 (
            .O(N__27632),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    InMux I__5282 (
            .O(N__27627),
            .I(N__27622));
    InMux I__5281 (
            .O(N__27626),
            .I(N__27619));
    InMux I__5280 (
            .O(N__27625),
            .I(N__27616));
    LocalMux I__5279 (
            .O(N__27622),
            .I(\b2v_inst6.curr_state_RNIKIRD1Z0Z_0 ));
    LocalMux I__5278 (
            .O(N__27619),
            .I(\b2v_inst6.curr_state_RNIKIRD1Z0Z_0 ));
    LocalMux I__5277 (
            .O(N__27616),
            .I(\b2v_inst6.curr_state_RNIKIRD1Z0Z_0 ));
    CascadeMux I__5276 (
            .O(N__27609),
            .I(\b2v_inst6.un2_count_1_axb_9_cascade_ ));
    InMux I__5275 (
            .O(N__27606),
            .I(N__27600));
    InMux I__5274 (
            .O(N__27605),
            .I(N__27600));
    LocalMux I__5273 (
            .O(N__27600),
            .I(\b2v_inst6.count_rst_6 ));
    InMux I__5272 (
            .O(N__27597),
            .I(N__27591));
    InMux I__5271 (
            .O(N__27596),
            .I(N__27591));
    LocalMux I__5270 (
            .O(N__27591),
            .I(\b2v_inst6.count_rst_5 ));
    CascadeMux I__5269 (
            .O(N__27588),
            .I(\b2v_inst6.countZ0Z_8_cascade_ ));
    InMux I__5268 (
            .O(N__27585),
            .I(N__27579));
    InMux I__5267 (
            .O(N__27584),
            .I(N__27579));
    LocalMux I__5266 (
            .O(N__27579),
            .I(\b2v_inst6.count_0_9 ));
    InMux I__5265 (
            .O(N__27576),
            .I(N__27570));
    InMux I__5264 (
            .O(N__27575),
            .I(N__27570));
    LocalMux I__5263 (
            .O(N__27570),
            .I(\b2v_inst6.count_0_8 ));
    InMux I__5262 (
            .O(N__27567),
            .I(N__27559));
    InMux I__5261 (
            .O(N__27566),
            .I(N__27552));
    InMux I__5260 (
            .O(N__27565),
            .I(N__27552));
    InMux I__5259 (
            .O(N__27564),
            .I(N__27552));
    InMux I__5258 (
            .O(N__27563),
            .I(N__27547));
    InMux I__5257 (
            .O(N__27562),
            .I(N__27547));
    LocalMux I__5256 (
            .O(N__27559),
            .I(N__27530));
    LocalMux I__5255 (
            .O(N__27552),
            .I(N__27527));
    LocalMux I__5254 (
            .O(N__27547),
            .I(N__27524));
    CEMux I__5253 (
            .O(N__27546),
            .I(N__27489));
    CEMux I__5252 (
            .O(N__27545),
            .I(N__27489));
    CEMux I__5251 (
            .O(N__27544),
            .I(N__27489));
    CEMux I__5250 (
            .O(N__27543),
            .I(N__27489));
    CEMux I__5249 (
            .O(N__27542),
            .I(N__27489));
    CEMux I__5248 (
            .O(N__27541),
            .I(N__27489));
    CEMux I__5247 (
            .O(N__27540),
            .I(N__27489));
    CEMux I__5246 (
            .O(N__27539),
            .I(N__27489));
    CEMux I__5245 (
            .O(N__27538),
            .I(N__27489));
    CEMux I__5244 (
            .O(N__27537),
            .I(N__27489));
    CEMux I__5243 (
            .O(N__27536),
            .I(N__27489));
    CEMux I__5242 (
            .O(N__27535),
            .I(N__27489));
    CEMux I__5241 (
            .O(N__27534),
            .I(N__27489));
    CEMux I__5240 (
            .O(N__27533),
            .I(N__27489));
    Glb2LocalMux I__5239 (
            .O(N__27530),
            .I(N__27489));
    Glb2LocalMux I__5238 (
            .O(N__27527),
            .I(N__27489));
    Glb2LocalMux I__5237 (
            .O(N__27524),
            .I(N__27489));
    GlobalMux I__5236 (
            .O(N__27489),
            .I(N__27486));
    gio2CtrlBuf I__5235 (
            .O(N__27486),
            .I(N_607_g));
    CascadeMux I__5234 (
            .O(N__27483),
            .I(\b2v_inst6.N_394_cascade_ ));
    InMux I__5233 (
            .O(N__27480),
            .I(N__27477));
    LocalMux I__5232 (
            .O(N__27477),
            .I(N__27474));
    Odrv4 I__5231 (
            .O(N__27474),
            .I(\b2v_inst6.curr_state_1_1 ));
    CascadeMux I__5230 (
            .O(N__27471),
            .I(\b2v_inst6.m6_i_a3_cascade_ ));
    CascadeMux I__5229 (
            .O(N__27468),
            .I(N__27462));
    InMux I__5228 (
            .O(N__27467),
            .I(N__27457));
    InMux I__5227 (
            .O(N__27466),
            .I(N__27457));
    InMux I__5226 (
            .O(N__27465),
            .I(N__27452));
    InMux I__5225 (
            .O(N__27462),
            .I(N__27452));
    LocalMux I__5224 (
            .O(N__27457),
            .I(N__27449));
    LocalMux I__5223 (
            .O(N__27452),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    Odrv4 I__5222 (
            .O(N__27449),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    CascadeMux I__5221 (
            .O(N__27444),
            .I(\b2v_inst6.curr_stateZ0Z_1_cascade_ ));
    InMux I__5220 (
            .O(N__27441),
            .I(\b2v_inst11.CO2 ));
    CascadeMux I__5219 (
            .O(N__27438),
            .I(N__27434));
    InMux I__5218 (
            .O(N__27437),
            .I(N__27431));
    InMux I__5217 (
            .O(N__27434),
            .I(N__27428));
    LocalMux I__5216 (
            .O(N__27431),
            .I(\b2v_inst11.mult1_un61_sum ));
    LocalMux I__5215 (
            .O(N__27428),
            .I(\b2v_inst11.mult1_un61_sum ));
    InMux I__5214 (
            .O(N__27423),
            .I(N__27420));
    LocalMux I__5213 (
            .O(N__27420),
            .I(\b2v_inst11.mult1_un61_sum_i ));
    CascadeMux I__5212 (
            .O(N__27417),
            .I(N__27414));
    InMux I__5211 (
            .O(N__27414),
            .I(N__27411));
    LocalMux I__5210 (
            .O(N__27411),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_13 ));
    InMux I__5209 (
            .O(N__27408),
            .I(N__27404));
    InMux I__5208 (
            .O(N__27407),
            .I(N__27401));
    LocalMux I__5207 (
            .O(N__27404),
            .I(N__27398));
    LocalMux I__5206 (
            .O(N__27401),
            .I(\b2v_inst11.mult1_un47_sum_6 ));
    Odrv4 I__5205 (
            .O(N__27398),
            .I(\b2v_inst11.mult1_un47_sum_6 ));
    CascadeMux I__5204 (
            .O(N__27393),
            .I(N__27390));
    InMux I__5203 (
            .O(N__27390),
            .I(N__27386));
    InMux I__5202 (
            .O(N__27389),
            .I(N__27383));
    LocalMux I__5201 (
            .O(N__27386),
            .I(N__27380));
    LocalMux I__5200 (
            .O(N__27383),
            .I(\b2v_inst11.mult1_un89_sum ));
    Odrv12 I__5199 (
            .O(N__27380),
            .I(\b2v_inst11.mult1_un89_sum ));
    InMux I__5198 (
            .O(N__27375),
            .I(N__27372));
    LocalMux I__5197 (
            .O(N__27372),
            .I(N__27369));
    Odrv4 I__5196 (
            .O(N__27369),
            .I(\b2v_inst11.mult1_un89_sum_i ));
    CascadeMux I__5195 (
            .O(N__27366),
            .I(\b2v_inst6.un2_count_1_axb_8_cascade_ ));
    InMux I__5194 (
            .O(N__27363),
            .I(bfn_8_15_0_));
    InMux I__5193 (
            .O(N__27360),
            .I(N__27356));
    InMux I__5192 (
            .O(N__27359),
            .I(N__27353));
    LocalMux I__5191 (
            .O(N__27356),
            .I(N__27348));
    LocalMux I__5190 (
            .O(N__27353),
            .I(N__27348));
    Span4Mux_v I__5189 (
            .O(N__27348),
            .I(N__27345));
    Odrv4 I__5188 (
            .O(N__27345),
            .I(\b2v_inst11.mult1_un82_sum ));
    InMux I__5187 (
            .O(N__27342),
            .I(\b2v_inst11.un1_dutycycle_53_cry_8 ));
    InMux I__5186 (
            .O(N__27339),
            .I(N__27336));
    LocalMux I__5185 (
            .O(N__27336),
            .I(N__27332));
    InMux I__5184 (
            .O(N__27335),
            .I(N__27329));
    Span4Mux_v I__5183 (
            .O(N__27332),
            .I(N__27326));
    LocalMux I__5182 (
            .O(N__27329),
            .I(N__27323));
    Odrv4 I__5181 (
            .O(N__27326),
            .I(\b2v_inst11.mult1_un75_sum ));
    Odrv4 I__5180 (
            .O(N__27323),
            .I(\b2v_inst11.mult1_un75_sum ));
    InMux I__5179 (
            .O(N__27318),
            .I(\b2v_inst11.un1_dutycycle_53_cry_9 ));
    InMux I__5178 (
            .O(N__27315),
            .I(N__27312));
    LocalMux I__5177 (
            .O(N__27312),
            .I(N__27308));
    CascadeMux I__5176 (
            .O(N__27311),
            .I(N__27305));
    Span4Mux_v I__5175 (
            .O(N__27308),
            .I(N__27302));
    InMux I__5174 (
            .O(N__27305),
            .I(N__27299));
    Odrv4 I__5173 (
            .O(N__27302),
            .I(\b2v_inst11.mult1_un68_sum ));
    LocalMux I__5172 (
            .O(N__27299),
            .I(\b2v_inst11.mult1_un68_sum ));
    InMux I__5171 (
            .O(N__27294),
            .I(\b2v_inst11.un1_dutycycle_53_cry_10 ));
    InMux I__5170 (
            .O(N__27291),
            .I(\b2v_inst11.un1_dutycycle_53_cry_11 ));
    CascadeMux I__5169 (
            .O(N__27288),
            .I(N__27285));
    InMux I__5168 (
            .O(N__27285),
            .I(N__27281));
    CascadeMux I__5167 (
            .O(N__27284),
            .I(N__27278));
    LocalMux I__5166 (
            .O(N__27281),
            .I(N__27275));
    InMux I__5165 (
            .O(N__27278),
            .I(N__27272));
    Odrv4 I__5164 (
            .O(N__27275),
            .I(\b2v_inst11.mult1_un47_sum_1 ));
    LocalMux I__5163 (
            .O(N__27272),
            .I(\b2v_inst11.mult1_un47_sum_1 ));
    InMux I__5162 (
            .O(N__27267),
            .I(\b2v_inst11.un1_dutycycle_53_cry_12 ));
    InMux I__5161 (
            .O(N__27264),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13 ));
    InMux I__5160 (
            .O(N__27261),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14 ));
    InMux I__5159 (
            .O(N__27258),
            .I(bfn_8_16_0_));
    CascadeMux I__5158 (
            .O(N__27255),
            .I(N__27252));
    InMux I__5157 (
            .O(N__27252),
            .I(N__27249));
    LocalMux I__5156 (
            .O(N__27249),
            .I(N__27245));
    InMux I__5155 (
            .O(N__27248),
            .I(N__27242));
    Span4Mux_h I__5154 (
            .O(N__27245),
            .I(N__27239));
    LocalMux I__5153 (
            .O(N__27242),
            .I(\b2v_inst11.un1_dutycycle_53_axb_0 ));
    Odrv4 I__5152 (
            .O(N__27239),
            .I(\b2v_inst11.un1_dutycycle_53_axb_0 ));
    CascadeMux I__5151 (
            .O(N__27234),
            .I(N__27231));
    InMux I__5150 (
            .O(N__27231),
            .I(N__27228));
    LocalMux I__5149 (
            .O(N__27228),
            .I(N__27225));
    Odrv12 I__5148 (
            .O(N__27225),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_0 ));
    InMux I__5147 (
            .O(N__27222),
            .I(N__27218));
    InMux I__5146 (
            .O(N__27221),
            .I(N__27215));
    LocalMux I__5145 (
            .O(N__27218),
            .I(N__27212));
    LocalMux I__5144 (
            .O(N__27215),
            .I(N__27209));
    Span4Mux_v I__5143 (
            .O(N__27212),
            .I(N__27206));
    Span4Mux_v I__5142 (
            .O(N__27209),
            .I(N__27203));
    Span4Mux_h I__5141 (
            .O(N__27206),
            .I(N__27200));
    Odrv4 I__5140 (
            .O(N__27203),
            .I(\b2v_inst11.mult1_un138_sum ));
    Odrv4 I__5139 (
            .O(N__27200),
            .I(\b2v_inst11.mult1_un138_sum ));
    InMux I__5138 (
            .O(N__27195),
            .I(\b2v_inst11.un1_dutycycle_53_cry_0 ));
    InMux I__5137 (
            .O(N__27192),
            .I(N__27189));
    LocalMux I__5136 (
            .O(N__27189),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_2 ));
    InMux I__5135 (
            .O(N__27186),
            .I(N__27182));
    InMux I__5134 (
            .O(N__27185),
            .I(N__27179));
    LocalMux I__5133 (
            .O(N__27182),
            .I(N__27176));
    LocalMux I__5132 (
            .O(N__27179),
            .I(N__27173));
    Span4Mux_s2_v I__5131 (
            .O(N__27176),
            .I(N__27170));
    Odrv4 I__5130 (
            .O(N__27173),
            .I(\b2v_inst11.mult1_un131_sum ));
    Odrv4 I__5129 (
            .O(N__27170),
            .I(\b2v_inst11.mult1_un131_sum ));
    InMux I__5128 (
            .O(N__27165),
            .I(\b2v_inst11.un1_dutycycle_53_cry_1 ));
    CascadeMux I__5127 (
            .O(N__27162),
            .I(N__27159));
    InMux I__5126 (
            .O(N__27159),
            .I(N__27156));
    LocalMux I__5125 (
            .O(N__27156),
            .I(N__27153));
    Span4Mux_v I__5124 (
            .O(N__27153),
            .I(N__27150));
    Odrv4 I__5123 (
            .O(N__27150),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_2 ));
    InMux I__5122 (
            .O(N__27147),
            .I(N__27143));
    InMux I__5121 (
            .O(N__27146),
            .I(N__27140));
    LocalMux I__5120 (
            .O(N__27143),
            .I(N__27137));
    LocalMux I__5119 (
            .O(N__27140),
            .I(N__27134));
    Span4Mux_v I__5118 (
            .O(N__27137),
            .I(N__27129));
    Span4Mux_s2_v I__5117 (
            .O(N__27134),
            .I(N__27129));
    Odrv4 I__5116 (
            .O(N__27129),
            .I(\b2v_inst11.mult1_un124_sum ));
    InMux I__5115 (
            .O(N__27126),
            .I(\b2v_inst11.un1_dutycycle_53_cry_2 ));
    CascadeMux I__5114 (
            .O(N__27123),
            .I(N__27120));
    InMux I__5113 (
            .O(N__27120),
            .I(N__27117));
    LocalMux I__5112 (
            .O(N__27117),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5 ));
    InMux I__5111 (
            .O(N__27114),
            .I(N__27111));
    LocalMux I__5110 (
            .O(N__27111),
            .I(N__27107));
    InMux I__5109 (
            .O(N__27110),
            .I(N__27104));
    Span4Mux_s2_v I__5108 (
            .O(N__27107),
            .I(N__27101));
    LocalMux I__5107 (
            .O(N__27104),
            .I(N__27098));
    Odrv4 I__5106 (
            .O(N__27101),
            .I(\b2v_inst11.mult1_un117_sum ));
    Odrv12 I__5105 (
            .O(N__27098),
            .I(\b2v_inst11.mult1_un117_sum ));
    InMux I__5104 (
            .O(N__27093),
            .I(\b2v_inst11.un1_dutycycle_53_cry_3 ));
    InMux I__5103 (
            .O(N__27090),
            .I(N__27087));
    LocalMux I__5102 (
            .O(N__27087),
            .I(N__27083));
    InMux I__5101 (
            .O(N__27086),
            .I(N__27080));
    Span4Mux_v I__5100 (
            .O(N__27083),
            .I(N__27075));
    LocalMux I__5099 (
            .O(N__27080),
            .I(N__27075));
    Odrv4 I__5098 (
            .O(N__27075),
            .I(\b2v_inst11.mult1_un110_sum ));
    InMux I__5097 (
            .O(N__27072),
            .I(\b2v_inst11.un1_dutycycle_53_cry_4 ));
    InMux I__5096 (
            .O(N__27069),
            .I(N__27065));
    InMux I__5095 (
            .O(N__27068),
            .I(N__27062));
    LocalMux I__5094 (
            .O(N__27065),
            .I(N__27059));
    LocalMux I__5093 (
            .O(N__27062),
            .I(N__27056));
    Span4Mux_s3_h I__5092 (
            .O(N__27059),
            .I(N__27053));
    Span4Mux_h I__5091 (
            .O(N__27056),
            .I(N__27050));
    Span4Mux_h I__5090 (
            .O(N__27053),
            .I(N__27047));
    Odrv4 I__5089 (
            .O(N__27050),
            .I(\b2v_inst11.mult1_un103_sum ));
    Odrv4 I__5088 (
            .O(N__27047),
            .I(\b2v_inst11.mult1_un103_sum ));
    InMux I__5087 (
            .O(N__27042),
            .I(\b2v_inst11.un1_dutycycle_53_cry_5 ));
    InMux I__5086 (
            .O(N__27039),
            .I(N__27035));
    InMux I__5085 (
            .O(N__27038),
            .I(N__27032));
    LocalMux I__5084 (
            .O(N__27035),
            .I(N__27029));
    LocalMux I__5083 (
            .O(N__27032),
            .I(N__27026));
    Span4Mux_v I__5082 (
            .O(N__27029),
            .I(N__27021));
    Span4Mux_s2_v I__5081 (
            .O(N__27026),
            .I(N__27021));
    Odrv4 I__5080 (
            .O(N__27021),
            .I(\b2v_inst11.mult1_un96_sum ));
    InMux I__5079 (
            .O(N__27018),
            .I(\b2v_inst11.un1_dutycycle_53_cry_6 ));
    InMux I__5078 (
            .O(N__27015),
            .I(N__27009));
    InMux I__5077 (
            .O(N__27014),
            .I(N__27009));
    LocalMux I__5076 (
            .O(N__27009),
            .I(\b2v_inst11.dutycycle_RNI_10Z0Z_0 ));
    CascadeMux I__5075 (
            .O(N__27006),
            .I(\b2v_inst11.dutycycle_RNIPKS23Z0Z_4_cascade_ ));
    InMux I__5074 (
            .O(N__27003),
            .I(N__27000));
    LocalMux I__5073 (
            .O(N__27000),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08UZ0 ));
    CascadeMux I__5072 (
            .O(N__26997),
            .I(N__26992));
    InMux I__5071 (
            .O(N__26996),
            .I(N__26985));
    InMux I__5070 (
            .O(N__26995),
            .I(N__26985));
    InMux I__5069 (
            .O(N__26992),
            .I(N__26985));
    LocalMux I__5068 (
            .O(N__26985),
            .I(\b2v_inst11.dutycycleZ1Z_4 ));
    InMux I__5067 (
            .O(N__26982),
            .I(N__26976));
    InMux I__5066 (
            .O(N__26981),
            .I(N__26976));
    LocalMux I__5065 (
            .O(N__26976),
            .I(\b2v_inst11.dutycycle_RNI5AV24Z0Z_4 ));
    InMux I__5064 (
            .O(N__26973),
            .I(N__26970));
    LocalMux I__5063 (
            .O(N__26970),
            .I(\b2v_inst11.dutycycle_RNIPKS23Z0Z_4 ));
    CascadeMux I__5062 (
            .O(N__26967),
            .I(\b2v_inst11.dutycycleZ0Z_6_cascade_ ));
    CascadeMux I__5061 (
            .O(N__26964),
            .I(\b2v_inst11.un1_i3_mux_cascade_ ));
    InMux I__5060 (
            .O(N__26961),
            .I(N__26958));
    LocalMux I__5059 (
            .O(N__26958),
            .I(\b2v_inst11.d_i3_mux ));
    CascadeMux I__5058 (
            .O(N__26955),
            .I(\b2v_inst11.un1_dutycycle_172_m4_rn_0_cascade_ ));
    InMux I__5057 (
            .O(N__26952),
            .I(N__26949));
    LocalMux I__5056 (
            .O(N__26949),
            .I(\b2v_inst11.un1_dutycycle_172_m4 ));
    InMux I__5055 (
            .O(N__26946),
            .I(N__26943));
    LocalMux I__5054 (
            .O(N__26943),
            .I(\b2v_inst11.N_3057_0 ));
    InMux I__5053 (
            .O(N__26940),
            .I(N__26934));
    InMux I__5052 (
            .O(N__26939),
            .I(N__26934));
    LocalMux I__5051 (
            .O(N__26934),
            .I(\b2v_inst11.g1_0_0_0 ));
    InMux I__5050 (
            .O(N__26931),
            .I(N__26928));
    LocalMux I__5049 (
            .O(N__26928),
            .I(\b2v_inst11.N_3055_0_0 ));
    CascadeMux I__5048 (
            .O(N__26925),
            .I(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_1_cascade_ ));
    InMux I__5047 (
            .O(N__26922),
            .I(N__26919));
    LocalMux I__5046 (
            .O(N__26919),
            .I(\b2v_inst11.g0_0_1 ));
    InMux I__5045 (
            .O(N__26916),
            .I(N__26910));
    InMux I__5044 (
            .O(N__26915),
            .I(N__26910));
    LocalMux I__5043 (
            .O(N__26910),
            .I(\b2v_inst11.g1_0_1_0 ));
    InMux I__5042 (
            .O(N__26907),
            .I(N__26904));
    LocalMux I__5041 (
            .O(N__26904),
            .I(\b2v_inst11.g0_3_2 ));
    CascadeMux I__5040 (
            .O(N__26901),
            .I(\b2v_inst11.g2_1_0_1_cascade_ ));
    InMux I__5039 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__5038 (
            .O(N__26895),
            .I(\b2v_inst11.g2_1_0 ));
    InMux I__5037 (
            .O(N__26892),
            .I(N__26889));
    LocalMux I__5036 (
            .O(N__26889),
            .I(\b2v_inst11.dutycycle_RNI_9Z0Z_0 ));
    CascadeMux I__5035 (
            .O(N__26886),
            .I(\b2v_inst11.un1_dutycycle_172_m3_d_ns_1_0_cascade_ ));
    InMux I__5034 (
            .O(N__26883),
            .I(N__26880));
    LocalMux I__5033 (
            .O(N__26880),
            .I(\b2v_inst11.g1_1 ));
    InMux I__5032 (
            .O(N__26877),
            .I(N__26874));
    LocalMux I__5031 (
            .O(N__26874),
            .I(\b2v_inst11.dutycycle_RNIDQ4A1Z0Z_5 ));
    CascadeMux I__5030 (
            .O(N__26871),
            .I(\b2v_inst11.un1_dutycycle_172_m4_rn_1_cascade_ ));
    InMux I__5029 (
            .O(N__26868),
            .I(N__26865));
    LocalMux I__5028 (
            .O(N__26865),
            .I(\b2v_inst11.dutycycle_RNI_11Z0Z_0 ));
    InMux I__5027 (
            .O(N__26862),
            .I(N__26856));
    InMux I__5026 (
            .O(N__26861),
            .I(N__26856));
    LocalMux I__5025 (
            .O(N__26856),
            .I(N__26851));
    InMux I__5024 (
            .O(N__26855),
            .I(N__26848));
    InMux I__5023 (
            .O(N__26854),
            .I(N__26845));
    Odrv4 I__5022 (
            .O(N__26851),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ));
    LocalMux I__5021 (
            .O(N__26848),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ));
    LocalMux I__5020 (
            .O(N__26845),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ));
    CascadeMux I__5019 (
            .O(N__26838),
            .I(\b2v_inst11.dutycycleZ1Z_5_cascade_ ));
    CascadeMux I__5018 (
            .O(N__26835),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_5_cascade_ ));
    InMux I__5017 (
            .O(N__26832),
            .I(N__26829));
    LocalMux I__5016 (
            .O(N__26829),
            .I(N__26826));
    Odrv4 I__5015 (
            .O(N__26826),
            .I(\b2v_inst11.N_293 ));
    CascadeMux I__5014 (
            .O(N__26823),
            .I(N__26820));
    InMux I__5013 (
            .O(N__26820),
            .I(N__26814));
    InMux I__5012 (
            .O(N__26819),
            .I(N__26814));
    LocalMux I__5011 (
            .O(N__26814),
            .I(N__26810));
    InMux I__5010 (
            .O(N__26813),
            .I(N__26807));
    Span4Mux_h I__5009 (
            .O(N__26810),
            .I(N__26804));
    LocalMux I__5008 (
            .O(N__26807),
            .I(\b2v_inst11.N_365 ));
    Odrv4 I__5007 (
            .O(N__26804),
            .I(\b2v_inst11.N_365 ));
    CascadeMux I__5006 (
            .O(N__26799),
            .I(\b2v_inst11.N_159_cascade_ ));
    CascadeMux I__5005 (
            .O(N__26796),
            .I(\b2v_inst11.func_state_1_m2_0_cascade_ ));
    CascadeMux I__5004 (
            .O(N__26793),
            .I(\b2v_inst11.func_stateZ0Z_0_cascade_ ));
    InMux I__5003 (
            .O(N__26790),
            .I(N__26787));
    LocalMux I__5002 (
            .O(N__26787),
            .I(\b2v_inst11.func_state_1_m2_0 ));
    InMux I__5001 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__5000 (
            .O(N__26781),
            .I(N__26778));
    Span4Mux_v I__4999 (
            .O(N__26778),
            .I(N__26770));
    InMux I__4998 (
            .O(N__26777),
            .I(N__26767));
    InMux I__4997 (
            .O(N__26776),
            .I(N__26762));
    InMux I__4996 (
            .O(N__26775),
            .I(N__26762));
    InMux I__4995 (
            .O(N__26774),
            .I(N__26757));
    InMux I__4994 (
            .O(N__26773),
            .I(N__26757));
    Odrv4 I__4993 (
            .O(N__26770),
            .I(VCCST_EN_i_0_o3_0));
    LocalMux I__4992 (
            .O(N__26767),
            .I(VCCST_EN_i_0_o3_0));
    LocalMux I__4991 (
            .O(N__26762),
            .I(VCCST_EN_i_0_o3_0));
    LocalMux I__4990 (
            .O(N__26757),
            .I(VCCST_EN_i_0_o3_0));
    InMux I__4989 (
            .O(N__26748),
            .I(N__26742));
    InMux I__4988 (
            .O(N__26747),
            .I(N__26742));
    LocalMux I__4987 (
            .O(N__26742),
            .I(\b2v_inst11.func_stateZ1Z_0 ));
    CascadeMux I__4986 (
            .O(N__26739),
            .I(N__26736));
    InMux I__4985 (
            .O(N__26736),
            .I(N__26725));
    InMux I__4984 (
            .O(N__26735),
            .I(N__26725));
    InMux I__4983 (
            .O(N__26734),
            .I(N__26725));
    InMux I__4982 (
            .O(N__26733),
            .I(N__26720));
    InMux I__4981 (
            .O(N__26732),
            .I(N__26720));
    LocalMux I__4980 (
            .O(N__26725),
            .I(\b2v_inst11.count_clk_en_0 ));
    LocalMux I__4979 (
            .O(N__26720),
            .I(\b2v_inst11.count_clk_en_0 ));
    CascadeMux I__4978 (
            .O(N__26715),
            .I(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1_cascade_ ));
    InMux I__4977 (
            .O(N__26712),
            .I(N__26709));
    LocalMux I__4976 (
            .O(N__26709),
            .I(\b2v_inst11.un1_dutycycle_53_axb_3_1 ));
    CascadeMux I__4975 (
            .O(N__26706),
            .I(N__26703));
    InMux I__4974 (
            .O(N__26703),
            .I(N__26700));
    LocalMux I__4973 (
            .O(N__26700),
            .I(\b2v_inst11.d_N_5 ));
    CascadeMux I__4972 (
            .O(N__26697),
            .I(N__26694));
    InMux I__4971 (
            .O(N__26694),
            .I(N__26682));
    InMux I__4970 (
            .O(N__26693),
            .I(N__26682));
    InMux I__4969 (
            .O(N__26692),
            .I(N__26682));
    InMux I__4968 (
            .O(N__26691),
            .I(N__26682));
    LocalMux I__4967 (
            .O(N__26682),
            .I(N__26677));
    InMux I__4966 (
            .O(N__26681),
            .I(N__26674));
    CascadeMux I__4965 (
            .O(N__26680),
            .I(N__26666));
    Span4Mux_h I__4964 (
            .O(N__26677),
            .I(N__26661));
    LocalMux I__4963 (
            .O(N__26674),
            .I(N__26661));
    InMux I__4962 (
            .O(N__26673),
            .I(N__26658));
    CascadeMux I__4961 (
            .O(N__26672),
            .I(N__26655));
    InMux I__4960 (
            .O(N__26671),
            .I(N__26645));
    InMux I__4959 (
            .O(N__26670),
            .I(N__26645));
    InMux I__4958 (
            .O(N__26669),
            .I(N__26645));
    InMux I__4957 (
            .O(N__26666),
            .I(N__26645));
    Span4Mux_h I__4956 (
            .O(N__26661),
            .I(N__26640));
    LocalMux I__4955 (
            .O(N__26658),
            .I(N__26640));
    InMux I__4954 (
            .O(N__26655),
            .I(N__26635));
    InMux I__4953 (
            .O(N__26654),
            .I(N__26635));
    LocalMux I__4952 (
            .O(N__26645),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv4 I__4951 (
            .O(N__26640),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    LocalMux I__4950 (
            .O(N__26635),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    InMux I__4949 (
            .O(N__26628),
            .I(N__26622));
    InMux I__4948 (
            .O(N__26627),
            .I(N__26622));
    LocalMux I__4947 (
            .O(N__26622),
            .I(\b2v_inst11.func_state_1_ss0_i_0_o3_0 ));
    InMux I__4946 (
            .O(N__26619),
            .I(N__26616));
    LocalMux I__4945 (
            .O(N__26616),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_331_N ));
    CascadeMux I__4944 (
            .O(N__26613),
            .I(\b2v_inst11.un1_func_state25_6_0_a3_0_1_cascade_ ));
    InMux I__4943 (
            .O(N__26610),
            .I(N__26607));
    LocalMux I__4942 (
            .O(N__26607),
            .I(N__26604));
    Odrv4 I__4941 (
            .O(N__26604),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_332_N ));
    CascadeMux I__4940 (
            .O(N__26601),
            .I(N__26598));
    InMux I__4939 (
            .O(N__26598),
            .I(N__26594));
    InMux I__4938 (
            .O(N__26597),
            .I(N__26591));
    LocalMux I__4937 (
            .O(N__26594),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    LocalMux I__4936 (
            .O(N__26591),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    CascadeMux I__4935 (
            .O(N__26586),
            .I(\b2v_inst11.N_337_cascade_ ));
    InMux I__4934 (
            .O(N__26583),
            .I(N__26580));
    LocalMux I__4933 (
            .O(N__26580),
            .I(\b2v_inst11.func_state_1_m2s2_i_1 ));
    InMux I__4932 (
            .O(N__26577),
            .I(N__26574));
    LocalMux I__4931 (
            .O(N__26574),
            .I(\b2v_inst11.N_76 ));
    InMux I__4930 (
            .O(N__26571),
            .I(N__26568));
    LocalMux I__4929 (
            .O(N__26568),
            .I(\b2v_inst11.func_state_RNI6IFF4_0Z0Z_1 ));
    CascadeMux I__4928 (
            .O(N__26565),
            .I(\b2v_inst11.N_428_cascade_ ));
    InMux I__4927 (
            .O(N__26562),
            .I(N__26559));
    LocalMux I__4926 (
            .O(N__26559),
            .I(\b2v_inst11.count_clk_RNITV5AUZ0Z_7 ));
    CascadeMux I__4925 (
            .O(N__26556),
            .I(N__26549));
    CascadeMux I__4924 (
            .O(N__26555),
            .I(N__26544));
    CascadeMux I__4923 (
            .O(N__26554),
            .I(N__26541));
    CascadeMux I__4922 (
            .O(N__26553),
            .I(N__26538));
    InMux I__4921 (
            .O(N__26552),
            .I(N__26517));
    InMux I__4920 (
            .O(N__26549),
            .I(N__26517));
    InMux I__4919 (
            .O(N__26548),
            .I(N__26506));
    InMux I__4918 (
            .O(N__26547),
            .I(N__26506));
    InMux I__4917 (
            .O(N__26544),
            .I(N__26506));
    InMux I__4916 (
            .O(N__26541),
            .I(N__26506));
    InMux I__4915 (
            .O(N__26538),
            .I(N__26506));
    InMux I__4914 (
            .O(N__26537),
            .I(N__26489));
    InMux I__4913 (
            .O(N__26536),
            .I(N__26489));
    InMux I__4912 (
            .O(N__26535),
            .I(N__26489));
    InMux I__4911 (
            .O(N__26534),
            .I(N__26489));
    InMux I__4910 (
            .O(N__26533),
            .I(N__26489));
    InMux I__4909 (
            .O(N__26532),
            .I(N__26489));
    InMux I__4908 (
            .O(N__26531),
            .I(N__26489));
    InMux I__4907 (
            .O(N__26530),
            .I(N__26489));
    InMux I__4906 (
            .O(N__26529),
            .I(N__26474));
    InMux I__4905 (
            .O(N__26528),
            .I(N__26474));
    InMux I__4904 (
            .O(N__26527),
            .I(N__26474));
    InMux I__4903 (
            .O(N__26526),
            .I(N__26474));
    InMux I__4902 (
            .O(N__26525),
            .I(N__26474));
    InMux I__4901 (
            .O(N__26524),
            .I(N__26474));
    InMux I__4900 (
            .O(N__26523),
            .I(N__26474));
    CascadeMux I__4899 (
            .O(N__26522),
            .I(N__26468));
    LocalMux I__4898 (
            .O(N__26517),
            .I(N__26461));
    LocalMux I__4897 (
            .O(N__26506),
            .I(N__26461));
    LocalMux I__4896 (
            .O(N__26489),
            .I(N__26452));
    LocalMux I__4895 (
            .O(N__26474),
            .I(N__26452));
    InMux I__4894 (
            .O(N__26473),
            .I(N__26439));
    InMux I__4893 (
            .O(N__26472),
            .I(N__26439));
    InMux I__4892 (
            .O(N__26471),
            .I(N__26439));
    InMux I__4891 (
            .O(N__26468),
            .I(N__26439));
    InMux I__4890 (
            .O(N__26467),
            .I(N__26439));
    InMux I__4889 (
            .O(N__26466),
            .I(N__26439));
    Span4Mux_h I__4888 (
            .O(N__26461),
            .I(N__26436));
    InMux I__4887 (
            .O(N__26460),
            .I(N__26427));
    InMux I__4886 (
            .O(N__26459),
            .I(N__26427));
    InMux I__4885 (
            .O(N__26458),
            .I(N__26427));
    InMux I__4884 (
            .O(N__26457),
            .I(N__26427));
    Span4Mux_h I__4883 (
            .O(N__26452),
            .I(N__26424));
    LocalMux I__4882 (
            .O(N__26439),
            .I(N__26421));
    Odrv4 I__4881 (
            .O(N__26436),
            .I(\b2v_inst11.count_clk_RNILG61T1Z0Z_5 ));
    LocalMux I__4880 (
            .O(N__26427),
            .I(\b2v_inst11.count_clk_RNILG61T1Z0Z_5 ));
    Odrv4 I__4879 (
            .O(N__26424),
            .I(\b2v_inst11.count_clk_RNILG61T1Z0Z_5 ));
    Odrv4 I__4878 (
            .O(N__26421),
            .I(\b2v_inst11.count_clk_RNILG61T1Z0Z_5 ));
    CascadeMux I__4877 (
            .O(N__26412),
            .I(\b2v_inst11.un1_func_state25_4_i_a2_sxZ0_cascade_ ));
    CascadeMux I__4876 (
            .O(N__26409),
            .I(rsmrstn_cascade_));
    InMux I__4875 (
            .O(N__26406),
            .I(N__26403));
    LocalMux I__4874 (
            .O(N__26403),
            .I(N__26400));
    Span4Mux_h I__4873 (
            .O(N__26400),
            .I(N__26397));
    Odrv4 I__4872 (
            .O(N__26397),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_0_2 ));
    CascadeMux I__4871 (
            .O(N__26394),
            .I(N__26391));
    InMux I__4870 (
            .O(N__26391),
            .I(N__26388));
    LocalMux I__4869 (
            .O(N__26388),
            .I(N__26385));
    Span4Mux_v I__4868 (
            .O(N__26385),
            .I(N__26382));
    Span4Mux_v I__4867 (
            .O(N__26382),
            .I(N__26379));
    Sp12to4 I__4866 (
            .O(N__26379),
            .I(N__26376));
    Odrv12 I__4865 (
            .O(N__26376),
            .I(vr_ready_vccin));
    CascadeMux I__4864 (
            .O(N__26373),
            .I(\b2v_inst6.N_192_cascade_ ));
    CascadeMux I__4863 (
            .O(N__26370),
            .I(\b2v_inst6.N_241_cascade_ ));
    CascadeMux I__4862 (
            .O(N__26367),
            .I(\b2v_inst11.count_clk_RNIG8KAHZ0Z_7_cascade_ ));
    CascadeMux I__4861 (
            .O(N__26364),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_ ));
    InMux I__4860 (
            .O(N__26361),
            .I(N__26358));
    LocalMux I__4859 (
            .O(N__26358),
            .I(\b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1 ));
    CascadeMux I__4858 (
            .O(N__26355),
            .I(\b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1_cascade_ ));
    InMux I__4857 (
            .O(N__26352),
            .I(N__26346));
    InMux I__4856 (
            .O(N__26351),
            .I(N__26346));
    LocalMux I__4855 (
            .O(N__26346),
            .I(\b2v_inst5.count_1_10 ));
    CascadeMux I__4854 (
            .O(N__26343),
            .I(\b2v_inst5.count_rst_4_cascade_ ));
    InMux I__4853 (
            .O(N__26340),
            .I(N__26337));
    LocalMux I__4852 (
            .O(N__26337),
            .I(N__26334));
    Span4Mux_v I__4851 (
            .O(N__26334),
            .I(N__26331));
    Odrv4 I__4850 (
            .O(N__26331),
            .I(\b2v_inst5.un12_clk_100khz_4 ));
    InMux I__4849 (
            .O(N__26328),
            .I(N__26325));
    LocalMux I__4848 (
            .O(N__26325),
            .I(\b2v_inst5.un12_clk_100khz_11 ));
    CascadeMux I__4847 (
            .O(N__26322),
            .I(\b2v_inst5.un12_clk_100khz_5_cascade_ ));
    InMux I__4846 (
            .O(N__26319),
            .I(N__26316));
    LocalMux I__4845 (
            .O(N__26316),
            .I(\b2v_inst5.un12_clk_100khz_12 ));
    CascadeMux I__4844 (
            .O(N__26313),
            .I(\b2v_inst5.N_1_i_cascade_ ));
    CEMux I__4843 (
            .O(N__26310),
            .I(N__26307));
    LocalMux I__4842 (
            .O(N__26307),
            .I(N__26303));
    CEMux I__4841 (
            .O(N__26306),
            .I(N__26300));
    Span4Mux_s0_v I__4840 (
            .O(N__26303),
            .I(N__26295));
    LocalMux I__4839 (
            .O(N__26300),
            .I(N__26295));
    Span4Mux_v I__4838 (
            .O(N__26295),
            .I(N__26291));
    CEMux I__4837 (
            .O(N__26294),
            .I(N__26288));
    Span4Mux_h I__4836 (
            .O(N__26291),
            .I(N__26282));
    LocalMux I__4835 (
            .O(N__26288),
            .I(N__26282));
    CEMux I__4834 (
            .O(N__26287),
            .I(N__26279));
    Span4Mux_h I__4833 (
            .O(N__26282),
            .I(N__26271));
    LocalMux I__4832 (
            .O(N__26279),
            .I(N__26271));
    CascadeMux I__4831 (
            .O(N__26278),
            .I(N__26267));
    CascadeMux I__4830 (
            .O(N__26277),
            .I(N__26259));
    CEMux I__4829 (
            .O(N__26276),
            .I(N__26247));
    Span4Mux_v I__4828 (
            .O(N__26271),
            .I(N__26244));
    CEMux I__4827 (
            .O(N__26270),
            .I(N__26233));
    InMux I__4826 (
            .O(N__26267),
            .I(N__26233));
    InMux I__4825 (
            .O(N__26266),
            .I(N__26233));
    InMux I__4824 (
            .O(N__26265),
            .I(N__26233));
    InMux I__4823 (
            .O(N__26264),
            .I(N__26233));
    InMux I__4822 (
            .O(N__26263),
            .I(N__26224));
    InMux I__4821 (
            .O(N__26262),
            .I(N__26224));
    InMux I__4820 (
            .O(N__26259),
            .I(N__26224));
    InMux I__4819 (
            .O(N__26258),
            .I(N__26224));
    InMux I__4818 (
            .O(N__26257),
            .I(N__26216));
    InMux I__4817 (
            .O(N__26256),
            .I(N__26216));
    InMux I__4816 (
            .O(N__26255),
            .I(N__26209));
    InMux I__4815 (
            .O(N__26254),
            .I(N__26209));
    InMux I__4814 (
            .O(N__26253),
            .I(N__26209));
    InMux I__4813 (
            .O(N__26252),
            .I(N__26202));
    InMux I__4812 (
            .O(N__26251),
            .I(N__26202));
    InMux I__4811 (
            .O(N__26250),
            .I(N__26202));
    LocalMux I__4810 (
            .O(N__26247),
            .I(N__26193));
    Span4Mux_s0_v I__4809 (
            .O(N__26244),
            .I(N__26193));
    LocalMux I__4808 (
            .O(N__26233),
            .I(N__26193));
    LocalMux I__4807 (
            .O(N__26224),
            .I(N__26193));
    InMux I__4806 (
            .O(N__26223),
            .I(N__26190));
    InMux I__4805 (
            .O(N__26222),
            .I(N__26185));
    InMux I__4804 (
            .O(N__26221),
            .I(N__26185));
    LocalMux I__4803 (
            .O(N__26216),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__4802 (
            .O(N__26209),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__4801 (
            .O(N__26202),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    Odrv4 I__4800 (
            .O(N__26193),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__4799 (
            .O(N__26190),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    LocalMux I__4798 (
            .O(N__26185),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ));
    CascadeMux I__4797 (
            .O(N__26172),
            .I(N__26169));
    InMux I__4796 (
            .O(N__26169),
            .I(N__26166));
    LocalMux I__4795 (
            .O(N__26166),
            .I(\b2v_inst5.count_1_9 ));
    CascadeMux I__4794 (
            .O(N__26163),
            .I(N__26159));
    InMux I__4793 (
            .O(N__26162),
            .I(N__26156));
    InMux I__4792 (
            .O(N__26159),
            .I(N__26152));
    LocalMux I__4791 (
            .O(N__26156),
            .I(N__26149));
    InMux I__4790 (
            .O(N__26155),
            .I(N__26146));
    LocalMux I__4789 (
            .O(N__26152),
            .I(N__26143));
    Odrv4 I__4788 (
            .O(N__26149),
            .I(\b2v_inst5.countZ0Z_13 ));
    LocalMux I__4787 (
            .O(N__26146),
            .I(\b2v_inst5.countZ0Z_13 ));
    Odrv4 I__4786 (
            .O(N__26143),
            .I(\b2v_inst5.countZ0Z_13 ));
    InMux I__4785 (
            .O(N__26136),
            .I(N__26132));
    InMux I__4784 (
            .O(N__26135),
            .I(N__26129));
    LocalMux I__4783 (
            .O(N__26132),
            .I(N__26126));
    LocalMux I__4782 (
            .O(N__26129),
            .I(N__26123));
    Odrv4 I__4781 (
            .O(N__26126),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    Odrv12 I__4780 (
            .O(N__26123),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    InMux I__4779 (
            .O(N__26118),
            .I(N__26115));
    LocalMux I__4778 (
            .O(N__26115),
            .I(N__26112));
    Odrv4 I__4777 (
            .O(N__26112),
            .I(\b2v_inst5.count_rst_1 ));
    CascadeMux I__4776 (
            .O(N__26109),
            .I(N__26105));
    InMux I__4775 (
            .O(N__26108),
            .I(N__26091));
    InMux I__4774 (
            .O(N__26105),
            .I(N__26091));
    InMux I__4773 (
            .O(N__26104),
            .I(N__26091));
    InMux I__4772 (
            .O(N__26103),
            .I(N__26091));
    InMux I__4771 (
            .O(N__26102),
            .I(N__26091));
    LocalMux I__4770 (
            .O(N__26091),
            .I(N__26082));
    InMux I__4769 (
            .O(N__26090),
            .I(N__26078));
    InMux I__4768 (
            .O(N__26089),
            .I(N__26075));
    InMux I__4767 (
            .O(N__26088),
            .I(N__26070));
    InMux I__4766 (
            .O(N__26087),
            .I(N__26070));
    InMux I__4765 (
            .O(N__26086),
            .I(N__26065));
    InMux I__4764 (
            .O(N__26085),
            .I(N__26065));
    Span4Mux_h I__4763 (
            .O(N__26082),
            .I(N__26062));
    InMux I__4762 (
            .O(N__26081),
            .I(N__26059));
    LocalMux I__4761 (
            .O(N__26078),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__4760 (
            .O(N__26075),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__4759 (
            .O(N__26070),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__4758 (
            .O(N__26065),
            .I(\b2v_inst5.N_1_i ));
    Odrv4 I__4757 (
            .O(N__26062),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__4756 (
            .O(N__26059),
            .I(\b2v_inst5.N_1_i ));
    InMux I__4755 (
            .O(N__26046),
            .I(N__26042));
    InMux I__4754 (
            .O(N__26045),
            .I(N__26039));
    LocalMux I__4753 (
            .O(N__26042),
            .I(N__26036));
    LocalMux I__4752 (
            .O(N__26039),
            .I(N__26031));
    Span4Mux_s3_v I__4751 (
            .O(N__26036),
            .I(N__26031));
    Odrv4 I__4750 (
            .O(N__26031),
            .I(\b2v_inst5.un2_count_1_cry_8_THRU_CO ));
    InMux I__4749 (
            .O(N__26028),
            .I(N__26024));
    CascadeMux I__4748 (
            .O(N__26027),
            .I(N__26021));
    LocalMux I__4747 (
            .O(N__26024),
            .I(N__26018));
    InMux I__4746 (
            .O(N__26021),
            .I(N__26013));
    Span4Mux_h I__4745 (
            .O(N__26018),
            .I(N__26010));
    InMux I__4744 (
            .O(N__26017),
            .I(N__26005));
    InMux I__4743 (
            .O(N__26016),
            .I(N__26005));
    LocalMux I__4742 (
            .O(N__26013),
            .I(\b2v_inst5.countZ0Z_9 ));
    Odrv4 I__4741 (
            .O(N__26010),
            .I(\b2v_inst5.countZ0Z_9 ));
    LocalMux I__4740 (
            .O(N__26005),
            .I(\b2v_inst5.countZ0Z_9 ));
    SRMux I__4739 (
            .O(N__25998),
            .I(N__25995));
    LocalMux I__4738 (
            .O(N__25995),
            .I(N__25992));
    Span4Mux_v I__4737 (
            .O(N__25992),
            .I(N__25985));
    SRMux I__4736 (
            .O(N__25991),
            .I(N__25982));
    SRMux I__4735 (
            .O(N__25990),
            .I(N__25971));
    CascadeMux I__4734 (
            .O(N__25989),
            .I(N__25967));
    SRMux I__4733 (
            .O(N__25988),
            .I(N__25955));
    Span4Mux_h I__4732 (
            .O(N__25985),
            .I(N__25950));
    LocalMux I__4731 (
            .O(N__25982),
            .I(N__25950));
    InMux I__4730 (
            .O(N__25981),
            .I(N__25947));
    SRMux I__4729 (
            .O(N__25980),
            .I(N__25944));
    InMux I__4728 (
            .O(N__25979),
            .I(N__25937));
    InMux I__4727 (
            .O(N__25978),
            .I(N__25937));
    SRMux I__4726 (
            .O(N__25977),
            .I(N__25937));
    InMux I__4725 (
            .O(N__25976),
            .I(N__25934));
    InMux I__4724 (
            .O(N__25975),
            .I(N__25929));
    InMux I__4723 (
            .O(N__25974),
            .I(N__25929));
    LocalMux I__4722 (
            .O(N__25971),
            .I(N__25926));
    InMux I__4721 (
            .O(N__25970),
            .I(N__25915));
    InMux I__4720 (
            .O(N__25967),
            .I(N__25915));
    InMux I__4719 (
            .O(N__25966),
            .I(N__25915));
    InMux I__4718 (
            .O(N__25965),
            .I(N__25915));
    InMux I__4717 (
            .O(N__25964),
            .I(N__25915));
    InMux I__4716 (
            .O(N__25963),
            .I(N__25904));
    InMux I__4715 (
            .O(N__25962),
            .I(N__25904));
    InMux I__4714 (
            .O(N__25961),
            .I(N__25904));
    InMux I__4713 (
            .O(N__25960),
            .I(N__25904));
    InMux I__4712 (
            .O(N__25959),
            .I(N__25904));
    CascadeMux I__4711 (
            .O(N__25958),
            .I(N__25899));
    LocalMux I__4710 (
            .O(N__25955),
            .I(N__25893));
    Span4Mux_h I__4709 (
            .O(N__25950),
            .I(N__25884));
    LocalMux I__4708 (
            .O(N__25947),
            .I(N__25884));
    LocalMux I__4707 (
            .O(N__25944),
            .I(N__25884));
    LocalMux I__4706 (
            .O(N__25937),
            .I(N__25884));
    LocalMux I__4705 (
            .O(N__25934),
            .I(N__25879));
    LocalMux I__4704 (
            .O(N__25929),
            .I(N__25876));
    Span4Mux_s1_v I__4703 (
            .O(N__25926),
            .I(N__25869));
    LocalMux I__4702 (
            .O(N__25915),
            .I(N__25869));
    LocalMux I__4701 (
            .O(N__25904),
            .I(N__25869));
    InMux I__4700 (
            .O(N__25903),
            .I(N__25858));
    InMux I__4699 (
            .O(N__25902),
            .I(N__25858));
    InMux I__4698 (
            .O(N__25899),
            .I(N__25858));
    InMux I__4697 (
            .O(N__25898),
            .I(N__25858));
    InMux I__4696 (
            .O(N__25897),
            .I(N__25858));
    CascadeMux I__4695 (
            .O(N__25896),
            .I(N__25850));
    Span4Mux_s1_v I__4694 (
            .O(N__25893),
            .I(N__25846));
    Span4Mux_v I__4693 (
            .O(N__25884),
            .I(N__25843));
    InMux I__4692 (
            .O(N__25883),
            .I(N__25840));
    InMux I__4691 (
            .O(N__25882),
            .I(N__25837));
    Span4Mux_s2_v I__4690 (
            .O(N__25879),
            .I(N__25832));
    Span4Mux_h I__4689 (
            .O(N__25876),
            .I(N__25832));
    Span4Mux_h I__4688 (
            .O(N__25869),
            .I(N__25827));
    LocalMux I__4687 (
            .O(N__25858),
            .I(N__25827));
    InMux I__4686 (
            .O(N__25857),
            .I(N__25816));
    InMux I__4685 (
            .O(N__25856),
            .I(N__25816));
    InMux I__4684 (
            .O(N__25855),
            .I(N__25816));
    InMux I__4683 (
            .O(N__25854),
            .I(N__25816));
    InMux I__4682 (
            .O(N__25853),
            .I(N__25816));
    InMux I__4681 (
            .O(N__25850),
            .I(N__25811));
    InMux I__4680 (
            .O(N__25849),
            .I(N__25811));
    Odrv4 I__4679 (
            .O(N__25846),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__4678 (
            .O(N__25843),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__4677 (
            .O(N__25840),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__4676 (
            .O(N__25837),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__4675 (
            .O(N__25832),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__4674 (
            .O(N__25827),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__4673 (
            .O(N__25816),
            .I(\b2v_inst5.count_0_sqmuxa ));
    LocalMux I__4672 (
            .O(N__25811),
            .I(\b2v_inst5.count_0_sqmuxa ));
    InMux I__4671 (
            .O(N__25794),
            .I(N__25791));
    LocalMux I__4670 (
            .O(N__25791),
            .I(\b2v_inst5.count_rst_5 ));
    InMux I__4669 (
            .O(N__25788),
            .I(N__25785));
    LocalMux I__4668 (
            .O(N__25785),
            .I(N__25782));
    Sp12to4 I__4667 (
            .O(N__25782),
            .I(N__25779));
    Span12Mux_v I__4666 (
            .O(N__25779),
            .I(N__25776));
    Odrv12 I__4665 (
            .O(N__25776),
            .I(v33a_ok));
    InMux I__4664 (
            .O(N__25773),
            .I(N__25770));
    LocalMux I__4663 (
            .O(N__25770),
            .I(N__25767));
    Span4Mux_v I__4662 (
            .O(N__25767),
            .I(N__25764));
    Odrv4 I__4661 (
            .O(N__25764),
            .I(vccst_cpu_ok));
    CascadeMux I__4660 (
            .O(N__25761),
            .I(N__25758));
    InMux I__4659 (
            .O(N__25758),
            .I(N__25755));
    LocalMux I__4658 (
            .O(N__25755),
            .I(N__25752));
    Span4Mux_h I__4657 (
            .O(N__25752),
            .I(N__25749));
    Sp12to4 I__4656 (
            .O(N__25749),
            .I(N__25746));
    Span12Mux_s11_v I__4655 (
            .O(N__25746),
            .I(N__25743));
    Odrv12 I__4654 (
            .O(N__25743),
            .I(v1p8a_ok));
    InMux I__4653 (
            .O(N__25740),
            .I(N__25737));
    LocalMux I__4652 (
            .O(N__25737),
            .I(N__25734));
    Span12Mux_s4_v I__4651 (
            .O(N__25734),
            .I(N__25731));
    Odrv12 I__4650 (
            .O(N__25731),
            .I(v5a_ok));
    InMux I__4649 (
            .O(N__25728),
            .I(N__25725));
    LocalMux I__4648 (
            .O(N__25725),
            .I(N__25722));
    Span4Mux_v I__4647 (
            .O(N__25722),
            .I(N__25719));
    Span4Mux_h I__4646 (
            .O(N__25719),
            .I(N__25716));
    Odrv4 I__4645 (
            .O(N__25716),
            .I(vr_ready_vccinaux));
    InMux I__4644 (
            .O(N__25713),
            .I(N__25704));
    InMux I__4643 (
            .O(N__25712),
            .I(N__25704));
    InMux I__4642 (
            .O(N__25711),
            .I(N__25704));
    LocalMux I__4641 (
            .O(N__25704),
            .I(N__25701));
    Span4Mux_s3_v I__4640 (
            .O(N__25701),
            .I(N__25698));
    Odrv4 I__4639 (
            .O(N__25698),
            .I(\b2v_inst5.count_rst_3 ));
    InMux I__4638 (
            .O(N__25695),
            .I(N__25691));
    InMux I__4637 (
            .O(N__25694),
            .I(N__25688));
    LocalMux I__4636 (
            .O(N__25691),
            .I(\b2v_inst5.count_1_11 ));
    LocalMux I__4635 (
            .O(N__25688),
            .I(\b2v_inst5.count_1_11 ));
    CascadeMux I__4634 (
            .O(N__25683),
            .I(\b2v_inst5.countZ0Z_7_cascade_ ));
    InMux I__4633 (
            .O(N__25680),
            .I(N__25674));
    InMux I__4632 (
            .O(N__25679),
            .I(N__25674));
    LocalMux I__4631 (
            .O(N__25674),
            .I(N__25671));
    Span4Mux_s2_v I__4630 (
            .O(N__25671),
            .I(N__25668));
    Odrv4 I__4629 (
            .O(N__25668),
            .I(\b2v_inst5.un2_count_1_cry_1_c_RNIMEQZ0Z9 ));
    CascadeMux I__4628 (
            .O(N__25665),
            .I(N__25662));
    InMux I__4627 (
            .O(N__25662),
            .I(N__25659));
    LocalMux I__4626 (
            .O(N__25659),
            .I(\b2v_inst5.count_1_2 ));
    InMux I__4625 (
            .O(N__25656),
            .I(N__25652));
    InMux I__4624 (
            .O(N__25655),
            .I(N__25649));
    LocalMux I__4623 (
            .O(N__25652),
            .I(N__25646));
    LocalMux I__4622 (
            .O(N__25649),
            .I(N__25643));
    Span4Mux_h I__4621 (
            .O(N__25646),
            .I(N__25640));
    Odrv4 I__4620 (
            .O(N__25643),
            .I(\b2v_inst5.countZ0Z_2 ));
    Odrv4 I__4619 (
            .O(N__25640),
            .I(\b2v_inst5.countZ0Z_2 ));
    InMux I__4618 (
            .O(N__25635),
            .I(N__25632));
    LocalMux I__4617 (
            .O(N__25632),
            .I(N__25628));
    InMux I__4616 (
            .O(N__25631),
            .I(N__25625));
    Span4Mux_h I__4615 (
            .O(N__25628),
            .I(N__25622));
    LocalMux I__4614 (
            .O(N__25625),
            .I(N__25619));
    Odrv4 I__4613 (
            .O(N__25622),
            .I(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ));
    Odrv4 I__4612 (
            .O(N__25619),
            .I(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ));
    CascadeMux I__4611 (
            .O(N__25614),
            .I(N__25611));
    InMux I__4610 (
            .O(N__25611),
            .I(N__25608));
    LocalMux I__4609 (
            .O(N__25608),
            .I(\b2v_inst5.count_1_3 ));
    CascadeMux I__4608 (
            .O(N__25605),
            .I(\b2v_inst5.un2_count_1_axb_10_cascade_ ));
    InMux I__4607 (
            .O(N__25602),
            .I(N__25599));
    LocalMux I__4606 (
            .O(N__25599),
            .I(\b2v_inst5.un12_clk_100khz_9 ));
    InMux I__4605 (
            .O(N__25596),
            .I(N__25592));
    InMux I__4604 (
            .O(N__25595),
            .I(N__25589));
    LocalMux I__4603 (
            .O(N__25592),
            .I(\b2v_inst5.countZ0Z_5 ));
    LocalMux I__4602 (
            .O(N__25589),
            .I(\b2v_inst5.countZ0Z_5 ));
    CascadeMux I__4601 (
            .O(N__25584),
            .I(N__25581));
    InMux I__4600 (
            .O(N__25581),
            .I(N__25578));
    LocalMux I__4599 (
            .O(N__25578),
            .I(\b2v_inst5.un12_clk_100khz_1 ));
    InMux I__4598 (
            .O(N__25575),
            .I(N__25572));
    LocalMux I__4597 (
            .O(N__25572),
            .I(N__25568));
    InMux I__4596 (
            .O(N__25571),
            .I(N__25565));
    Odrv4 I__4595 (
            .O(N__25568),
            .I(\b2v_inst5.countZ0Z_6 ));
    LocalMux I__4594 (
            .O(N__25565),
            .I(\b2v_inst5.countZ0Z_6 ));
    InMux I__4593 (
            .O(N__25560),
            .I(N__25557));
    LocalMux I__4592 (
            .O(N__25557),
            .I(N__25553));
    InMux I__4591 (
            .O(N__25556),
            .I(N__25550));
    Span4Mux_h I__4590 (
            .O(N__25553),
            .I(N__25547));
    LocalMux I__4589 (
            .O(N__25550),
            .I(\b2v_inst5.un2_count_1_axb_10 ));
    Odrv4 I__4588 (
            .O(N__25547),
            .I(\b2v_inst5.un2_count_1_axb_10 ));
    CascadeMux I__4587 (
            .O(N__25542),
            .I(N__25538));
    InMux I__4586 (
            .O(N__25541),
            .I(N__25533));
    InMux I__4585 (
            .O(N__25538),
            .I(N__25533));
    LocalMux I__4584 (
            .O(N__25533),
            .I(N__25530));
    Span4Mux_h I__4583 (
            .O(N__25530),
            .I(N__25527));
    Odrv4 I__4582 (
            .O(N__25527),
            .I(\b2v_inst5.un2_count_1_cry_9_THRU_CO ));
    InMux I__4581 (
            .O(N__25524),
            .I(N__25521));
    LocalMux I__4580 (
            .O(N__25521),
            .I(\b2v_inst5.count_rst_4 ));
    CascadeMux I__4579 (
            .O(N__25518),
            .I(\b2v_inst6.count_rst_10_cascade_ ));
    InMux I__4578 (
            .O(N__25515),
            .I(N__25512));
    LocalMux I__4577 (
            .O(N__25512),
            .I(\b2v_inst6.count_rst_11 ));
    InMux I__4576 (
            .O(N__25509),
            .I(N__25503));
    InMux I__4575 (
            .O(N__25508),
            .I(N__25503));
    LocalMux I__4574 (
            .O(N__25503),
            .I(\b2v_inst6.count_0_3 ));
    InMux I__4573 (
            .O(N__25500),
            .I(N__25497));
    LocalMux I__4572 (
            .O(N__25497),
            .I(\b2v_inst6.count_rst_10 ));
    CascadeMux I__4571 (
            .O(N__25494),
            .I(\b2v_inst6.countZ0Z_3_cascade_ ));
    InMux I__4570 (
            .O(N__25491),
            .I(N__25485));
    InMux I__4569 (
            .O(N__25490),
            .I(N__25485));
    LocalMux I__4568 (
            .O(N__25485),
            .I(\b2v_inst6.count_0_4 ));
    InMux I__4567 (
            .O(N__25482),
            .I(N__25479));
    LocalMux I__4566 (
            .O(N__25479),
            .I(N__25476));
    Span4Mux_v I__4565 (
            .O(N__25476),
            .I(N__25473));
    Odrv4 I__4564 (
            .O(N__25473),
            .I(\b2v_inst5.un2_count_1_axb_11 ));
    InMux I__4563 (
            .O(N__25470),
            .I(N__25467));
    LocalMux I__4562 (
            .O(N__25467),
            .I(\b2v_inst5.count_1_7 ));
    InMux I__4561 (
            .O(N__25464),
            .I(N__25458));
    InMux I__4560 (
            .O(N__25463),
            .I(N__25458));
    LocalMux I__4559 (
            .O(N__25458),
            .I(N__25455));
    Span4Mux_s2_v I__4558 (
            .O(N__25455),
            .I(N__25452));
    Odrv4 I__4557 (
            .O(N__25452),
            .I(\b2v_inst5.un2_count_1_cry_6_c_RNIROVZ0Z9 ));
    InMux I__4556 (
            .O(N__25449),
            .I(N__25446));
    LocalMux I__4555 (
            .O(N__25446),
            .I(N__25443));
    Span4Mux_h I__4554 (
            .O(N__25443),
            .I(N__25440));
    Odrv4 I__4553 (
            .O(N__25440),
            .I(\b2v_inst5.countZ0Z_7 ));
    CascadeMux I__4552 (
            .O(N__25437),
            .I(N__25434));
    InMux I__4551 (
            .O(N__25434),
            .I(N__25431));
    LocalMux I__4550 (
            .O(N__25431),
            .I(\b2v_inst11.mult1_un68_sum_cry_4_s ));
    InMux I__4549 (
            .O(N__25428),
            .I(\b2v_inst11.mult1_un68_sum_cry_3 ));
    CascadeMux I__4548 (
            .O(N__25425),
            .I(N__25422));
    InMux I__4547 (
            .O(N__25422),
            .I(N__25419));
    LocalMux I__4546 (
            .O(N__25419),
            .I(\b2v_inst11.mult1_un61_sum_cry_4_s ));
    InMux I__4545 (
            .O(N__25416),
            .I(N__25413));
    LocalMux I__4544 (
            .O(N__25413),
            .I(\b2v_inst11.mult1_un68_sum_cry_5_s ));
    InMux I__4543 (
            .O(N__25410),
            .I(\b2v_inst11.mult1_un68_sum_cry_4 ));
    InMux I__4542 (
            .O(N__25407),
            .I(N__25404));
    LocalMux I__4541 (
            .O(N__25404),
            .I(\b2v_inst11.mult1_un61_sum_cry_5_s ));
    InMux I__4540 (
            .O(N__25401),
            .I(N__25398));
    LocalMux I__4539 (
            .O(N__25398),
            .I(\b2v_inst11.mult1_un68_sum_cry_6_s ));
    InMux I__4538 (
            .O(N__25395),
            .I(\b2v_inst11.mult1_un68_sum_cry_5 ));
    InMux I__4537 (
            .O(N__25392),
            .I(N__25389));
    LocalMux I__4536 (
            .O(N__25389),
            .I(\b2v_inst11.mult1_un61_sum_cry_6_s ));
    CascadeMux I__4535 (
            .O(N__25386),
            .I(N__25383));
    InMux I__4534 (
            .O(N__25383),
            .I(N__25380));
    LocalMux I__4533 (
            .O(N__25380),
            .I(\b2v_inst11.mult1_un75_sum_axb_8 ));
    InMux I__4532 (
            .O(N__25377),
            .I(\b2v_inst11.mult1_un68_sum_cry_6 ));
    CascadeMux I__4531 (
            .O(N__25374),
            .I(N__25371));
    InMux I__4530 (
            .O(N__25371),
            .I(N__25368));
    LocalMux I__4529 (
            .O(N__25368),
            .I(\b2v_inst11.mult1_un68_sum_axb_8 ));
    InMux I__4528 (
            .O(N__25365),
            .I(\b2v_inst11.mult1_un68_sum_cry_7 ));
    InMux I__4527 (
            .O(N__25362),
            .I(N__25359));
    LocalMux I__4526 (
            .O(N__25359),
            .I(N__25356));
    Span4Mux_s2_h I__4525 (
            .O(N__25356),
            .I(N__25352));
    CascadeMux I__4524 (
            .O(N__25355),
            .I(N__25348));
    Span4Mux_h I__4523 (
            .O(N__25352),
            .I(N__25343));
    InMux I__4522 (
            .O(N__25351),
            .I(N__25340));
    InMux I__4521 (
            .O(N__25348),
            .I(N__25333));
    InMux I__4520 (
            .O(N__25347),
            .I(N__25333));
    InMux I__4519 (
            .O(N__25346),
            .I(N__25333));
    Odrv4 I__4518 (
            .O(N__25343),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__4517 (
            .O(N__25340),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__4516 (
            .O(N__25333),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    InMux I__4515 (
            .O(N__25326),
            .I(N__25322));
    CascadeMux I__4514 (
            .O(N__25325),
            .I(N__25318));
    LocalMux I__4513 (
            .O(N__25322),
            .I(N__25313));
    InMux I__4512 (
            .O(N__25321),
            .I(N__25310));
    InMux I__4511 (
            .O(N__25318),
            .I(N__25303));
    InMux I__4510 (
            .O(N__25317),
            .I(N__25303));
    InMux I__4509 (
            .O(N__25316),
            .I(N__25303));
    Odrv12 I__4508 (
            .O(N__25313),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__4507 (
            .O(N__25310),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__4506 (
            .O(N__25303),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    CascadeMux I__4505 (
            .O(N__25296),
            .I(N__25292));
    CascadeMux I__4504 (
            .O(N__25295),
            .I(N__25288));
    InMux I__4503 (
            .O(N__25292),
            .I(N__25281));
    InMux I__4502 (
            .O(N__25291),
            .I(N__25281));
    InMux I__4501 (
            .O(N__25288),
            .I(N__25281));
    LocalMux I__4500 (
            .O(N__25281),
            .I(\b2v_inst11.mult1_un61_sum_i_0_8 ));
    CascadeMux I__4499 (
            .O(N__25278),
            .I(\b2v_inst6.count_rst_11_cascade_ ));
    CascadeMux I__4498 (
            .O(N__25275),
            .I(\b2v_inst6.un2_count_1_axb_3_cascade_ ));
    InMux I__4497 (
            .O(N__25272),
            .I(N__25269));
    LocalMux I__4496 (
            .O(N__25269),
            .I(\b2v_inst11.mult1_un54_sum_cry_3_s ));
    CascadeMux I__4495 (
            .O(N__25266),
            .I(N__25263));
    InMux I__4494 (
            .O(N__25263),
            .I(N__25256));
    InMux I__4493 (
            .O(N__25262),
            .I(N__25256));
    InMux I__4492 (
            .O(N__25261),
            .I(N__25253));
    LocalMux I__4491 (
            .O(N__25256),
            .I(\b2v_inst11.mult1_un54_sum_cry_7_THRU_CO ));
    LocalMux I__4490 (
            .O(N__25253),
            .I(\b2v_inst11.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__4489 (
            .O(N__25248),
            .I(\b2v_inst11.mult1_un61_sum_cry_3 ));
    CascadeMux I__4488 (
            .O(N__25245),
            .I(N__25242));
    InMux I__4487 (
            .O(N__25242),
            .I(N__25239));
    LocalMux I__4486 (
            .O(N__25239),
            .I(\b2v_inst11.mult1_un54_sum_cry_4_s ));
    InMux I__4485 (
            .O(N__25236),
            .I(\b2v_inst11.mult1_un61_sum_cry_4 ));
    InMux I__4484 (
            .O(N__25233),
            .I(N__25230));
    LocalMux I__4483 (
            .O(N__25230),
            .I(\b2v_inst11.mult1_un54_sum_cry_5_s ));
    InMux I__4482 (
            .O(N__25227),
            .I(\b2v_inst11.mult1_un61_sum_cry_5 ));
    InMux I__4481 (
            .O(N__25224),
            .I(N__25221));
    LocalMux I__4480 (
            .O(N__25221),
            .I(\b2v_inst11.mult1_un54_sum_cry_6_s ));
    InMux I__4479 (
            .O(N__25218),
            .I(\b2v_inst11.mult1_un61_sum_cry_6 ));
    InMux I__4478 (
            .O(N__25215),
            .I(N__25212));
    LocalMux I__4477 (
            .O(N__25212),
            .I(\b2v_inst11.mult1_un54_sum_cry_6_THRU_CO ));
    InMux I__4476 (
            .O(N__25209),
            .I(\b2v_inst11.mult1_un61_sum_cry_7 ));
    CascadeMux I__4475 (
            .O(N__25206),
            .I(N__25202));
    CascadeMux I__4474 (
            .O(N__25205),
            .I(N__25199));
    InMux I__4473 (
            .O(N__25202),
            .I(N__25188));
    InMux I__4472 (
            .O(N__25199),
            .I(N__25188));
    InMux I__4471 (
            .O(N__25198),
            .I(N__25188));
    InMux I__4470 (
            .O(N__25197),
            .I(N__25188));
    LocalMux I__4469 (
            .O(N__25188),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    CascadeMux I__4468 (
            .O(N__25185),
            .I(N__25182));
    InMux I__4467 (
            .O(N__25182),
            .I(N__25179));
    LocalMux I__4466 (
            .O(N__25179),
            .I(\b2v_inst11.mult1_un54_sum_i_8 ));
    CascadeMux I__4465 (
            .O(N__25176),
            .I(N__25173));
    InMux I__4464 (
            .O(N__25173),
            .I(N__25170));
    LocalMux I__4463 (
            .O(N__25170),
            .I(\b2v_inst11.mult1_un68_sum_cry_3_s ));
    InMux I__4462 (
            .O(N__25167),
            .I(\b2v_inst11.mult1_un68_sum_cry_2 ));
    CascadeMux I__4461 (
            .O(N__25164),
            .I(N__25161));
    InMux I__4460 (
            .O(N__25161),
            .I(N__25158));
    LocalMux I__4459 (
            .O(N__25158),
            .I(\b2v_inst11.mult1_un61_sum_cry_3_s ));
    CascadeMux I__4458 (
            .O(N__25155),
            .I(N__25152));
    InMux I__4457 (
            .O(N__25152),
            .I(N__25149));
    LocalMux I__4456 (
            .O(N__25149),
            .I(\b2v_inst11.mult1_un54_sum_s_3_sf ));
    InMux I__4455 (
            .O(N__25146),
            .I(\b2v_inst11.mult1_un54_sum_cry_2 ));
    InMux I__4454 (
            .O(N__25143),
            .I(\b2v_inst11.mult1_un54_sum_cry_3 ));
    InMux I__4453 (
            .O(N__25140),
            .I(\b2v_inst11.mult1_un54_sum_cry_4 ));
    InMux I__4452 (
            .O(N__25137),
            .I(\b2v_inst11.mult1_un54_sum_cry_5 ));
    InMux I__4451 (
            .O(N__25134),
            .I(\b2v_inst11.mult1_un54_sum_cry_6 ));
    InMux I__4450 (
            .O(N__25131),
            .I(\b2v_inst11.mult1_un54_sum_cry_7 ));
    CascadeMux I__4449 (
            .O(N__25128),
            .I(N__25125));
    InMux I__4448 (
            .O(N__25125),
            .I(N__25122));
    LocalMux I__4447 (
            .O(N__25122),
            .I(N__25119));
    Odrv4 I__4446 (
            .O(N__25119),
            .I(\b2v_inst11.mult1_un47_sum_i_1 ));
    InMux I__4445 (
            .O(N__25116),
            .I(\b2v_inst11.mult1_un61_sum_cry_2 ));
    InMux I__4444 (
            .O(N__25113),
            .I(N__25110));
    LocalMux I__4443 (
            .O(N__25110),
            .I(\b2v_inst11.g0_3_2_0 ));
    CascadeMux I__4442 (
            .O(N__25107),
            .I(\b2v_inst11.un2_count_clk_17_0_a2_1_4_cascade_ ));
    CascadeMux I__4441 (
            .O(N__25104),
            .I(\b2v_inst11.N_363_cascade_ ));
    InMux I__4440 (
            .O(N__25101),
            .I(N__25098));
    LocalMux I__4439 (
            .O(N__25098),
            .I(N__25095));
    Odrv4 I__4438 (
            .O(N__25095),
            .I(\b2v_inst11.mult1_un145_sum_i ));
    InMux I__4437 (
            .O(N__25092),
            .I(N__25089));
    LocalMux I__4436 (
            .O(N__25089),
            .I(N__25086));
    Odrv12 I__4435 (
            .O(N__25086),
            .I(\b2v_inst11.mult1_un131_sum_i ));
    CascadeMux I__4434 (
            .O(N__25083),
            .I(\b2v_inst11.N_3055_0_cascade_ ));
    InMux I__4433 (
            .O(N__25080),
            .I(N__25077));
    LocalMux I__4432 (
            .O(N__25077),
            .I(\b2v_inst11.dutycycle_RNI_14Z0Z_0 ));
    CascadeMux I__4431 (
            .O(N__25074),
            .I(\b2v_inst11.un1_dutycycle_172_m3_0_cascade_ ));
    InMux I__4430 (
            .O(N__25071),
            .I(N__25068));
    LocalMux I__4429 (
            .O(N__25068),
            .I(\b2v_inst11.un1_dutycycle_172_0 ));
    CascadeMux I__4428 (
            .O(N__25065),
            .I(\b2v_inst11.N_19_i_cascade_ ));
    CascadeMux I__4427 (
            .O(N__25062),
            .I(\b2v_inst11.un1_dutycycle_172_m0_ns_1_cascade_ ));
    InMux I__4426 (
            .O(N__25059),
            .I(N__25056));
    LocalMux I__4425 (
            .O(N__25056),
            .I(\b2v_inst11.un1_dutycycle_172_m0 ));
    CascadeMux I__4424 (
            .O(N__25053),
            .I(\b2v_inst11.g0_4_1_cascade_ ));
    InMux I__4423 (
            .O(N__25050),
            .I(N__25047));
    LocalMux I__4422 (
            .O(N__25047),
            .I(\b2v_inst11.N_293_0 ));
    CascadeMux I__4421 (
            .O(N__25044),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVKZ0_cascade_ ));
    InMux I__4420 (
            .O(N__25041),
            .I(N__25038));
    LocalMux I__4419 (
            .O(N__25038),
            .I(\b2v_inst11.N_236 ));
    CascadeMux I__4418 (
            .O(N__25035),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ));
    InMux I__4417 (
            .O(N__25032),
            .I(N__25029));
    LocalMux I__4416 (
            .O(N__25029),
            .I(\b2v_inst11.N_295 ));
    InMux I__4415 (
            .O(N__25026),
            .I(N__25023));
    LocalMux I__4414 (
            .O(N__25023),
            .I(\b2v_inst11.mult1_un152_sum_i ));
    CascadeMux I__4413 (
            .O(N__25020),
            .I(v5s_enn_cascade_));
    InMux I__4412 (
            .O(N__25017),
            .I(N__25014));
    LocalMux I__4411 (
            .O(N__25014),
            .I(N__25009));
    InMux I__4410 (
            .O(N__25013),
            .I(N__25006));
    CascadeMux I__4409 (
            .O(N__25012),
            .I(N__25003));
    Span4Mux_v I__4408 (
            .O(N__25009),
            .I(N__24999));
    LocalMux I__4407 (
            .O(N__25006),
            .I(N__24996));
    InMux I__4406 (
            .O(N__25003),
            .I(N__24991));
    InMux I__4405 (
            .O(N__25002),
            .I(N__24991));
    Odrv4 I__4404 (
            .O(N__24999),
            .I(\b2v_inst20.counterZ0Z_0 ));
    Odrv4 I__4403 (
            .O(N__24996),
            .I(\b2v_inst20.counterZ0Z_0 ));
    LocalMux I__4402 (
            .O(N__24991),
            .I(\b2v_inst20.counterZ0Z_0 ));
    InMux I__4401 (
            .O(N__24984),
            .I(N__24981));
    LocalMux I__4400 (
            .O(N__24981),
            .I(\b2v_inst20.un4_counter_0_and ));
    InMux I__4399 (
            .O(N__24978),
            .I(N__24975));
    LocalMux I__4398 (
            .O(N__24975),
            .I(N__24972));
    Odrv12 I__4397 (
            .O(N__24972),
            .I(\b2v_inst20.counter_1_cry_1_THRU_CO ));
    InMux I__4396 (
            .O(N__24969),
            .I(N__24965));
    CascadeMux I__4395 (
            .O(N__24968),
            .I(N__24962));
    LocalMux I__4394 (
            .O(N__24965),
            .I(N__24958));
    InMux I__4393 (
            .O(N__24962),
            .I(N__24953));
    InMux I__4392 (
            .O(N__24961),
            .I(N__24953));
    Odrv4 I__4391 (
            .O(N__24958),
            .I(\b2v_inst20.counterZ0Z_2 ));
    LocalMux I__4390 (
            .O(N__24953),
            .I(\b2v_inst20.counterZ0Z_2 ));
    InMux I__4389 (
            .O(N__24948),
            .I(N__24945));
    LocalMux I__4388 (
            .O(N__24945),
            .I(N__24942));
    Odrv12 I__4387 (
            .O(N__24942),
            .I(\b2v_inst20.counter_1_cry_2_THRU_CO ));
    InMux I__4386 (
            .O(N__24939),
            .I(N__24935));
    CascadeMux I__4385 (
            .O(N__24938),
            .I(N__24931));
    LocalMux I__4384 (
            .O(N__24935),
            .I(N__24928));
    InMux I__4383 (
            .O(N__24934),
            .I(N__24923));
    InMux I__4382 (
            .O(N__24931),
            .I(N__24923));
    Odrv12 I__4381 (
            .O(N__24928),
            .I(\b2v_inst20.counterZ0Z_3 ));
    LocalMux I__4380 (
            .O(N__24923),
            .I(\b2v_inst20.counterZ0Z_3 ));
    InMux I__4379 (
            .O(N__24918),
            .I(N__24915));
    LocalMux I__4378 (
            .O(N__24915),
            .I(N__24912));
    Odrv12 I__4377 (
            .O(N__24912),
            .I(\b2v_inst20.counter_1_cry_3_THRU_CO ));
    InMux I__4376 (
            .O(N__24909),
            .I(N__24906));
    LocalMux I__4375 (
            .O(N__24906),
            .I(N__24901));
    InMux I__4374 (
            .O(N__24905),
            .I(N__24896));
    InMux I__4373 (
            .O(N__24904),
            .I(N__24896));
    Odrv4 I__4372 (
            .O(N__24901),
            .I(\b2v_inst20.counterZ0Z_4 ));
    LocalMux I__4371 (
            .O(N__24896),
            .I(\b2v_inst20.counterZ0Z_4 ));
    CascadeMux I__4370 (
            .O(N__24891),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_1_cascade_ ));
    CascadeMux I__4369 (
            .O(N__24888),
            .I(N__24885));
    InMux I__4368 (
            .O(N__24885),
            .I(N__24882));
    LocalMux I__4367 (
            .O(N__24882),
            .I(\b2v_inst11.func_state_1_m2_1 ));
    InMux I__4366 (
            .O(N__24879),
            .I(N__24873));
    InMux I__4365 (
            .O(N__24878),
            .I(N__24873));
    LocalMux I__4364 (
            .O(N__24873),
            .I(\b2v_inst11.func_stateZ0Z_1 ));
    CascadeMux I__4363 (
            .O(N__24870),
            .I(\b2v_inst11.un1_clk_100khz_51_and_i_a3_0_1_cascade_ ));
    InMux I__4362 (
            .O(N__24867),
            .I(N__24864));
    LocalMux I__4361 (
            .O(N__24864),
            .I(N__24861));
    Span4Mux_v I__4360 (
            .O(N__24861),
            .I(N__24858));
    Span4Mux_v I__4359 (
            .O(N__24858),
            .I(N__24855));
    Span4Mux_h I__4358 (
            .O(N__24855),
            .I(N__24852));
    Odrv4 I__4357 (
            .O(N__24852),
            .I(vpp_ok));
    CascadeMux I__4356 (
            .O(N__24849),
            .I(VCCST_EN_i_0_o3_0_cascade_));
    IoInMux I__4355 (
            .O(N__24846),
            .I(N__24843));
    LocalMux I__4354 (
            .O(N__24843),
            .I(N__24840));
    IoSpan4Mux I__4353 (
            .O(N__24840),
            .I(N__24837));
    Span4Mux_s2_h I__4352 (
            .O(N__24837),
            .I(N__24834));
    Span4Mux_h I__4351 (
            .O(N__24834),
            .I(N__24831));
    Span4Mux_v I__4350 (
            .O(N__24831),
            .I(N__24828));
    Odrv4 I__4349 (
            .O(N__24828),
            .I(vddq_en));
    CascadeMux I__4348 (
            .O(N__24825),
            .I(\b2v_inst11.count_clk_en_0_xZ0Z1_cascade_ ));
    InMux I__4347 (
            .O(N__24822),
            .I(N__24819));
    LocalMux I__4346 (
            .O(N__24819),
            .I(N__24816));
    Odrv4 I__4345 (
            .O(N__24816),
            .I(\b2v_inst11.N_335 ));
    InMux I__4344 (
            .O(N__24813),
            .I(N__24810));
    LocalMux I__4343 (
            .O(N__24810),
            .I(N__24807));
    Span4Mux_v I__4342 (
            .O(N__24807),
            .I(N__24803));
    InMux I__4341 (
            .O(N__24806),
            .I(N__24800));
    Odrv4 I__4340 (
            .O(N__24803),
            .I(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ));
    LocalMux I__4339 (
            .O(N__24800),
            .I(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ));
    InMux I__4338 (
            .O(N__24795),
            .I(N__24792));
    LocalMux I__4337 (
            .O(N__24792),
            .I(N__24789));
    Span4Mux_h I__4336 (
            .O(N__24789),
            .I(N__24786));
    Odrv4 I__4335 (
            .O(N__24786),
            .I(\b2v_inst11.count_off_0_9 ));
    CascadeMux I__4334 (
            .O(N__24783),
            .I(\b2v_inst11.N_76_cascade_ ));
    InMux I__4333 (
            .O(N__24780),
            .I(N__24777));
    LocalMux I__4332 (
            .O(N__24777),
            .I(\b2v_inst11.func_state_RNICMPB4Z0Z_0 ));
    CascadeMux I__4331 (
            .O(N__24774),
            .I(\b2v_inst11.func_state_1_m2_1_cascade_ ));
    CascadeMux I__4330 (
            .O(N__24771),
            .I(\b2v_inst11.func_state_cascade_ ));
    InMux I__4329 (
            .O(N__24768),
            .I(N__24765));
    LocalMux I__4328 (
            .O(N__24765),
            .I(\b2v_inst11.N_339 ));
    CascadeMux I__4327 (
            .O(N__24762),
            .I(\b2v_inst11.N_339_cascade_ ));
    InMux I__4326 (
            .O(N__24759),
            .I(N__24756));
    LocalMux I__4325 (
            .O(N__24756),
            .I(\b2v_inst11.func_state_RNI6IFF4Z0Z_1 ));
    InMux I__4324 (
            .O(N__24753),
            .I(N__24750));
    LocalMux I__4323 (
            .O(N__24750),
            .I(N__24747));
    Span4Mux_v I__4322 (
            .O(N__24747),
            .I(N__24744));
    Odrv4 I__4321 (
            .O(N__24744),
            .I(\b2v_inst36.DSW_PWROK_0 ));
    InMux I__4320 (
            .O(N__24741),
            .I(N__24738));
    LocalMux I__4319 (
            .O(N__24738),
            .I(\b2v_inst36.curr_state_RNI3E27Z0Z_0 ));
    IoInMux I__4318 (
            .O(N__24735),
            .I(N__24732));
    LocalMux I__4317 (
            .O(N__24732),
            .I(N__24729));
    Span4Mux_s2_h I__4316 (
            .O(N__24729),
            .I(N__24726));
    Span4Mux_h I__4315 (
            .O(N__24726),
            .I(N__24723));
    Odrv4 I__4314 (
            .O(N__24723),
            .I(dsw_pwrok));
    CascadeMux I__4313 (
            .O(N__24720),
            .I(curr_state_RNID8DP1_0_0_cascade_));
    InMux I__4312 (
            .O(N__24717),
            .I(N__24708));
    InMux I__4311 (
            .O(N__24716),
            .I(N__24708));
    InMux I__4310 (
            .O(N__24715),
            .I(N__24708));
    LocalMux I__4309 (
            .O(N__24708),
            .I(N_413));
    InMux I__4308 (
            .O(N__24705),
            .I(N__24702));
    LocalMux I__4307 (
            .O(N__24702),
            .I(\b2v_inst5.curr_state_0_0 ));
    CascadeMux I__4306 (
            .O(N__24699),
            .I(N__24695));
    CascadeMux I__4305 (
            .O(N__24698),
            .I(N__24691));
    InMux I__4304 (
            .O(N__24695),
            .I(N__24684));
    InMux I__4303 (
            .O(N__24694),
            .I(N__24684));
    InMux I__4302 (
            .O(N__24691),
            .I(N__24684));
    LocalMux I__4301 (
            .O(N__24684),
            .I(\b2v_inst5.curr_stateZ0Z_0 ));
    InMux I__4300 (
            .O(N__24681),
            .I(N__24674));
    InMux I__4299 (
            .O(N__24680),
            .I(N__24674));
    InMux I__4298 (
            .O(N__24679),
            .I(N__24671));
    LocalMux I__4297 (
            .O(N__24674),
            .I(\b2v_inst5.N_2856_i ));
    LocalMux I__4296 (
            .O(N__24671),
            .I(\b2v_inst5.N_2856_i ));
    InMux I__4295 (
            .O(N__24666),
            .I(N__24659));
    InMux I__4294 (
            .O(N__24665),
            .I(N__24650));
    InMux I__4293 (
            .O(N__24664),
            .I(N__24650));
    InMux I__4292 (
            .O(N__24663),
            .I(N__24650));
    InMux I__4291 (
            .O(N__24662),
            .I(N__24650));
    LocalMux I__4290 (
            .O(N__24659),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1 ));
    LocalMux I__4289 (
            .O(N__24650),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1 ));
    CascadeMux I__4288 (
            .O(N__24645),
            .I(\b2v_inst5.N_2856_i_cascade_ ));
    InMux I__4287 (
            .O(N__24642),
            .I(N__24639));
    LocalMux I__4286 (
            .O(N__24639),
            .I(N__24636));
    Odrv4 I__4285 (
            .O(N__24636),
            .I(\b2v_inst11.count_off_0_7 ));
    CascadeMux I__4284 (
            .O(N__24633),
            .I(N__24629));
    InMux I__4283 (
            .O(N__24632),
            .I(N__24626));
    InMux I__4282 (
            .O(N__24629),
            .I(N__24623));
    LocalMux I__4281 (
            .O(N__24626),
            .I(N__24620));
    LocalMux I__4280 (
            .O(N__24623),
            .I(N__24617));
    Span4Mux_h I__4279 (
            .O(N__24620),
            .I(N__24614));
    Odrv4 I__4278 (
            .O(N__24617),
            .I(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ));
    Odrv4 I__4277 (
            .O(N__24614),
            .I(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ));
    CascadeMux I__4276 (
            .O(N__24609),
            .I(N__24606));
    InMux I__4275 (
            .O(N__24606),
            .I(N__24602));
    InMux I__4274 (
            .O(N__24605),
            .I(N__24599));
    LocalMux I__4273 (
            .O(N__24602),
            .I(N__24596));
    LocalMux I__4272 (
            .O(N__24599),
            .I(\b2v_inst11.count_offZ0Z_7 ));
    Odrv4 I__4271 (
            .O(N__24596),
            .I(\b2v_inst11.count_offZ0Z_7 ));
    InMux I__4270 (
            .O(N__24591),
            .I(N__24588));
    LocalMux I__4269 (
            .O(N__24588),
            .I(N__24585));
    Span4Mux_h I__4268 (
            .O(N__24585),
            .I(N__24582));
    Odrv4 I__4267 (
            .O(N__24582),
            .I(\b2v_inst11.un34_clk_100khz_11 ));
    InMux I__4266 (
            .O(N__24579),
            .I(N__24576));
    LocalMux I__4265 (
            .O(N__24576),
            .I(\b2v_inst11.un34_clk_100khz_9 ));
    CascadeMux I__4264 (
            .O(N__24573),
            .I(N__24570));
    InMux I__4263 (
            .O(N__24570),
            .I(N__24567));
    LocalMux I__4262 (
            .O(N__24567),
            .I(N__24564));
    Span4Mux_h I__4261 (
            .O(N__24564),
            .I(N__24561));
    Odrv4 I__4260 (
            .O(N__24561),
            .I(\b2v_inst11.un34_clk_100khz_10 ));
    InMux I__4259 (
            .O(N__24558),
            .I(N__24555));
    LocalMux I__4258 (
            .O(N__24555),
            .I(\b2v_inst11.un34_clk_100khz_8 ));
    CascadeMux I__4257 (
            .O(N__24552),
            .I(\b2v_inst11.count_off_RNI_1Z0Z_1_cascade_ ));
    CascadeMux I__4256 (
            .O(N__24549),
            .I(\b2v_inst11.func_state_1_m0_0_0_1_cascade_ ));
    InMux I__4255 (
            .O(N__24546),
            .I(N__24540));
    InMux I__4254 (
            .O(N__24545),
            .I(N__24540));
    LocalMux I__4253 (
            .O(N__24540),
            .I(N__24537));
    Odrv4 I__4252 (
            .O(N__24537),
            .I(\b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ));
    CascadeMux I__4251 (
            .O(N__24534),
            .I(N__24531));
    InMux I__4250 (
            .O(N__24531),
            .I(N__24528));
    LocalMux I__4249 (
            .O(N__24528),
            .I(\b2v_inst11.count_off_0_8 ));
    InMux I__4248 (
            .O(N__24525),
            .I(N__24522));
    LocalMux I__4247 (
            .O(N__24522),
            .I(N__24518));
    InMux I__4246 (
            .O(N__24521),
            .I(N__24515));
    Odrv4 I__4245 (
            .O(N__24518),
            .I(\b2v_inst11.count_offZ0Z_8 ));
    LocalMux I__4244 (
            .O(N__24515),
            .I(\b2v_inst11.count_offZ0Z_8 ));
    CascadeMux I__4243 (
            .O(N__24510),
            .I(\b2v_inst5.curr_stateZ0Z_1_cascade_ ));
    InMux I__4242 (
            .O(N__24507),
            .I(N__24501));
    InMux I__4241 (
            .O(N__24506),
            .I(N__24501));
    LocalMux I__4240 (
            .O(N__24501),
            .I(\b2v_inst5.count_1_0 ));
    CascadeMux I__4239 (
            .O(N__24498),
            .I(N__24495));
    InMux I__4238 (
            .O(N__24495),
            .I(N__24489));
    InMux I__4237 (
            .O(N__24494),
            .I(N__24489));
    LocalMux I__4236 (
            .O(N__24489),
            .I(\b2v_inst5.count_rst_14 ));
    InMux I__4235 (
            .O(N__24486),
            .I(N__24479));
    InMux I__4234 (
            .O(N__24485),
            .I(N__24479));
    InMux I__4233 (
            .O(N__24484),
            .I(N__24476));
    LocalMux I__4232 (
            .O(N__24479),
            .I(\b2v_inst5.count_i_0 ));
    LocalMux I__4231 (
            .O(N__24476),
            .I(\b2v_inst5.count_i_0 ));
    InMux I__4230 (
            .O(N__24471),
            .I(N__24468));
    LocalMux I__4229 (
            .O(N__24468),
            .I(\b2v_inst5.curr_stateZ0Z_1 ));
    InMux I__4228 (
            .O(N__24465),
            .I(N__24462));
    LocalMux I__4227 (
            .O(N__24462),
            .I(N__24459));
    Odrv12 I__4226 (
            .O(N__24459),
            .I(\b2v_inst5.count_1_15 ));
    InMux I__4225 (
            .O(N__24456),
            .I(N__24453));
    LocalMux I__4224 (
            .O(N__24453),
            .I(N__24450));
    Span4Mux_s0_v I__4223 (
            .O(N__24450),
            .I(N__24446));
    InMux I__4222 (
            .O(N__24449),
            .I(N__24443));
    Odrv4 I__4221 (
            .O(N__24446),
            .I(\b2v_inst5.count_rst ));
    LocalMux I__4220 (
            .O(N__24443),
            .I(\b2v_inst5.count_rst ));
    InMux I__4219 (
            .O(N__24438),
            .I(N__24435));
    LocalMux I__4218 (
            .O(N__24435),
            .I(N__24431));
    InMux I__4217 (
            .O(N__24434),
            .I(N__24428));
    Odrv4 I__4216 (
            .O(N__24431),
            .I(\b2v_inst5.countZ0Z_15 ));
    LocalMux I__4215 (
            .O(N__24428),
            .I(\b2v_inst5.countZ0Z_15 ));
    CascadeMux I__4214 (
            .O(N__24423),
            .I(\b2v_inst5.curr_stateZ0Z_0_cascade_ ));
    InMux I__4213 (
            .O(N__24420),
            .I(N__24414));
    InMux I__4212 (
            .O(N__24419),
            .I(N__24414));
    LocalMux I__4211 (
            .O(N__24414),
            .I(\b2v_inst5.N_51 ));
    InMux I__4210 (
            .O(N__24411),
            .I(N__24408));
    LocalMux I__4209 (
            .O(N__24408),
            .I(\b2v_inst5.m4_0 ));
    InMux I__4208 (
            .O(N__24405),
            .I(N__24399));
    InMux I__4207 (
            .O(N__24404),
            .I(N__24399));
    LocalMux I__4206 (
            .O(N__24399),
            .I(\b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2 ));
    CascadeMux I__4205 (
            .O(N__24396),
            .I(N__24393));
    InMux I__4204 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__4203 (
            .O(N__24390),
            .I(\b2v_inst5.count_1_12 ));
    InMux I__4202 (
            .O(N__24387),
            .I(N__24384));
    LocalMux I__4201 (
            .O(N__24384),
            .I(\b2v_inst5.count_1_14 ));
    InMux I__4200 (
            .O(N__24381),
            .I(N__24375));
    InMux I__4199 (
            .O(N__24380),
            .I(N__24375));
    LocalMux I__4198 (
            .O(N__24375),
            .I(\b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ));
    InMux I__4197 (
            .O(N__24372),
            .I(N__24369));
    LocalMux I__4196 (
            .O(N__24369),
            .I(\b2v_inst5.countZ0Z_14 ));
    CascadeMux I__4195 (
            .O(N__24366),
            .I(\b2v_inst5.countZ0Z_14_cascade_ ));
    InMux I__4194 (
            .O(N__24363),
            .I(N__24359));
    InMux I__4193 (
            .O(N__24362),
            .I(N__24356));
    LocalMux I__4192 (
            .O(N__24359),
            .I(\b2v_inst5.countZ0Z_12 ));
    LocalMux I__4191 (
            .O(N__24356),
            .I(\b2v_inst5.countZ0Z_12 ));
    CascadeMux I__4190 (
            .O(N__24351),
            .I(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_ ));
    InMux I__4189 (
            .O(N__24348),
            .I(N__24345));
    LocalMux I__4188 (
            .O(N__24345),
            .I(\b2v_inst5.un2_count_1_axb_0 ));
    InMux I__4187 (
            .O(N__24342),
            .I(N__24339));
    LocalMux I__4186 (
            .O(N__24339),
            .I(\b2v_inst5.curr_state_0_1 ));
    InMux I__4185 (
            .O(N__24336),
            .I(N__24330));
    InMux I__4184 (
            .O(N__24335),
            .I(N__24330));
    LocalMux I__4183 (
            .O(N__24330),
            .I(\b2v_inst5.un2_count_1_cry_4_c_RNIPKTZ0Z9 ));
    CascadeMux I__4182 (
            .O(N__24327),
            .I(N__24324));
    InMux I__4181 (
            .O(N__24324),
            .I(N__24321));
    LocalMux I__4180 (
            .O(N__24321),
            .I(\b2v_inst5.count_1_5 ));
    InMux I__4179 (
            .O(N__24318),
            .I(N__24314));
    InMux I__4178 (
            .O(N__24317),
            .I(N__24311));
    LocalMux I__4177 (
            .O(N__24314),
            .I(\b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9 ));
    LocalMux I__4176 (
            .O(N__24311),
            .I(\b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9 ));
    CascadeMux I__4175 (
            .O(N__24306),
            .I(N__24303));
    InMux I__4174 (
            .O(N__24303),
            .I(N__24300));
    LocalMux I__4173 (
            .O(N__24300),
            .I(\b2v_inst5.count_1_6 ));
    CascadeMux I__4172 (
            .O(N__24297),
            .I(\b2v_inst5.countZ0Z_13_cascade_ ));
    InMux I__4171 (
            .O(N__24294),
            .I(N__24291));
    LocalMux I__4170 (
            .O(N__24291),
            .I(\b2v_inst5.count_1_13 ));
    InMux I__4169 (
            .O(N__24288),
            .I(N__24285));
    LocalMux I__4168 (
            .O(N__24285),
            .I(\b2v_inst5.countZ0Z_3 ));
    CascadeMux I__4167 (
            .O(N__24282),
            .I(\b2v_inst5.countZ0Z_3_cascade_ ));
    InMux I__4166 (
            .O(N__24279),
            .I(N__24276));
    LocalMux I__4165 (
            .O(N__24276),
            .I(N__24272));
    InMux I__4164 (
            .O(N__24275),
            .I(N__24269));
    Odrv4 I__4163 (
            .O(N__24272),
            .I(\b2v_inst5.countZ0Z_1 ));
    LocalMux I__4162 (
            .O(N__24269),
            .I(\b2v_inst5.countZ0Z_1 ));
    InMux I__4161 (
            .O(N__24264),
            .I(N__24258));
    InMux I__4160 (
            .O(N__24263),
            .I(N__24258));
    LocalMux I__4159 (
            .O(N__24258),
            .I(N__24255));
    Odrv4 I__4158 (
            .O(N__24255),
            .I(\b2v_inst5.un2_count_1_cry_0_c_RNILCPZ0Z9 ));
    CascadeMux I__4157 (
            .O(N__24252),
            .I(N__24249));
    InMux I__4156 (
            .O(N__24249),
            .I(N__24246));
    LocalMux I__4155 (
            .O(N__24246),
            .I(\b2v_inst5.count_1_1 ));
    CascadeMux I__4154 (
            .O(N__24243),
            .I(N__24240));
    InMux I__4153 (
            .O(N__24240),
            .I(N__24237));
    LocalMux I__4152 (
            .O(N__24237),
            .I(\b2v_inst11.mult1_un75_sum_cry_4_s ));
    InMux I__4151 (
            .O(N__24234),
            .I(\b2v_inst11.mult1_un75_sum_cry_3 ));
    InMux I__4150 (
            .O(N__24231),
            .I(N__24228));
    LocalMux I__4149 (
            .O(N__24228),
            .I(\b2v_inst11.mult1_un75_sum_cry_5_s ));
    InMux I__4148 (
            .O(N__24225),
            .I(\b2v_inst11.mult1_un75_sum_cry_4 ));
    InMux I__4147 (
            .O(N__24222),
            .I(N__24219));
    LocalMux I__4146 (
            .O(N__24219),
            .I(\b2v_inst11.mult1_un75_sum_cry_6_s ));
    InMux I__4145 (
            .O(N__24216),
            .I(\b2v_inst11.mult1_un75_sum_cry_5 ));
    CascadeMux I__4144 (
            .O(N__24213),
            .I(N__24210));
    InMux I__4143 (
            .O(N__24210),
            .I(N__24207));
    LocalMux I__4142 (
            .O(N__24207),
            .I(\b2v_inst11.mult1_un82_sum_axb_8 ));
    InMux I__4141 (
            .O(N__24204),
            .I(\b2v_inst11.mult1_un75_sum_cry_6 ));
    InMux I__4140 (
            .O(N__24201),
            .I(\b2v_inst11.mult1_un75_sum_cry_7 ));
    InMux I__4139 (
            .O(N__24198),
            .I(N__24195));
    LocalMux I__4138 (
            .O(N__24195),
            .I(N__24191));
    CascadeMux I__4137 (
            .O(N__24194),
            .I(N__24187));
    Span4Mux_s3_h I__4136 (
            .O(N__24191),
            .I(N__24182));
    InMux I__4135 (
            .O(N__24190),
            .I(N__24179));
    InMux I__4134 (
            .O(N__24187),
            .I(N__24172));
    InMux I__4133 (
            .O(N__24186),
            .I(N__24172));
    InMux I__4132 (
            .O(N__24185),
            .I(N__24172));
    Odrv4 I__4131 (
            .O(N__24182),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__4130 (
            .O(N__24179),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__4129 (
            .O(N__24172),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    CascadeMux I__4128 (
            .O(N__24165),
            .I(N__24161));
    CascadeMux I__4127 (
            .O(N__24164),
            .I(N__24157));
    InMux I__4126 (
            .O(N__24161),
            .I(N__24150));
    InMux I__4125 (
            .O(N__24160),
            .I(N__24150));
    InMux I__4124 (
            .O(N__24157),
            .I(N__24150));
    LocalMux I__4123 (
            .O(N__24150),
            .I(\b2v_inst11.mult1_un68_sum_i_0_8 ));
    CascadeMux I__4122 (
            .O(N__24147),
            .I(N__24144));
    InMux I__4121 (
            .O(N__24144),
            .I(N__24141));
    LocalMux I__4120 (
            .O(N__24141),
            .I(\b2v_inst11.mult1_un82_sum_cry_4_s ));
    InMux I__4119 (
            .O(N__24138),
            .I(\b2v_inst11.mult1_un82_sum_cry_3 ));
    InMux I__4118 (
            .O(N__24135),
            .I(N__24132));
    LocalMux I__4117 (
            .O(N__24132),
            .I(\b2v_inst11.mult1_un82_sum_cry_5_s ));
    InMux I__4116 (
            .O(N__24129),
            .I(\b2v_inst11.mult1_un82_sum_cry_4 ));
    InMux I__4115 (
            .O(N__24126),
            .I(N__24123));
    LocalMux I__4114 (
            .O(N__24123),
            .I(\b2v_inst11.mult1_un82_sum_cry_6_s ));
    InMux I__4113 (
            .O(N__24120),
            .I(\b2v_inst11.mult1_un82_sum_cry_5 ));
    CascadeMux I__4112 (
            .O(N__24117),
            .I(N__24114));
    InMux I__4111 (
            .O(N__24114),
            .I(N__24111));
    LocalMux I__4110 (
            .O(N__24111),
            .I(\b2v_inst11.mult1_un89_sum_axb_8 ));
    InMux I__4109 (
            .O(N__24108),
            .I(\b2v_inst11.mult1_un82_sum_cry_6 ));
    InMux I__4108 (
            .O(N__24105),
            .I(\b2v_inst11.mult1_un82_sum_cry_7 ));
    InMux I__4107 (
            .O(N__24102),
            .I(N__24099));
    LocalMux I__4106 (
            .O(N__24099),
            .I(N__24095));
    CascadeMux I__4105 (
            .O(N__24098),
            .I(N__24091));
    Span4Mux_s2_v I__4104 (
            .O(N__24095),
            .I(N__24086));
    InMux I__4103 (
            .O(N__24094),
            .I(N__24083));
    InMux I__4102 (
            .O(N__24091),
            .I(N__24076));
    InMux I__4101 (
            .O(N__24090),
            .I(N__24076));
    InMux I__4100 (
            .O(N__24089),
            .I(N__24076));
    Odrv4 I__4099 (
            .O(N__24086),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__4098 (
            .O(N__24083),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__4097 (
            .O(N__24076),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    CascadeMux I__4096 (
            .O(N__24069),
            .I(N__24065));
    CascadeMux I__4095 (
            .O(N__24068),
            .I(N__24061));
    InMux I__4094 (
            .O(N__24065),
            .I(N__24054));
    InMux I__4093 (
            .O(N__24064),
            .I(N__24054));
    InMux I__4092 (
            .O(N__24061),
            .I(N__24054));
    LocalMux I__4091 (
            .O(N__24054),
            .I(\b2v_inst11.mult1_un75_sum_i_0_8 ));
    InMux I__4090 (
            .O(N__24051),
            .I(N__24048));
    LocalMux I__4089 (
            .O(N__24048),
            .I(N__24045));
    Odrv4 I__4088 (
            .O(N__24045),
            .I(\b2v_inst11.mult1_un68_sum_i ));
    CascadeMux I__4087 (
            .O(N__24042),
            .I(N__24039));
    InMux I__4086 (
            .O(N__24039),
            .I(N__24036));
    LocalMux I__4085 (
            .O(N__24036),
            .I(\b2v_inst11.mult1_un75_sum_cry_3_s ));
    InMux I__4084 (
            .O(N__24033),
            .I(\b2v_inst11.mult1_un75_sum_cry_2 ));
    InMux I__4083 (
            .O(N__24030),
            .I(\b2v_inst11.mult1_un152_sum_cry_7 ));
    InMux I__4082 (
            .O(N__24027),
            .I(N__24024));
    LocalMux I__4081 (
            .O(N__24024),
            .I(N__24021));
    Span4Mux_s2_h I__4080 (
            .O(N__24021),
            .I(N__24017));
    CascadeMux I__4079 (
            .O(N__24020),
            .I(N__24013));
    Span4Mux_h I__4078 (
            .O(N__24017),
            .I(N__24009));
    InMux I__4077 (
            .O(N__24016),
            .I(N__24004));
    InMux I__4076 (
            .O(N__24013),
            .I(N__24004));
    InMux I__4075 (
            .O(N__24012),
            .I(N__24001));
    Odrv4 I__4074 (
            .O(N__24009),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__4073 (
            .O(N__24004),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__4072 (
            .O(N__24001),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    CascadeMux I__4071 (
            .O(N__23994),
            .I(\b2v_inst11.mult1_un152_sum_s_8_cascade_ ));
    CascadeMux I__4070 (
            .O(N__23991),
            .I(N__23987));
    CascadeMux I__4069 (
            .O(N__23990),
            .I(N__23983));
    InMux I__4068 (
            .O(N__23987),
            .I(N__23976));
    InMux I__4067 (
            .O(N__23986),
            .I(N__23976));
    InMux I__4066 (
            .O(N__23983),
            .I(N__23976));
    LocalMux I__4065 (
            .O(N__23976),
            .I(\b2v_inst11.mult1_un152_sum_i_0_8 ));
    InMux I__4064 (
            .O(N__23973),
            .I(N__23970));
    LocalMux I__4063 (
            .O(N__23970),
            .I(N__23967));
    Odrv4 I__4062 (
            .O(N__23967),
            .I(\b2v_inst11.mult1_un82_sum_i ));
    InMux I__4061 (
            .O(N__23964),
            .I(N__23961));
    LocalMux I__4060 (
            .O(N__23961),
            .I(N__23958));
    Span4Mux_h I__4059 (
            .O(N__23958),
            .I(N__23955));
    Odrv4 I__4058 (
            .O(N__23955),
            .I(\b2v_inst11.mult1_un96_sum_i ));
    IoInMux I__4057 (
            .O(N__23952),
            .I(N__23949));
    LocalMux I__4056 (
            .O(N__23949),
            .I(N__23946));
    Span4Mux_s3_h I__4055 (
            .O(N__23946),
            .I(N__23942));
    IoInMux I__4054 (
            .O(N__23945),
            .I(N__23938));
    Span4Mux_v I__4053 (
            .O(N__23942),
            .I(N__23935));
    IoInMux I__4052 (
            .O(N__23941),
            .I(N__23932));
    LocalMux I__4051 (
            .O(N__23938),
            .I(N__23929));
    Sp12to4 I__4050 (
            .O(N__23935),
            .I(N__23926));
    LocalMux I__4049 (
            .O(N__23932),
            .I(N__23923));
    IoSpan4Mux I__4048 (
            .O(N__23929),
            .I(N__23920));
    Span12Mux_s5_h I__4047 (
            .O(N__23926),
            .I(N__23915));
    Span12Mux_s5_v I__4046 (
            .O(N__23923),
            .I(N__23915));
    Sp12to4 I__4045 (
            .O(N__23920),
            .I(N__23912));
    Odrv12 I__4044 (
            .O(N__23915),
            .I(pch_pwrok));
    Odrv12 I__4043 (
            .O(N__23912),
            .I(pch_pwrok));
    InMux I__4042 (
            .O(N__23907),
            .I(N__23904));
    LocalMux I__4041 (
            .O(N__23904),
            .I(N__23901));
    Odrv4 I__4040 (
            .O(N__23901),
            .I(\b2v_inst11.mult1_un75_sum_i ));
    CascadeMux I__4039 (
            .O(N__23898),
            .I(N__23895));
    InMux I__4038 (
            .O(N__23895),
            .I(N__23892));
    LocalMux I__4037 (
            .O(N__23892),
            .I(\b2v_inst11.mult1_un82_sum_cry_3_s ));
    InMux I__4036 (
            .O(N__23889),
            .I(\b2v_inst11.mult1_un82_sum_cry_2 ));
    InMux I__4035 (
            .O(N__23886),
            .I(N__23882));
    CascadeMux I__4034 (
            .O(N__23885),
            .I(N__23879));
    LocalMux I__4033 (
            .O(N__23882),
            .I(N__23874));
    InMux I__4032 (
            .O(N__23879),
            .I(N__23866));
    InMux I__4031 (
            .O(N__23878),
            .I(N__23866));
    InMux I__4030 (
            .O(N__23877),
            .I(N__23866));
    Span4Mux_h I__4029 (
            .O(N__23874),
            .I(N__23863));
    InMux I__4028 (
            .O(N__23873),
            .I(N__23860));
    LocalMux I__4027 (
            .O(N__23866),
            .I(N__23857));
    Odrv4 I__4026 (
            .O(N__23863),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    LocalMux I__4025 (
            .O(N__23860),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    Odrv4 I__4024 (
            .O(N__23857),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    InMux I__4023 (
            .O(N__23850),
            .I(N__23847));
    LocalMux I__4022 (
            .O(N__23847),
            .I(N__23844));
    Odrv4 I__4021 (
            .O(N__23844),
            .I(\b2v_inst11.mult1_un159_sum_i ));
    CascadeMux I__4020 (
            .O(N__23841),
            .I(N__23838));
    InMux I__4019 (
            .O(N__23838),
            .I(N__23835));
    LocalMux I__4018 (
            .O(N__23835),
            .I(\b2v_inst11.mult1_un145_sum_i_0_8 ));
    CascadeMux I__4017 (
            .O(N__23832),
            .I(N__23829));
    InMux I__4016 (
            .O(N__23829),
            .I(N__23826));
    LocalMux I__4015 (
            .O(N__23826),
            .I(\b2v_inst11.mult1_un152_sum_cry_3_s ));
    InMux I__4014 (
            .O(N__23823),
            .I(\b2v_inst11.mult1_un152_sum_cry_2 ));
    InMux I__4013 (
            .O(N__23820),
            .I(N__23816));
    InMux I__4012 (
            .O(N__23819),
            .I(N__23813));
    LocalMux I__4011 (
            .O(N__23816),
            .I(N__23810));
    LocalMux I__4010 (
            .O(N__23813),
            .I(\b2v_inst11.mult1_un145_sum_cry_3_s ));
    Odrv12 I__4009 (
            .O(N__23810),
            .I(\b2v_inst11.mult1_un145_sum_cry_3_s ));
    CascadeMux I__4008 (
            .O(N__23805),
            .I(N__23802));
    InMux I__4007 (
            .O(N__23802),
            .I(N__23799));
    LocalMux I__4006 (
            .O(N__23799),
            .I(\b2v_inst11.mult1_un152_sum_axb_4_l_fx ));
    InMux I__4005 (
            .O(N__23796),
            .I(N__23793));
    LocalMux I__4004 (
            .O(N__23793),
            .I(\b2v_inst11.mult1_un152_sum_cry_4_s ));
    InMux I__4003 (
            .O(N__23790),
            .I(\b2v_inst11.mult1_un152_sum_cry_3 ));
    InMux I__4002 (
            .O(N__23787),
            .I(N__23784));
    LocalMux I__4001 (
            .O(N__23784),
            .I(N__23781));
    Odrv4 I__4000 (
            .O(N__23781),
            .I(\b2v_inst11.mult1_un145_sum_cry_4_s ));
    CascadeMux I__3999 (
            .O(N__23778),
            .I(N__23775));
    InMux I__3998 (
            .O(N__23775),
            .I(N__23772));
    LocalMux I__3997 (
            .O(N__23772),
            .I(\b2v_inst11.mult1_un152_sum_cry_5_s ));
    InMux I__3996 (
            .O(N__23769),
            .I(\b2v_inst11.mult1_un152_sum_cry_4 ));
    InMux I__3995 (
            .O(N__23766),
            .I(N__23762));
    CascadeMux I__3994 (
            .O(N__23765),
            .I(N__23758));
    LocalMux I__3993 (
            .O(N__23762),
            .I(N__23755));
    InMux I__3992 (
            .O(N__23761),
            .I(N__23750));
    InMux I__3991 (
            .O(N__23758),
            .I(N__23750));
    Span4Mux_v I__3990 (
            .O(N__23755),
            .I(N__23741));
    LocalMux I__3989 (
            .O(N__23750),
            .I(N__23741));
    InMux I__3988 (
            .O(N__23749),
            .I(N__23738));
    InMux I__3987 (
            .O(N__23748),
            .I(N__23735));
    InMux I__3986 (
            .O(N__23747),
            .I(N__23730));
    InMux I__3985 (
            .O(N__23746),
            .I(N__23730));
    Odrv4 I__3984 (
            .O(N__23741),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__3983 (
            .O(N__23738),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__3982 (
            .O(N__23735),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__3981 (
            .O(N__23730),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    CascadeMux I__3980 (
            .O(N__23721),
            .I(N__23718));
    InMux I__3979 (
            .O(N__23718),
            .I(N__23715));
    LocalMux I__3978 (
            .O(N__23715),
            .I(N__23712));
    Odrv4 I__3977 (
            .O(N__23712),
            .I(\b2v_inst11.mult1_un145_sum_cry_5_s ));
    InMux I__3976 (
            .O(N__23709),
            .I(N__23706));
    LocalMux I__3975 (
            .O(N__23706),
            .I(\b2v_inst11.mult1_un152_sum_cry_6_s ));
    InMux I__3974 (
            .O(N__23703),
            .I(\b2v_inst11.mult1_un152_sum_cry_5 ));
    InMux I__3973 (
            .O(N__23700),
            .I(N__23696));
    InMux I__3972 (
            .O(N__23699),
            .I(N__23693));
    LocalMux I__3971 (
            .O(N__23696),
            .I(N__23690));
    LocalMux I__3970 (
            .O(N__23693),
            .I(\b2v_inst11.mult1_un145_sum_cry_6_s ));
    Odrv4 I__3969 (
            .O(N__23690),
            .I(\b2v_inst11.mult1_un145_sum_cry_6_s ));
    CascadeMux I__3968 (
            .O(N__23685),
            .I(N__23682));
    InMux I__3967 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__3966 (
            .O(N__23679),
            .I(\b2v_inst11.mult1_un152_sum_axb_7_l_fx ));
    CascadeMux I__3965 (
            .O(N__23676),
            .I(N__23673));
    InMux I__3964 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__3963 (
            .O(N__23670),
            .I(\b2v_inst11.mult1_un159_sum_axb_7 ));
    InMux I__3962 (
            .O(N__23667),
            .I(\b2v_inst11.mult1_un152_sum_cry_6 ));
    CascadeMux I__3961 (
            .O(N__23664),
            .I(N__23661));
    InMux I__3960 (
            .O(N__23661),
            .I(N__23658));
    LocalMux I__3959 (
            .O(N__23658),
            .I(N__23655));
    Odrv4 I__3958 (
            .O(N__23655),
            .I(\b2v_inst11.mult1_un152_sum_axb_8 ));
    InMux I__3957 (
            .O(N__23652),
            .I(N__23648));
    InMux I__3956 (
            .O(N__23651),
            .I(N__23645));
    LocalMux I__3955 (
            .O(N__23648),
            .I(\b2v_inst20.counterZ0Z_24 ));
    LocalMux I__3954 (
            .O(N__23645),
            .I(\b2v_inst20.counterZ0Z_24 ));
    InMux I__3953 (
            .O(N__23640),
            .I(N__23636));
    InMux I__3952 (
            .O(N__23639),
            .I(N__23633));
    LocalMux I__3951 (
            .O(N__23636),
            .I(N__23630));
    LocalMux I__3950 (
            .O(N__23633),
            .I(\b2v_inst20.counterZ0Z_26 ));
    Odrv4 I__3949 (
            .O(N__23630),
            .I(\b2v_inst20.counterZ0Z_26 ));
    CascadeMux I__3948 (
            .O(N__23625),
            .I(N__23622));
    InMux I__3947 (
            .O(N__23622),
            .I(N__23618));
    InMux I__3946 (
            .O(N__23621),
            .I(N__23615));
    LocalMux I__3945 (
            .O(N__23618),
            .I(N__23612));
    LocalMux I__3944 (
            .O(N__23615),
            .I(\b2v_inst20.counterZ0Z_25 ));
    Odrv4 I__3943 (
            .O(N__23612),
            .I(\b2v_inst20.counterZ0Z_25 ));
    InMux I__3942 (
            .O(N__23607),
            .I(N__23603));
    InMux I__3941 (
            .O(N__23606),
            .I(N__23600));
    LocalMux I__3940 (
            .O(N__23603),
            .I(N__23597));
    LocalMux I__3939 (
            .O(N__23600),
            .I(\b2v_inst20.counterZ0Z_27 ));
    Odrv4 I__3938 (
            .O(N__23597),
            .I(\b2v_inst20.counterZ0Z_27 ));
    InMux I__3937 (
            .O(N__23592),
            .I(N__23589));
    LocalMux I__3936 (
            .O(N__23589),
            .I(\b2v_inst20.un4_counter_6_and ));
    CascadeMux I__3935 (
            .O(N__23586),
            .I(N__23583));
    InMux I__3934 (
            .O(N__23583),
            .I(N__23580));
    LocalMux I__3933 (
            .O(N__23580),
            .I(N__23577));
    Odrv4 I__3932 (
            .O(N__23577),
            .I(\b2v_inst11.mult1_un159_sum_cry_2_s ));
    InMux I__3931 (
            .O(N__23574),
            .I(\b2v_inst11.mult1_un159_sum_cry_1 ));
    CascadeMux I__3930 (
            .O(N__23571),
            .I(N__23568));
    InMux I__3929 (
            .O(N__23568),
            .I(N__23565));
    LocalMux I__3928 (
            .O(N__23565),
            .I(N__23562));
    Odrv4 I__3927 (
            .O(N__23562),
            .I(\b2v_inst11.mult1_un159_sum_cry_3_s ));
    InMux I__3926 (
            .O(N__23559),
            .I(\b2v_inst11.mult1_un159_sum_cry_2 ));
    InMux I__3925 (
            .O(N__23556),
            .I(N__23553));
    LocalMux I__3924 (
            .O(N__23553),
            .I(N__23550));
    Odrv4 I__3923 (
            .O(N__23550),
            .I(\b2v_inst11.mult1_un159_sum_cry_4_s ));
    InMux I__3922 (
            .O(N__23547),
            .I(\b2v_inst11.mult1_un159_sum_cry_3 ));
    InMux I__3921 (
            .O(N__23544),
            .I(N__23541));
    LocalMux I__3920 (
            .O(N__23541),
            .I(N__23538));
    Odrv4 I__3919 (
            .O(N__23538),
            .I(\b2v_inst11.mult1_un159_sum_cry_5_s ));
    InMux I__3918 (
            .O(N__23535),
            .I(\b2v_inst11.mult1_un159_sum_cry_4 ));
    InMux I__3917 (
            .O(N__23532),
            .I(N__23529));
    LocalMux I__3916 (
            .O(N__23529),
            .I(N__23526));
    Odrv4 I__3915 (
            .O(N__23526),
            .I(\b2v_inst11.mult1_un166_sum_axb_6 ));
    InMux I__3914 (
            .O(N__23523),
            .I(\b2v_inst11.mult1_un159_sum_cry_5 ));
    InMux I__3913 (
            .O(N__23520),
            .I(\b2v_inst11.mult1_un159_sum_cry_6 ));
    InMux I__3912 (
            .O(N__23517),
            .I(N__23514));
    LocalMux I__3911 (
            .O(N__23514),
            .I(N__23511));
    Span4Mux_h I__3910 (
            .O(N__23511),
            .I(N__23508));
    Odrv4 I__3909 (
            .O(N__23508),
            .I(\b2v_inst20.un4_counter_5_and ));
    InMux I__3908 (
            .O(N__23505),
            .I(N__23502));
    LocalMux I__3907 (
            .O(N__23502),
            .I(\b2v_inst20.un4_counter_7_and ));
    InMux I__3906 (
            .O(N__23499),
            .I(bfn_6_10_0_));
    InMux I__3905 (
            .O(N__23496),
            .I(N__23492));
    InMux I__3904 (
            .O(N__23495),
            .I(N__23489));
    LocalMux I__3903 (
            .O(N__23492),
            .I(\b2v_inst20.counterZ0Z_16 ));
    LocalMux I__3902 (
            .O(N__23489),
            .I(\b2v_inst20.counterZ0Z_16 ));
    InMux I__3901 (
            .O(N__23484),
            .I(N__23480));
    InMux I__3900 (
            .O(N__23483),
            .I(N__23477));
    LocalMux I__3899 (
            .O(N__23480),
            .I(\b2v_inst20.counterZ0Z_17 ));
    LocalMux I__3898 (
            .O(N__23477),
            .I(\b2v_inst20.counterZ0Z_17 ));
    CascadeMux I__3897 (
            .O(N__23472),
            .I(N__23468));
    InMux I__3896 (
            .O(N__23471),
            .I(N__23465));
    InMux I__3895 (
            .O(N__23468),
            .I(N__23462));
    LocalMux I__3894 (
            .O(N__23465),
            .I(\b2v_inst20.counterZ0Z_18 ));
    LocalMux I__3893 (
            .O(N__23462),
            .I(\b2v_inst20.counterZ0Z_18 ));
    InMux I__3892 (
            .O(N__23457),
            .I(N__23453));
    InMux I__3891 (
            .O(N__23456),
            .I(N__23450));
    LocalMux I__3890 (
            .O(N__23453),
            .I(\b2v_inst20.counterZ0Z_19 ));
    LocalMux I__3889 (
            .O(N__23450),
            .I(\b2v_inst20.counterZ0Z_19 ));
    InMux I__3888 (
            .O(N__23445),
            .I(N__23442));
    LocalMux I__3887 (
            .O(N__23442),
            .I(\b2v_inst20.un4_counter_4_and ));
    InMux I__3886 (
            .O(N__23439),
            .I(N__23435));
    InMux I__3885 (
            .O(N__23438),
            .I(N__23432));
    LocalMux I__3884 (
            .O(N__23435),
            .I(\b2v_inst20.counterZ0Z_15 ));
    LocalMux I__3883 (
            .O(N__23432),
            .I(\b2v_inst20.counterZ0Z_15 ));
    InMux I__3882 (
            .O(N__23427),
            .I(N__23423));
    InMux I__3881 (
            .O(N__23426),
            .I(N__23420));
    LocalMux I__3880 (
            .O(N__23423),
            .I(\b2v_inst20.counterZ0Z_13 ));
    LocalMux I__3879 (
            .O(N__23420),
            .I(\b2v_inst20.counterZ0Z_13 ));
    CascadeMux I__3878 (
            .O(N__23415),
            .I(N__23411));
    InMux I__3877 (
            .O(N__23414),
            .I(N__23408));
    InMux I__3876 (
            .O(N__23411),
            .I(N__23405));
    LocalMux I__3875 (
            .O(N__23408),
            .I(\b2v_inst20.counterZ0Z_14 ));
    LocalMux I__3874 (
            .O(N__23405),
            .I(\b2v_inst20.counterZ0Z_14 ));
    InMux I__3873 (
            .O(N__23400),
            .I(N__23396));
    InMux I__3872 (
            .O(N__23399),
            .I(N__23393));
    LocalMux I__3871 (
            .O(N__23396),
            .I(\b2v_inst20.counterZ0Z_12 ));
    LocalMux I__3870 (
            .O(N__23393),
            .I(\b2v_inst20.counterZ0Z_12 ));
    InMux I__3869 (
            .O(N__23388),
            .I(N__23385));
    LocalMux I__3868 (
            .O(N__23385),
            .I(\b2v_inst20.un4_counter_3_and ));
    InMux I__3867 (
            .O(N__23382),
            .I(N__23379));
    LocalMux I__3866 (
            .O(N__23379),
            .I(\b2v_inst11.count_off_0_5 ));
    CascadeMux I__3865 (
            .O(N__23376),
            .I(N__23373));
    InMux I__3864 (
            .O(N__23373),
            .I(N__23367));
    InMux I__3863 (
            .O(N__23372),
            .I(N__23367));
    LocalMux I__3862 (
            .O(N__23367),
            .I(N__23364));
    Odrv4 I__3861 (
            .O(N__23364),
            .I(\b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ));
    CascadeMux I__3860 (
            .O(N__23361),
            .I(N__23357));
    InMux I__3859 (
            .O(N__23360),
            .I(N__23354));
    InMux I__3858 (
            .O(N__23357),
            .I(N__23351));
    LocalMux I__3857 (
            .O(N__23354),
            .I(N__23346));
    LocalMux I__3856 (
            .O(N__23351),
            .I(N__23346));
    Odrv4 I__3855 (
            .O(N__23346),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    InMux I__3854 (
            .O(N__23343),
            .I(N__23340));
    LocalMux I__3853 (
            .O(N__23340),
            .I(\b2v_inst11.count_off_0_6 ));
    CascadeMux I__3852 (
            .O(N__23337),
            .I(N__23334));
    InMux I__3851 (
            .O(N__23334),
            .I(N__23330));
    CascadeMux I__3850 (
            .O(N__23333),
            .I(N__23327));
    LocalMux I__3849 (
            .O(N__23330),
            .I(N__23324));
    InMux I__3848 (
            .O(N__23327),
            .I(N__23321));
    Span4Mux_v I__3847 (
            .O(N__23324),
            .I(N__23318));
    LocalMux I__3846 (
            .O(N__23321),
            .I(N__23315));
    Odrv4 I__3845 (
            .O(N__23318),
            .I(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ));
    Odrv4 I__3844 (
            .O(N__23315),
            .I(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ));
    CascadeMux I__3843 (
            .O(N__23310),
            .I(N__23307));
    InMux I__3842 (
            .O(N__23307),
            .I(N__23303));
    InMux I__3841 (
            .O(N__23306),
            .I(N__23300));
    LocalMux I__3840 (
            .O(N__23303),
            .I(N__23297));
    LocalMux I__3839 (
            .O(N__23300),
            .I(N__23294));
    Span4Mux_h I__3838 (
            .O(N__23297),
            .I(N__23291));
    Odrv4 I__3837 (
            .O(N__23294),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    Odrv4 I__3836 (
            .O(N__23291),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    InMux I__3835 (
            .O(N__23286),
            .I(N__23283));
    LocalMux I__3834 (
            .O(N__23283),
            .I(N__23280));
    Odrv4 I__3833 (
            .O(N__23280),
            .I(\b2v_inst20.un4_counter_1_and ));
    InMux I__3832 (
            .O(N__23277),
            .I(N__23274));
    LocalMux I__3831 (
            .O(N__23274),
            .I(N__23271));
    Span4Mux_v I__3830 (
            .O(N__23271),
            .I(N__23268));
    Odrv4 I__3829 (
            .O(N__23268),
            .I(\b2v_inst20.un4_counter_2_and ));
    InMux I__3828 (
            .O(N__23265),
            .I(N__23262));
    LocalMux I__3827 (
            .O(N__23262),
            .I(N__23259));
    Odrv4 I__3826 (
            .O(N__23259),
            .I(\b2v_inst20.counter_1_cry_4_THRU_CO ));
    CascadeMux I__3825 (
            .O(N__23256),
            .I(N__23253));
    InMux I__3824 (
            .O(N__23253),
            .I(N__23250));
    LocalMux I__3823 (
            .O(N__23250),
            .I(N__23245));
    InMux I__3822 (
            .O(N__23249),
            .I(N__23240));
    InMux I__3821 (
            .O(N__23248),
            .I(N__23240));
    Odrv4 I__3820 (
            .O(N__23245),
            .I(\b2v_inst20.counterZ0Z_5 ));
    LocalMux I__3819 (
            .O(N__23240),
            .I(\b2v_inst20.counterZ0Z_5 ));
    InMux I__3818 (
            .O(N__23235),
            .I(N__23232));
    LocalMux I__3817 (
            .O(N__23232),
            .I(N__23229));
    Odrv4 I__3816 (
            .O(N__23229),
            .I(\b2v_inst20.counter_1_cry_5_THRU_CO ));
    InMux I__3815 (
            .O(N__23226),
            .I(N__23222));
    CascadeMux I__3814 (
            .O(N__23225),
            .I(N__23218));
    LocalMux I__3813 (
            .O(N__23222),
            .I(N__23215));
    InMux I__3812 (
            .O(N__23221),
            .I(N__23210));
    InMux I__3811 (
            .O(N__23218),
            .I(N__23210));
    Odrv4 I__3810 (
            .O(N__23215),
            .I(\b2v_inst20.counterZ0Z_6 ));
    LocalMux I__3809 (
            .O(N__23210),
            .I(\b2v_inst20.counterZ0Z_6 ));
    CascadeMux I__3808 (
            .O(N__23205),
            .I(N__23202));
    InMux I__3807 (
            .O(N__23202),
            .I(N__23198));
    CascadeMux I__3806 (
            .O(N__23201),
            .I(N__23195));
    LocalMux I__3805 (
            .O(N__23198),
            .I(N__23192));
    InMux I__3804 (
            .O(N__23195),
            .I(N__23189));
    Span4Mux_v I__3803 (
            .O(N__23192),
            .I(N__23186));
    LocalMux I__3802 (
            .O(N__23189),
            .I(N__23183));
    Odrv4 I__3801 (
            .O(N__23186),
            .I(\b2v_inst11.count_offZ0Z_3 ));
    Odrv4 I__3800 (
            .O(N__23183),
            .I(\b2v_inst11.count_offZ0Z_3 ));
    CascadeMux I__3799 (
            .O(N__23178),
            .I(N__23175));
    InMux I__3798 (
            .O(N__23175),
            .I(N__23172));
    LocalMux I__3797 (
            .O(N__23172),
            .I(N__23169));
    Span4Mux_h I__3796 (
            .O(N__23169),
            .I(N__23164));
    InMux I__3795 (
            .O(N__23168),
            .I(N__23159));
    InMux I__3794 (
            .O(N__23167),
            .I(N__23159));
    Odrv4 I__3793 (
            .O(N__23164),
            .I(\b2v_inst20.counterZ0Z_1 ));
    LocalMux I__3792 (
            .O(N__23159),
            .I(\b2v_inst20.counterZ0Z_1 ));
    InMux I__3791 (
            .O(N__23154),
            .I(N__23134));
    InMux I__3790 (
            .O(N__23153),
            .I(N__23134));
    InMux I__3789 (
            .O(N__23152),
            .I(N__23134));
    InMux I__3788 (
            .O(N__23151),
            .I(N__23134));
    InMux I__3787 (
            .O(N__23150),
            .I(N__23134));
    InMux I__3786 (
            .O(N__23149),
            .I(N__23134));
    CascadeMux I__3785 (
            .O(N__23148),
            .I(N__23131));
    InMux I__3784 (
            .O(N__23147),
            .I(N__23128));
    LocalMux I__3783 (
            .O(N__23134),
            .I(N__23125));
    InMux I__3782 (
            .O(N__23131),
            .I(N__23122));
    LocalMux I__3781 (
            .O(N__23128),
            .I(N__23119));
    Span4Mux_v I__3780 (
            .O(N__23125),
            .I(N__23114));
    LocalMux I__3779 (
            .O(N__23122),
            .I(N__23114));
    Span4Mux_v I__3778 (
            .O(N__23119),
            .I(N__23111));
    Span4Mux_h I__3777 (
            .O(N__23114),
            .I(N__23108));
    Span4Mux_v I__3776 (
            .O(N__23111),
            .I(N__23105));
    Span4Mux_v I__3775 (
            .O(N__23108),
            .I(N__23102));
    Span4Mux_h I__3774 (
            .O(N__23105),
            .I(N__23099));
    Span4Mux_v I__3773 (
            .O(N__23102),
            .I(N__23096));
    Odrv4 I__3772 (
            .O(N__23099),
            .I(v33dsw_ok));
    Odrv4 I__3771 (
            .O(N__23096),
            .I(v33dsw_ok));
    InMux I__3770 (
            .O(N__23091),
            .I(N__23087));
    InMux I__3769 (
            .O(N__23090),
            .I(N__23083));
    LocalMux I__3768 (
            .O(N__23087),
            .I(N__23079));
    CascadeMux I__3767 (
            .O(N__23086),
            .I(N__23076));
    LocalMux I__3766 (
            .O(N__23083),
            .I(N__23073));
    CascadeMux I__3765 (
            .O(N__23082),
            .I(N__23069));
    Span4Mux_h I__3764 (
            .O(N__23079),
            .I(N__23064));
    InMux I__3763 (
            .O(N__23076),
            .I(N__23061));
    Span4Mux_s3_h I__3762 (
            .O(N__23073),
            .I(N__23058));
    InMux I__3761 (
            .O(N__23072),
            .I(N__23049));
    InMux I__3760 (
            .O(N__23069),
            .I(N__23049));
    InMux I__3759 (
            .O(N__23068),
            .I(N__23049));
    InMux I__3758 (
            .O(N__23067),
            .I(N__23049));
    Odrv4 I__3757 (
            .O(N__23064),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    LocalMux I__3756 (
            .O(N__23061),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    Odrv4 I__3755 (
            .O(N__23058),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    LocalMux I__3754 (
            .O(N__23049),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    InMux I__3753 (
            .O(N__23040),
            .I(N__23037));
    LocalMux I__3752 (
            .O(N__23037),
            .I(N__23033));
    InMux I__3751 (
            .O(N__23036),
            .I(N__23030));
    Span4Mux_v I__3750 (
            .O(N__23033),
            .I(N__23026));
    LocalMux I__3749 (
            .O(N__23030),
            .I(N__23023));
    CascadeMux I__3748 (
            .O(N__23029),
            .I(N__23017));
    Span4Mux_h I__3747 (
            .O(N__23026),
            .I(N__23013));
    Span4Mux_s3_h I__3746 (
            .O(N__23023),
            .I(N__23010));
    InMux I__3745 (
            .O(N__23022),
            .I(N__22999));
    InMux I__3744 (
            .O(N__23021),
            .I(N__22999));
    InMux I__3743 (
            .O(N__23020),
            .I(N__22999));
    InMux I__3742 (
            .O(N__23017),
            .I(N__22999));
    InMux I__3741 (
            .O(N__23016),
            .I(N__22999));
    Odrv4 I__3740 (
            .O(N__23013),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    Odrv4 I__3739 (
            .O(N__23010),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    LocalMux I__3738 (
            .O(N__22999),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    CascadeMux I__3737 (
            .O(N__22992),
            .I(N__22989));
    InMux I__3736 (
            .O(N__22989),
            .I(N__22985));
    InMux I__3735 (
            .O(N__22988),
            .I(N__22982));
    LocalMux I__3734 (
            .O(N__22985),
            .I(N__22979));
    LocalMux I__3733 (
            .O(N__22982),
            .I(\b2v_inst11.count_offZ0Z_4 ));
    Odrv4 I__3732 (
            .O(N__22979),
            .I(\b2v_inst11.count_offZ0Z_4 ));
    CascadeMux I__3731 (
            .O(N__22974),
            .I(N__22971));
    InMux I__3730 (
            .O(N__22971),
            .I(N__22965));
    InMux I__3729 (
            .O(N__22970),
            .I(N__22965));
    LocalMux I__3728 (
            .O(N__22965),
            .I(N__22962));
    Span4Mux_v I__3727 (
            .O(N__22962),
            .I(N__22959));
    Odrv4 I__3726 (
            .O(N__22959),
            .I(\b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ));
    InMux I__3725 (
            .O(N__22956),
            .I(N__22953));
    LocalMux I__3724 (
            .O(N__22953),
            .I(\b2v_inst11.count_off_0_4 ));
    InMux I__3723 (
            .O(N__22950),
            .I(N__22946));
    InMux I__3722 (
            .O(N__22949),
            .I(N__22943));
    LocalMux I__3721 (
            .O(N__22946),
            .I(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ));
    LocalMux I__3720 (
            .O(N__22943),
            .I(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ));
    InMux I__3719 (
            .O(N__22938),
            .I(N__22935));
    LocalMux I__3718 (
            .O(N__22935),
            .I(N__22932));
    Odrv12 I__3717 (
            .O(N__22932),
            .I(\b2v_inst11.count_off_0_15 ));
    InMux I__3716 (
            .O(N__22929),
            .I(N__22926));
    LocalMux I__3715 (
            .O(N__22926),
            .I(\b2v_inst11.count_off_0_2 ));
    InMux I__3714 (
            .O(N__22923),
            .I(N__22917));
    InMux I__3713 (
            .O(N__22922),
            .I(N__22917));
    LocalMux I__3712 (
            .O(N__22917),
            .I(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ));
    CascadeMux I__3711 (
            .O(N__22914),
            .I(N__22911));
    InMux I__3710 (
            .O(N__22911),
            .I(N__22908));
    LocalMux I__3709 (
            .O(N__22908),
            .I(\b2v_inst11.count_off_0_0 ));
    InMux I__3708 (
            .O(N__22905),
            .I(N__22902));
    LocalMux I__3707 (
            .O(N__22902),
            .I(N__22896));
    CascadeMux I__3706 (
            .O(N__22901),
            .I(N__22893));
    InMux I__3705 (
            .O(N__22900),
            .I(N__22888));
    InMux I__3704 (
            .O(N__22899),
            .I(N__22888));
    Span4Mux_h I__3703 (
            .O(N__22896),
            .I(N__22885));
    InMux I__3702 (
            .O(N__22893),
            .I(N__22882));
    LocalMux I__3701 (
            .O(N__22888),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    Odrv4 I__3700 (
            .O(N__22885),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    LocalMux I__3699 (
            .O(N__22882),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    CascadeMux I__3698 (
            .O(N__22875),
            .I(\b2v_inst11.count_offZ0Z_0_cascade_ ));
    InMux I__3697 (
            .O(N__22872),
            .I(N__22869));
    LocalMux I__3696 (
            .O(N__22869),
            .I(\b2v_inst11.count_off_RNIZ0Z_1 ));
    InMux I__3695 (
            .O(N__22866),
            .I(N__22863));
    LocalMux I__3694 (
            .O(N__22863),
            .I(\b2v_inst11.count_off_0_1 ));
    CascadeMux I__3693 (
            .O(N__22860),
            .I(\b2v_inst11.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__3692 (
            .O(N__22857),
            .I(N__22853));
    InMux I__3691 (
            .O(N__22856),
            .I(N__22850));
    LocalMux I__3690 (
            .O(N__22853),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    LocalMux I__3689 (
            .O(N__22850),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    CascadeMux I__3688 (
            .O(N__22845),
            .I(\b2v_inst11.count_offZ0Z_1_cascade_ ));
    CascadeMux I__3687 (
            .O(N__22842),
            .I(N__22838));
    InMux I__3686 (
            .O(N__22841),
            .I(N__22835));
    InMux I__3685 (
            .O(N__22838),
            .I(N__22832));
    LocalMux I__3684 (
            .O(N__22835),
            .I(\b2v_inst11.count_offZ0Z_2 ));
    LocalMux I__3683 (
            .O(N__22832),
            .I(\b2v_inst11.count_offZ0Z_2 ));
    InMux I__3682 (
            .O(N__22827),
            .I(N__22823));
    InMux I__3681 (
            .O(N__22826),
            .I(N__22820));
    LocalMux I__3680 (
            .O(N__22823),
            .I(N__22817));
    LocalMux I__3679 (
            .O(N__22820),
            .I(\b2v_inst20.counterZ0Z_7 ));
    Odrv4 I__3678 (
            .O(N__22817),
            .I(\b2v_inst20.counterZ0Z_7 ));
    InMux I__3677 (
            .O(N__22812),
            .I(\b2v_inst5.un2_count_1_cry_14 ));
    CascadeMux I__3676 (
            .O(N__22809),
            .I(\b2v_inst5.countZ0Z_4_cascade_ ));
    InMux I__3675 (
            .O(N__22806),
            .I(N__22803));
    LocalMux I__3674 (
            .O(N__22803),
            .I(\b2v_inst5.count_rst_6 ));
    CascadeMux I__3673 (
            .O(N__22800),
            .I(\b2v_inst5.count_rst_6_cascade_ ));
    CascadeMux I__3672 (
            .O(N__22797),
            .I(N__22793));
    CascadeMux I__3671 (
            .O(N__22796),
            .I(N__22790));
    InMux I__3670 (
            .O(N__22793),
            .I(N__22787));
    InMux I__3669 (
            .O(N__22790),
            .I(N__22784));
    LocalMux I__3668 (
            .O(N__22787),
            .I(\b2v_inst5.un2_count_1_axb_8 ));
    LocalMux I__3667 (
            .O(N__22784),
            .I(\b2v_inst5.un2_count_1_axb_8 ));
    InMux I__3666 (
            .O(N__22779),
            .I(N__22773));
    InMux I__3665 (
            .O(N__22778),
            .I(N__22773));
    LocalMux I__3664 (
            .O(N__22773),
            .I(\b2v_inst5.un2_count_1_cry_7_THRU_CO ));
    CascadeMux I__3663 (
            .O(N__22770),
            .I(\b2v_inst5.un2_count_1_axb_8_cascade_ ));
    InMux I__3662 (
            .O(N__22767),
            .I(N__22761));
    InMux I__3661 (
            .O(N__22766),
            .I(N__22761));
    LocalMux I__3660 (
            .O(N__22761),
            .I(\b2v_inst5.count_1_8 ));
    InMux I__3659 (
            .O(N__22758),
            .I(N__22755));
    LocalMux I__3658 (
            .O(N__22755),
            .I(\b2v_inst5.count_rst_10 ));
    InMux I__3657 (
            .O(N__22752),
            .I(N__22746));
    InMux I__3656 (
            .O(N__22751),
            .I(N__22746));
    LocalMux I__3655 (
            .O(N__22746),
            .I(N__22743));
    Odrv4 I__3654 (
            .O(N__22743),
            .I(\b2v_inst5.un2_count_1_cry_3_THRU_CO ));
    CascadeMux I__3653 (
            .O(N__22740),
            .I(N__22736));
    InMux I__3652 (
            .O(N__22739),
            .I(N__22732));
    InMux I__3651 (
            .O(N__22736),
            .I(N__22727));
    InMux I__3650 (
            .O(N__22735),
            .I(N__22727));
    LocalMux I__3649 (
            .O(N__22732),
            .I(N__22724));
    LocalMux I__3648 (
            .O(N__22727),
            .I(\b2v_inst5.countZ0Z_4 ));
    Odrv4 I__3647 (
            .O(N__22724),
            .I(\b2v_inst5.countZ0Z_4 ));
    InMux I__3646 (
            .O(N__22719),
            .I(N__22716));
    LocalMux I__3645 (
            .O(N__22716),
            .I(\b2v_inst5.count_1_4 ));
    InMux I__3644 (
            .O(N__22713),
            .I(\b2v_inst5.un2_count_1_cry_5 ));
    InMux I__3643 (
            .O(N__22710),
            .I(\b2v_inst5.un2_count_1_cry_6 ));
    InMux I__3642 (
            .O(N__22707),
            .I(bfn_6_4_0_));
    InMux I__3641 (
            .O(N__22704),
            .I(\b2v_inst5.un2_count_1_cry_8 ));
    InMux I__3640 (
            .O(N__22701),
            .I(\b2v_inst5.un2_count_1_cry_9 ));
    InMux I__3639 (
            .O(N__22698),
            .I(\b2v_inst5.un2_count_1_cry_10 ));
    InMux I__3638 (
            .O(N__22695),
            .I(\b2v_inst5.un2_count_1_cry_11 ));
    InMux I__3637 (
            .O(N__22692),
            .I(\b2v_inst5.un2_count_1_cry_12 ));
    InMux I__3636 (
            .O(N__22689),
            .I(\b2v_inst5.un2_count_1_cry_13 ));
    InMux I__3635 (
            .O(N__22686),
            .I(N__22682));
    InMux I__3634 (
            .O(N__22685),
            .I(N__22679));
    LocalMux I__3633 (
            .O(N__22682),
            .I(\b2v_inst200.count_1_6 ));
    LocalMux I__3632 (
            .O(N__22679),
            .I(\b2v_inst200.count_1_6 ));
    InMux I__3631 (
            .O(N__22674),
            .I(N__22671));
    LocalMux I__3630 (
            .O(N__22671),
            .I(\b2v_inst200.count_3_6 ));
    InMux I__3629 (
            .O(N__22668),
            .I(N__22664));
    InMux I__3628 (
            .O(N__22667),
            .I(N__22661));
    LocalMux I__3627 (
            .O(N__22664),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    LocalMux I__3626 (
            .O(N__22661),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    InMux I__3625 (
            .O(N__22656),
            .I(N__22653));
    LocalMux I__3624 (
            .O(N__22653),
            .I(\b2v_inst200.count_3_7 ));
    InMux I__3623 (
            .O(N__22650),
            .I(N__22646));
    InMux I__3622 (
            .O(N__22649),
            .I(N__22643));
    LocalMux I__3621 (
            .O(N__22646),
            .I(N__22640));
    LocalMux I__3620 (
            .O(N__22643),
            .I(\b2v_inst200.count_1_10 ));
    Odrv4 I__3619 (
            .O(N__22640),
            .I(\b2v_inst200.count_1_10 ));
    CascadeMux I__3618 (
            .O(N__22635),
            .I(N__22632));
    InMux I__3617 (
            .O(N__22632),
            .I(N__22629));
    LocalMux I__3616 (
            .O(N__22629),
            .I(\b2v_inst200.count_3_10 ));
    InMux I__3615 (
            .O(N__22626),
            .I(N__22590));
    InMux I__3614 (
            .O(N__22625),
            .I(N__22590));
    InMux I__3613 (
            .O(N__22624),
            .I(N__22590));
    InMux I__3612 (
            .O(N__22623),
            .I(N__22590));
    InMux I__3611 (
            .O(N__22622),
            .I(N__22590));
    InMux I__3610 (
            .O(N__22621),
            .I(N__22579));
    InMux I__3609 (
            .O(N__22620),
            .I(N__22579));
    InMux I__3608 (
            .O(N__22619),
            .I(N__22579));
    InMux I__3607 (
            .O(N__22618),
            .I(N__22579));
    InMux I__3606 (
            .O(N__22617),
            .I(N__22579));
    InMux I__3605 (
            .O(N__22616),
            .I(N__22574));
    InMux I__3604 (
            .O(N__22615),
            .I(N__22574));
    InMux I__3603 (
            .O(N__22614),
            .I(N__22565));
    InMux I__3602 (
            .O(N__22613),
            .I(N__22565));
    InMux I__3601 (
            .O(N__22612),
            .I(N__22565));
    InMux I__3600 (
            .O(N__22611),
            .I(N__22565));
    InMux I__3599 (
            .O(N__22610),
            .I(N__22552));
    InMux I__3598 (
            .O(N__22609),
            .I(N__22552));
    InMux I__3597 (
            .O(N__22608),
            .I(N__22552));
    InMux I__3596 (
            .O(N__22607),
            .I(N__22552));
    InMux I__3595 (
            .O(N__22606),
            .I(N__22552));
    InMux I__3594 (
            .O(N__22605),
            .I(N__22552));
    InMux I__3593 (
            .O(N__22604),
            .I(N__22543));
    InMux I__3592 (
            .O(N__22603),
            .I(N__22543));
    InMux I__3591 (
            .O(N__22602),
            .I(N__22543));
    InMux I__3590 (
            .O(N__22601),
            .I(N__22543));
    LocalMux I__3589 (
            .O(N__22590),
            .I(N__22534));
    LocalMux I__3588 (
            .O(N__22579),
            .I(N__22531));
    LocalMux I__3587 (
            .O(N__22574),
            .I(N__22528));
    LocalMux I__3586 (
            .O(N__22565),
            .I(N__22525));
    LocalMux I__3585 (
            .O(N__22552),
            .I(N__22522));
    LocalMux I__3584 (
            .O(N__22543),
            .I(N__22519));
    CEMux I__3583 (
            .O(N__22542),
            .I(N__22494));
    CEMux I__3582 (
            .O(N__22541),
            .I(N__22494));
    CEMux I__3581 (
            .O(N__22540),
            .I(N__22494));
    CEMux I__3580 (
            .O(N__22539),
            .I(N__22494));
    CEMux I__3579 (
            .O(N__22538),
            .I(N__22494));
    CEMux I__3578 (
            .O(N__22537),
            .I(N__22494));
    Glb2LocalMux I__3577 (
            .O(N__22534),
            .I(N__22494));
    Glb2LocalMux I__3576 (
            .O(N__22531),
            .I(N__22494));
    Glb2LocalMux I__3575 (
            .O(N__22528),
            .I(N__22494));
    Glb2LocalMux I__3574 (
            .O(N__22525),
            .I(N__22494));
    Glb2LocalMux I__3573 (
            .O(N__22522),
            .I(N__22494));
    Glb2LocalMux I__3572 (
            .O(N__22519),
            .I(N__22494));
    GlobalMux I__3571 (
            .O(N__22494),
            .I(N__22491));
    gio2CtrlBuf I__3570 (
            .O(N__22491),
            .I(\b2v_inst200.count_en_g ));
    InMux I__3569 (
            .O(N__22488),
            .I(\b2v_inst5.un2_count_1_cry_0 ));
    InMux I__3568 (
            .O(N__22485),
            .I(\b2v_inst5.un2_count_1_cry_1 ));
    InMux I__3567 (
            .O(N__22482),
            .I(\b2v_inst5.un2_count_1_cry_2 ));
    InMux I__3566 (
            .O(N__22479),
            .I(\b2v_inst5.un2_count_1_cry_3 ));
    InMux I__3565 (
            .O(N__22476),
            .I(\b2v_inst5.un2_count_1_cry_4 ));
    InMux I__3564 (
            .O(N__22473),
            .I(N__22467));
    InMux I__3563 (
            .O(N__22472),
            .I(N__22467));
    LocalMux I__3562 (
            .O(N__22467),
            .I(\b2v_inst200.count_3_15 ));
    CascadeMux I__3561 (
            .O(N__22464),
            .I(N__22461));
    InMux I__3560 (
            .O(N__22461),
            .I(N__22458));
    LocalMux I__3559 (
            .O(N__22458),
            .I(N__22454));
    InMux I__3558 (
            .O(N__22457),
            .I(N__22451));
    Odrv4 I__3557 (
            .O(N__22454),
            .I(\b2v_inst200.countZ0Z_6 ));
    LocalMux I__3556 (
            .O(N__22451),
            .I(\b2v_inst200.countZ0Z_6 ));
    InMux I__3555 (
            .O(N__22446),
            .I(N__22437));
    InMux I__3554 (
            .O(N__22445),
            .I(N__22437));
    InMux I__3553 (
            .O(N__22444),
            .I(N__22437));
    LocalMux I__3552 (
            .O(N__22437),
            .I(N__22434));
    Odrv4 I__3551 (
            .O(N__22434),
            .I(\b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71 ));
    InMux I__3550 (
            .O(N__22431),
            .I(N__22426));
    InMux I__3549 (
            .O(N__22430),
            .I(N__22421));
    InMux I__3548 (
            .O(N__22429),
            .I(N__22421));
    LocalMux I__3547 (
            .O(N__22426),
            .I(\b2v_inst200.count_1_8 ));
    LocalMux I__3546 (
            .O(N__22421),
            .I(\b2v_inst200.count_1_8 ));
    InMux I__3545 (
            .O(N__22416),
            .I(N__22412));
    InMux I__3544 (
            .O(N__22415),
            .I(N__22409));
    LocalMux I__3543 (
            .O(N__22412),
            .I(\b2v_inst200.count_3_8 ));
    LocalMux I__3542 (
            .O(N__22409),
            .I(\b2v_inst200.count_3_8 ));
    CascadeMux I__3541 (
            .O(N__22404),
            .I(N__22400));
    InMux I__3540 (
            .O(N__22403),
            .I(N__22397));
    InMux I__3539 (
            .O(N__22400),
            .I(N__22394));
    LocalMux I__3538 (
            .O(N__22397),
            .I(N__22391));
    LocalMux I__3537 (
            .O(N__22394),
            .I(\b2v_inst200.countZ0Z_10 ));
    Odrv4 I__3536 (
            .O(N__22391),
            .I(\b2v_inst200.countZ0Z_10 ));
    InMux I__3535 (
            .O(N__22386),
            .I(N__22383));
    LocalMux I__3534 (
            .O(N__22383),
            .I(N__22380));
    Span4Mux_h I__3533 (
            .O(N__22380),
            .I(N__22377));
    Odrv4 I__3532 (
            .O(N__22377),
            .I(\b2v_inst200.un25_clk_100khz_14 ));
    InMux I__3531 (
            .O(N__22374),
            .I(N__22371));
    LocalMux I__3530 (
            .O(N__22371),
            .I(\b2v_inst200.un25_clk_100khz_6 ));
    CascadeMux I__3529 (
            .O(N__22368),
            .I(\b2v_inst200.un25_clk_100khz_7_cascade_ ));
    InMux I__3528 (
            .O(N__22365),
            .I(N__22362));
    LocalMux I__3527 (
            .O(N__22362),
            .I(N__22359));
    Odrv4 I__3526 (
            .O(N__22359),
            .I(\b2v_inst200.un25_clk_100khz_13 ));
    InMux I__3525 (
            .O(N__22356),
            .I(N__22351));
    InMux I__3524 (
            .O(N__22355),
            .I(N__22348));
    InMux I__3523 (
            .O(N__22354),
            .I(N__22345));
    LocalMux I__3522 (
            .O(N__22351),
            .I(N__22336));
    LocalMux I__3521 (
            .O(N__22348),
            .I(N__22333));
    LocalMux I__3520 (
            .O(N__22345),
            .I(N__22330));
    InMux I__3519 (
            .O(N__22344),
            .I(N__22325));
    InMux I__3518 (
            .O(N__22343),
            .I(N__22325));
    InMux I__3517 (
            .O(N__22342),
            .I(N__22320));
    InMux I__3516 (
            .O(N__22341),
            .I(N__22320));
    InMux I__3515 (
            .O(N__22340),
            .I(N__22315));
    InMux I__3514 (
            .O(N__22339),
            .I(N__22315));
    Span4Mux_v I__3513 (
            .O(N__22336),
            .I(N__22309));
    Span4Mux_h I__3512 (
            .O(N__22333),
            .I(N__22309));
    Span4Mux_v I__3511 (
            .O(N__22330),
            .I(N__22300));
    LocalMux I__3510 (
            .O(N__22325),
            .I(N__22300));
    LocalMux I__3509 (
            .O(N__22320),
            .I(N__22300));
    LocalMux I__3508 (
            .O(N__22315),
            .I(N__22300));
    InMux I__3507 (
            .O(N__22314),
            .I(N__22297));
    Odrv4 I__3506 (
            .O(N__22309),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    Odrv4 I__3505 (
            .O(N__22300),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    LocalMux I__3504 (
            .O(N__22297),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8 ));
    CascadeMux I__3503 (
            .O(N__22290),
            .I(\b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_ ));
    InMux I__3502 (
            .O(N__22287),
            .I(N__22279));
    InMux I__3501 (
            .O(N__22286),
            .I(N__22276));
    InMux I__3500 (
            .O(N__22285),
            .I(N__22273));
    InMux I__3499 (
            .O(N__22284),
            .I(N__22266));
    InMux I__3498 (
            .O(N__22283),
            .I(N__22266));
    InMux I__3497 (
            .O(N__22282),
            .I(N__22266));
    LocalMux I__3496 (
            .O(N__22279),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__3495 (
            .O(N__22276),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__3494 (
            .O(N__22273),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__3493 (
            .O(N__22266),
            .I(\b2v_inst200.countZ0Z_0 ));
    InMux I__3492 (
            .O(N__22257),
            .I(N__22254));
    LocalMux I__3491 (
            .O(N__22254),
            .I(\b2v_inst200.count_3_0 ));
    InMux I__3490 (
            .O(N__22251),
            .I(N__22247));
    InMux I__3489 (
            .O(N__22250),
            .I(N__22244));
    LocalMux I__3488 (
            .O(N__22247),
            .I(\b2v_inst200.count_1_11 ));
    LocalMux I__3487 (
            .O(N__22244),
            .I(\b2v_inst200.count_1_11 ));
    InMux I__3486 (
            .O(N__22239),
            .I(N__22236));
    LocalMux I__3485 (
            .O(N__22236),
            .I(N__22233));
    Span4Mux_h I__3484 (
            .O(N__22233),
            .I(N__22230));
    Odrv4 I__3483 (
            .O(N__22230),
            .I(\b2v_inst200.count_3_11 ));
    InMux I__3482 (
            .O(N__22227),
            .I(N__22223));
    InMux I__3481 (
            .O(N__22226),
            .I(N__22220));
    LocalMux I__3480 (
            .O(N__22223),
            .I(N__22217));
    LocalMux I__3479 (
            .O(N__22220),
            .I(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ));
    Odrv4 I__3478 (
            .O(N__22217),
            .I(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ));
    InMux I__3477 (
            .O(N__22212),
            .I(N__22209));
    LocalMux I__3476 (
            .O(N__22209),
            .I(\b2v_inst200.count_3_14 ));
    InMux I__3475 (
            .O(N__22206),
            .I(N__22202));
    InMux I__3474 (
            .O(N__22205),
            .I(N__22199));
    LocalMux I__3473 (
            .O(N__22202),
            .I(N__22196));
    LocalMux I__3472 (
            .O(N__22199),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    Odrv4 I__3471 (
            .O(N__22196),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    InMux I__3470 (
            .O(N__22191),
            .I(N__22188));
    LocalMux I__3469 (
            .O(N__22188),
            .I(N__22185));
    Span4Mux_v I__3468 (
            .O(N__22185),
            .I(N__22182));
    Odrv4 I__3467 (
            .O(N__22182),
            .I(\b2v_inst200.count_3_2 ));
    InMux I__3466 (
            .O(N__22179),
            .I(N__22175));
    InMux I__3465 (
            .O(N__22178),
            .I(N__22172));
    LocalMux I__3464 (
            .O(N__22175),
            .I(N__22169));
    LocalMux I__3463 (
            .O(N__22172),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    Odrv4 I__3462 (
            .O(N__22169),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    InMux I__3461 (
            .O(N__22164),
            .I(N__22161));
    LocalMux I__3460 (
            .O(N__22161),
            .I(N__22158));
    Span4Mux_v I__3459 (
            .O(N__22158),
            .I(N__22155));
    Odrv4 I__3458 (
            .O(N__22155),
            .I(\b2v_inst200.count_3_4 ));
    InMux I__3457 (
            .O(N__22152),
            .I(N__22149));
    LocalMux I__3456 (
            .O(N__22149),
            .I(\b2v_inst11.mult1_un89_sum_cry_5_s ));
    InMux I__3455 (
            .O(N__22146),
            .I(N__22143));
    LocalMux I__3454 (
            .O(N__22143),
            .I(N__22140));
    Odrv4 I__3453 (
            .O(N__22140),
            .I(\b2v_inst11.mult1_un96_sum_cry_6_s ));
    InMux I__3452 (
            .O(N__22137),
            .I(\b2v_inst11.mult1_un96_sum_cry_5 ));
    InMux I__3451 (
            .O(N__22134),
            .I(N__22131));
    LocalMux I__3450 (
            .O(N__22131),
            .I(\b2v_inst11.mult1_un89_sum_cry_6_s ));
    CascadeMux I__3449 (
            .O(N__22128),
            .I(N__22125));
    InMux I__3448 (
            .O(N__22125),
            .I(N__22122));
    LocalMux I__3447 (
            .O(N__22122),
            .I(N__22119));
    Odrv4 I__3446 (
            .O(N__22119),
            .I(\b2v_inst11.mult1_un103_sum_axb_8 ));
    InMux I__3445 (
            .O(N__22116),
            .I(\b2v_inst11.mult1_un96_sum_cry_6 ));
    CascadeMux I__3444 (
            .O(N__22113),
            .I(N__22110));
    InMux I__3443 (
            .O(N__22110),
            .I(N__22107));
    LocalMux I__3442 (
            .O(N__22107),
            .I(\b2v_inst11.mult1_un96_sum_axb_8 ));
    InMux I__3441 (
            .O(N__22104),
            .I(\b2v_inst11.mult1_un96_sum_cry_7 ));
    InMux I__3440 (
            .O(N__22101),
            .I(N__22097));
    CascadeMux I__3439 (
            .O(N__22100),
            .I(N__22094));
    LocalMux I__3438 (
            .O(N__22097),
            .I(N__22088));
    InMux I__3437 (
            .O(N__22094),
            .I(N__22081));
    InMux I__3436 (
            .O(N__22093),
            .I(N__22081));
    InMux I__3435 (
            .O(N__22092),
            .I(N__22081));
    InMux I__3434 (
            .O(N__22091),
            .I(N__22078));
    Span4Mux_v I__3433 (
            .O(N__22088),
            .I(N__22073));
    LocalMux I__3432 (
            .O(N__22081),
            .I(N__22073));
    LocalMux I__3431 (
            .O(N__22078),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    Odrv4 I__3430 (
            .O(N__22073),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    InMux I__3429 (
            .O(N__22068),
            .I(N__22064));
    CascadeMux I__3428 (
            .O(N__22067),
            .I(N__22060));
    LocalMux I__3427 (
            .O(N__22064),
            .I(N__22055));
    InMux I__3426 (
            .O(N__22063),
            .I(N__22052));
    InMux I__3425 (
            .O(N__22060),
            .I(N__22045));
    InMux I__3424 (
            .O(N__22059),
            .I(N__22045));
    InMux I__3423 (
            .O(N__22058),
            .I(N__22045));
    Odrv4 I__3422 (
            .O(N__22055),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__3421 (
            .O(N__22052),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__3420 (
            .O(N__22045),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    CascadeMux I__3419 (
            .O(N__22038),
            .I(N__22034));
    CascadeMux I__3418 (
            .O(N__22037),
            .I(N__22030));
    InMux I__3417 (
            .O(N__22034),
            .I(N__22023));
    InMux I__3416 (
            .O(N__22033),
            .I(N__22023));
    InMux I__3415 (
            .O(N__22030),
            .I(N__22023));
    LocalMux I__3414 (
            .O(N__22023),
            .I(\b2v_inst11.mult1_un89_sum_i_0_8 ));
    CascadeMux I__3413 (
            .O(N__22020),
            .I(N__22017));
    InMux I__3412 (
            .O(N__22017),
            .I(N__22014));
    LocalMux I__3411 (
            .O(N__22014),
            .I(N__22011));
    Odrv4 I__3410 (
            .O(N__22011),
            .I(\b2v_inst200.un2_count_1_axb_15 ));
    InMux I__3409 (
            .O(N__22008),
            .I(N__22005));
    LocalMux I__3408 (
            .O(N__22005),
            .I(\b2v_inst200.un2_count_1_axb_8 ));
    InMux I__3407 (
            .O(N__22002),
            .I(\b2v_inst11.mult1_un89_sum_cry_4 ));
    InMux I__3406 (
            .O(N__21999),
            .I(\b2v_inst11.mult1_un89_sum_cry_5 ));
    InMux I__3405 (
            .O(N__21996),
            .I(\b2v_inst11.mult1_un89_sum_cry_6 ));
    InMux I__3404 (
            .O(N__21993),
            .I(\b2v_inst11.mult1_un89_sum_cry_7 ));
    CascadeMux I__3403 (
            .O(N__21990),
            .I(N__21986));
    CascadeMux I__3402 (
            .O(N__21989),
            .I(N__21982));
    InMux I__3401 (
            .O(N__21986),
            .I(N__21975));
    InMux I__3400 (
            .O(N__21985),
            .I(N__21975));
    InMux I__3399 (
            .O(N__21982),
            .I(N__21975));
    LocalMux I__3398 (
            .O(N__21975),
            .I(\b2v_inst11.mult1_un82_sum_i_0_8 ));
    CascadeMux I__3397 (
            .O(N__21972),
            .I(N__21969));
    InMux I__3396 (
            .O(N__21969),
            .I(N__21966));
    LocalMux I__3395 (
            .O(N__21966),
            .I(N__21963));
    Span4Mux_s2_h I__3394 (
            .O(N__21963),
            .I(N__21960));
    Odrv4 I__3393 (
            .O(N__21960),
            .I(\b2v_inst11.mult1_un96_sum_cry_3_s ));
    InMux I__3392 (
            .O(N__21957),
            .I(\b2v_inst11.mult1_un96_sum_cry_2 ));
    CascadeMux I__3391 (
            .O(N__21954),
            .I(N__21951));
    InMux I__3390 (
            .O(N__21951),
            .I(N__21948));
    LocalMux I__3389 (
            .O(N__21948),
            .I(\b2v_inst11.mult1_un89_sum_cry_3_s ));
    CascadeMux I__3388 (
            .O(N__21945),
            .I(N__21942));
    InMux I__3387 (
            .O(N__21942),
            .I(N__21939));
    LocalMux I__3386 (
            .O(N__21939),
            .I(N__21936));
    Odrv4 I__3385 (
            .O(N__21936),
            .I(\b2v_inst11.mult1_un96_sum_cry_4_s ));
    InMux I__3384 (
            .O(N__21933),
            .I(\b2v_inst11.mult1_un96_sum_cry_3 ));
    CascadeMux I__3383 (
            .O(N__21930),
            .I(N__21927));
    InMux I__3382 (
            .O(N__21927),
            .I(N__21924));
    LocalMux I__3381 (
            .O(N__21924),
            .I(\b2v_inst11.mult1_un89_sum_cry_4_s ));
    InMux I__3380 (
            .O(N__21921),
            .I(N__21918));
    LocalMux I__3379 (
            .O(N__21918),
            .I(N__21915));
    Odrv4 I__3378 (
            .O(N__21915),
            .I(\b2v_inst11.mult1_un96_sum_cry_5_s ));
    InMux I__3377 (
            .O(N__21912),
            .I(\b2v_inst11.mult1_un96_sum_cry_4 ));
    InMux I__3376 (
            .O(N__21909),
            .I(N__21906));
    LocalMux I__3375 (
            .O(N__21906),
            .I(N__21903));
    Span4Mux_v I__3374 (
            .O(N__21903),
            .I(N__21900));
    Odrv4 I__3373 (
            .O(N__21900),
            .I(\b2v_inst11.mult1_un103_sum_cry_4_s ));
    CascadeMux I__3372 (
            .O(N__21897),
            .I(N__21894));
    InMux I__3371 (
            .O(N__21894),
            .I(N__21891));
    LocalMux I__3370 (
            .O(N__21891),
            .I(\b2v_inst11.mult1_un110_sum_cry_5_s ));
    InMux I__3369 (
            .O(N__21888),
            .I(\b2v_inst11.mult1_un110_sum_cry_4 ));
    CascadeMux I__3368 (
            .O(N__21885),
            .I(N__21881));
    InMux I__3367 (
            .O(N__21884),
            .I(N__21876));
    InMux I__3366 (
            .O(N__21881),
            .I(N__21876));
    LocalMux I__3365 (
            .O(N__21876),
            .I(N__21872));
    InMux I__3364 (
            .O(N__21875),
            .I(N__21869));
    Span4Mux_s3_v I__3363 (
            .O(N__21872),
            .I(N__21862));
    LocalMux I__3362 (
            .O(N__21869),
            .I(N__21862));
    InMux I__3361 (
            .O(N__21868),
            .I(N__21859));
    InMux I__3360 (
            .O(N__21867),
            .I(N__21856));
    Span4Mux_h I__3359 (
            .O(N__21862),
            .I(N__21853));
    LocalMux I__3358 (
            .O(N__21859),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    LocalMux I__3357 (
            .O(N__21856),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    Odrv4 I__3356 (
            .O(N__21853),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    CascadeMux I__3355 (
            .O(N__21846),
            .I(N__21843));
    InMux I__3354 (
            .O(N__21843),
            .I(N__21840));
    LocalMux I__3353 (
            .O(N__21840),
            .I(N__21837));
    Span4Mux_v I__3352 (
            .O(N__21837),
            .I(N__21834));
    Odrv4 I__3351 (
            .O(N__21834),
            .I(\b2v_inst11.mult1_un103_sum_cry_5_s ));
    InMux I__3350 (
            .O(N__21831),
            .I(N__21828));
    LocalMux I__3349 (
            .O(N__21828),
            .I(\b2v_inst11.mult1_un110_sum_cry_6_s ));
    InMux I__3348 (
            .O(N__21825),
            .I(\b2v_inst11.mult1_un110_sum_cry_5 ));
    InMux I__3347 (
            .O(N__21822),
            .I(N__21819));
    LocalMux I__3346 (
            .O(N__21819),
            .I(N__21816));
    Span4Mux_h I__3345 (
            .O(N__21816),
            .I(N__21813));
    Odrv4 I__3344 (
            .O(N__21813),
            .I(\b2v_inst11.mult1_un103_sum_cry_6_s ));
    CascadeMux I__3343 (
            .O(N__21810),
            .I(N__21806));
    CascadeMux I__3342 (
            .O(N__21809),
            .I(N__21802));
    InMux I__3341 (
            .O(N__21806),
            .I(N__21795));
    InMux I__3340 (
            .O(N__21805),
            .I(N__21795));
    InMux I__3339 (
            .O(N__21802),
            .I(N__21795));
    LocalMux I__3338 (
            .O(N__21795),
            .I(\b2v_inst11.mult1_un103_sum_i_0_8 ));
    CascadeMux I__3337 (
            .O(N__21792),
            .I(N__21789));
    InMux I__3336 (
            .O(N__21789),
            .I(N__21786));
    LocalMux I__3335 (
            .O(N__21786),
            .I(\b2v_inst11.mult1_un117_sum_axb_8 ));
    InMux I__3334 (
            .O(N__21783),
            .I(\b2v_inst11.mult1_un110_sum_cry_6 ));
    CascadeMux I__3333 (
            .O(N__21780),
            .I(N__21777));
    InMux I__3332 (
            .O(N__21777),
            .I(N__21774));
    LocalMux I__3331 (
            .O(N__21774),
            .I(N__21771));
    Span4Mux_h I__3330 (
            .O(N__21771),
            .I(N__21768));
    Odrv4 I__3329 (
            .O(N__21768),
            .I(\b2v_inst11.mult1_un110_sum_axb_8 ));
    InMux I__3328 (
            .O(N__21765),
            .I(\b2v_inst11.mult1_un110_sum_cry_7 ));
    InMux I__3327 (
            .O(N__21762),
            .I(N__21758));
    CascadeMux I__3326 (
            .O(N__21761),
            .I(N__21754));
    LocalMux I__3325 (
            .O(N__21758),
            .I(N__21750));
    InMux I__3324 (
            .O(N__21757),
            .I(N__21745));
    InMux I__3323 (
            .O(N__21754),
            .I(N__21745));
    InMux I__3322 (
            .O(N__21753),
            .I(N__21742));
    Odrv4 I__3321 (
            .O(N__21750),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__3320 (
            .O(N__21745),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__3319 (
            .O(N__21742),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    CascadeMux I__3318 (
            .O(N__21735),
            .I(\b2v_inst11.mult1_un110_sum_s_8_cascade_ ));
    CascadeMux I__3317 (
            .O(N__21732),
            .I(N__21728));
    CascadeMux I__3316 (
            .O(N__21731),
            .I(N__21724));
    InMux I__3315 (
            .O(N__21728),
            .I(N__21717));
    InMux I__3314 (
            .O(N__21727),
            .I(N__21717));
    InMux I__3313 (
            .O(N__21724),
            .I(N__21717));
    LocalMux I__3312 (
            .O(N__21717),
            .I(\b2v_inst11.mult1_un110_sum_i_0_8 ));
    InMux I__3311 (
            .O(N__21714),
            .I(\b2v_inst11.mult1_un89_sum_cry_2 ));
    InMux I__3310 (
            .O(N__21711),
            .I(\b2v_inst11.mult1_un89_sum_cry_3 ));
    InMux I__3309 (
            .O(N__21708),
            .I(N__21705));
    LocalMux I__3308 (
            .O(N__21705),
            .I(\b2v_inst11.mult1_un138_sum_i ));
    InMux I__3307 (
            .O(N__21702),
            .I(N__21699));
    LocalMux I__3306 (
            .O(N__21699),
            .I(N__21696));
    Span4Mux_s1_v I__3305 (
            .O(N__21696),
            .I(N__21693));
    Odrv4 I__3304 (
            .O(N__21693),
            .I(\b2v_inst11.mult1_un124_sum_i ));
    InMux I__3303 (
            .O(N__21690),
            .I(N__21687));
    LocalMux I__3302 (
            .O(N__21687),
            .I(\b2v_inst11.mult1_un110_sum_i ));
    InMux I__3301 (
            .O(N__21684),
            .I(N__21681));
    LocalMux I__3300 (
            .O(N__21681),
            .I(\b2v_inst11.mult1_un103_sum_i ));
    CascadeMux I__3299 (
            .O(N__21678),
            .I(N__21675));
    InMux I__3298 (
            .O(N__21675),
            .I(N__21672));
    LocalMux I__3297 (
            .O(N__21672),
            .I(\b2v_inst11.mult1_un110_sum_cry_3_s ));
    InMux I__3296 (
            .O(N__21669),
            .I(\b2v_inst11.mult1_un110_sum_cry_2 ));
    CascadeMux I__3295 (
            .O(N__21666),
            .I(N__21663));
    InMux I__3294 (
            .O(N__21663),
            .I(N__21660));
    LocalMux I__3293 (
            .O(N__21660),
            .I(N__21657));
    Span4Mux_h I__3292 (
            .O(N__21657),
            .I(N__21654));
    Odrv4 I__3291 (
            .O(N__21654),
            .I(\b2v_inst11.mult1_un103_sum_cry_3_s ));
    InMux I__3290 (
            .O(N__21651),
            .I(N__21648));
    LocalMux I__3289 (
            .O(N__21648),
            .I(\b2v_inst11.mult1_un110_sum_cry_4_s ));
    InMux I__3288 (
            .O(N__21645),
            .I(\b2v_inst11.mult1_un110_sum_cry_3 ));
    InMux I__3287 (
            .O(N__21642),
            .I(bfn_5_12_0_));
    InMux I__3286 (
            .O(N__21639),
            .I(\b2v_inst20.counter_1_cry_25 ));
    InMux I__3285 (
            .O(N__21636),
            .I(\b2v_inst20.counter_1_cry_26 ));
    InMux I__3284 (
            .O(N__21633),
            .I(N__21629));
    InMux I__3283 (
            .O(N__21632),
            .I(N__21626));
    LocalMux I__3282 (
            .O(N__21629),
            .I(N__21623));
    LocalMux I__3281 (
            .O(N__21626),
            .I(\b2v_inst20.counterZ0Z_28 ));
    Odrv12 I__3280 (
            .O(N__21623),
            .I(\b2v_inst20.counterZ0Z_28 ));
    InMux I__3279 (
            .O(N__21618),
            .I(\b2v_inst20.counter_1_cry_27 ));
    InMux I__3278 (
            .O(N__21615),
            .I(N__21611));
    InMux I__3277 (
            .O(N__21614),
            .I(N__21608));
    LocalMux I__3276 (
            .O(N__21611),
            .I(N__21605));
    LocalMux I__3275 (
            .O(N__21608),
            .I(\b2v_inst20.counterZ0Z_29 ));
    Odrv12 I__3274 (
            .O(N__21605),
            .I(\b2v_inst20.counterZ0Z_29 ));
    InMux I__3273 (
            .O(N__21600),
            .I(\b2v_inst20.counter_1_cry_28 ));
    CascadeMux I__3272 (
            .O(N__21597),
            .I(N__21594));
    InMux I__3271 (
            .O(N__21594),
            .I(N__21590));
    InMux I__3270 (
            .O(N__21593),
            .I(N__21587));
    LocalMux I__3269 (
            .O(N__21590),
            .I(N__21584));
    LocalMux I__3268 (
            .O(N__21587),
            .I(\b2v_inst20.counterZ0Z_30 ));
    Odrv12 I__3267 (
            .O(N__21584),
            .I(\b2v_inst20.counterZ0Z_30 ));
    InMux I__3266 (
            .O(N__21579),
            .I(\b2v_inst20.counter_1_cry_29 ));
    InMux I__3265 (
            .O(N__21576),
            .I(\b2v_inst20.counter_1_cry_30 ));
    InMux I__3264 (
            .O(N__21573),
            .I(N__21569));
    InMux I__3263 (
            .O(N__21572),
            .I(N__21566));
    LocalMux I__3262 (
            .O(N__21569),
            .I(N__21563));
    LocalMux I__3261 (
            .O(N__21566),
            .I(\b2v_inst20.counterZ0Z_31 ));
    Odrv12 I__3260 (
            .O(N__21563),
            .I(\b2v_inst20.counterZ0Z_31 ));
    InMux I__3259 (
            .O(N__21558),
            .I(bfn_5_11_0_));
    InMux I__3258 (
            .O(N__21555),
            .I(\b2v_inst20.counter_1_cry_17 ));
    InMux I__3257 (
            .O(N__21552),
            .I(\b2v_inst20.counter_1_cry_18 ));
    InMux I__3256 (
            .O(N__21549),
            .I(N__21545));
    InMux I__3255 (
            .O(N__21548),
            .I(N__21542));
    LocalMux I__3254 (
            .O(N__21545),
            .I(\b2v_inst20.counterZ0Z_20 ));
    LocalMux I__3253 (
            .O(N__21542),
            .I(\b2v_inst20.counterZ0Z_20 ));
    InMux I__3252 (
            .O(N__21537),
            .I(\b2v_inst20.counter_1_cry_19 ));
    InMux I__3251 (
            .O(N__21534),
            .I(N__21530));
    InMux I__3250 (
            .O(N__21533),
            .I(N__21527));
    LocalMux I__3249 (
            .O(N__21530),
            .I(\b2v_inst20.counterZ0Z_21 ));
    LocalMux I__3248 (
            .O(N__21527),
            .I(\b2v_inst20.counterZ0Z_21 ));
    InMux I__3247 (
            .O(N__21522),
            .I(\b2v_inst20.counter_1_cry_20 ));
    CascadeMux I__3246 (
            .O(N__21519),
            .I(N__21515));
    InMux I__3245 (
            .O(N__21518),
            .I(N__21512));
    InMux I__3244 (
            .O(N__21515),
            .I(N__21509));
    LocalMux I__3243 (
            .O(N__21512),
            .I(\b2v_inst20.counterZ0Z_22 ));
    LocalMux I__3242 (
            .O(N__21509),
            .I(\b2v_inst20.counterZ0Z_22 ));
    InMux I__3241 (
            .O(N__21504),
            .I(\b2v_inst20.counter_1_cry_21 ));
    InMux I__3240 (
            .O(N__21501),
            .I(N__21497));
    InMux I__3239 (
            .O(N__21500),
            .I(N__21494));
    LocalMux I__3238 (
            .O(N__21497),
            .I(\b2v_inst20.counterZ0Z_23 ));
    LocalMux I__3237 (
            .O(N__21494),
            .I(\b2v_inst20.counterZ0Z_23 ));
    InMux I__3236 (
            .O(N__21489),
            .I(\b2v_inst20.counter_1_cry_22 ));
    InMux I__3235 (
            .O(N__21486),
            .I(\b2v_inst20.counter_1_cry_23 ));
    InMux I__3234 (
            .O(N__21483),
            .I(N__21479));
    InMux I__3233 (
            .O(N__21482),
            .I(N__21476));
    LocalMux I__3232 (
            .O(N__21479),
            .I(\b2v_inst20.counterZ0Z_8 ));
    LocalMux I__3231 (
            .O(N__21476),
            .I(\b2v_inst20.counterZ0Z_8 ));
    InMux I__3230 (
            .O(N__21471),
            .I(\b2v_inst20.counter_1_cry_7 ));
    InMux I__3229 (
            .O(N__21468),
            .I(N__21464));
    InMux I__3228 (
            .O(N__21467),
            .I(N__21461));
    LocalMux I__3227 (
            .O(N__21464),
            .I(\b2v_inst20.counterZ0Z_9 ));
    LocalMux I__3226 (
            .O(N__21461),
            .I(\b2v_inst20.counterZ0Z_9 ));
    InMux I__3225 (
            .O(N__21456),
            .I(bfn_5_10_0_));
    InMux I__3224 (
            .O(N__21453),
            .I(N__21449));
    InMux I__3223 (
            .O(N__21452),
            .I(N__21446));
    LocalMux I__3222 (
            .O(N__21449),
            .I(\b2v_inst20.counterZ0Z_10 ));
    LocalMux I__3221 (
            .O(N__21446),
            .I(\b2v_inst20.counterZ0Z_10 ));
    InMux I__3220 (
            .O(N__21441),
            .I(\b2v_inst20.counter_1_cry_9 ));
    CascadeMux I__3219 (
            .O(N__21438),
            .I(N__21434));
    InMux I__3218 (
            .O(N__21437),
            .I(N__21431));
    InMux I__3217 (
            .O(N__21434),
            .I(N__21428));
    LocalMux I__3216 (
            .O(N__21431),
            .I(\b2v_inst20.counterZ0Z_11 ));
    LocalMux I__3215 (
            .O(N__21428),
            .I(\b2v_inst20.counterZ0Z_11 ));
    InMux I__3214 (
            .O(N__21423),
            .I(\b2v_inst20.counter_1_cry_10 ));
    InMux I__3213 (
            .O(N__21420),
            .I(\b2v_inst20.counter_1_cry_11 ));
    InMux I__3212 (
            .O(N__21417),
            .I(\b2v_inst20.counter_1_cry_12 ));
    InMux I__3211 (
            .O(N__21414),
            .I(\b2v_inst20.counter_1_cry_13 ));
    InMux I__3210 (
            .O(N__21411),
            .I(\b2v_inst20.counter_1_cry_14 ));
    InMux I__3209 (
            .O(N__21408),
            .I(\b2v_inst20.counter_1_cry_15 ));
    InMux I__3208 (
            .O(N__21405),
            .I(N__21402));
    LocalMux I__3207 (
            .O(N__21402),
            .I(\b2v_inst200.HDA_SDO_ATP_0 ));
    CascadeMux I__3206 (
            .O(N__21399),
            .I(N__21396));
    InMux I__3205 (
            .O(N__21396),
            .I(N__21391));
    InMux I__3204 (
            .O(N__21395),
            .I(N__21386));
    InMux I__3203 (
            .O(N__21394),
            .I(N__21386));
    LocalMux I__3202 (
            .O(N__21391),
            .I(\b2v_inst200.N_205 ));
    LocalMux I__3201 (
            .O(N__21386),
            .I(\b2v_inst200.N_205 ));
    InMux I__3200 (
            .O(N__21381),
            .I(N__21372));
    InMux I__3199 (
            .O(N__21380),
            .I(N__21372));
    InMux I__3198 (
            .O(N__21379),
            .I(N__21372));
    LocalMux I__3197 (
            .O(N__21372),
            .I(\b2v_inst200.curr_state_i_2 ));
    IoInMux I__3196 (
            .O(N__21369),
            .I(N__21366));
    LocalMux I__3195 (
            .O(N__21366),
            .I(N__21363));
    Odrv12 I__3194 (
            .O(N__21363),
            .I(hda_sdo_atp));
    InMux I__3193 (
            .O(N__21360),
            .I(N__21351));
    InMux I__3192 (
            .O(N__21359),
            .I(N__21351));
    InMux I__3191 (
            .O(N__21358),
            .I(N__21351));
    LocalMux I__3190 (
            .O(N__21351),
            .I(N__21347));
    InMux I__3189 (
            .O(N__21350),
            .I(N__21344));
    Odrv12 I__3188 (
            .O(N__21347),
            .I(\b2v_inst200.N_282 ));
    LocalMux I__3187 (
            .O(N__21344),
            .I(\b2v_inst200.N_282 ));
    CascadeMux I__3186 (
            .O(N__21339),
            .I(N__21336));
    InMux I__3185 (
            .O(N__21336),
            .I(N__21332));
    CascadeMux I__3184 (
            .O(N__21335),
            .I(N__21329));
    LocalMux I__3183 (
            .O(N__21332),
            .I(N__21325));
    InMux I__3182 (
            .O(N__21329),
            .I(N__21320));
    InMux I__3181 (
            .O(N__21328),
            .I(N__21320));
    Odrv4 I__3180 (
            .O(N__21325),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__3179 (
            .O(N__21320),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    InMux I__3178 (
            .O(N__21315),
            .I(N__21309));
    InMux I__3177 (
            .O(N__21314),
            .I(N__21309));
    LocalMux I__3176 (
            .O(N__21309),
            .I(N__21304));
    InMux I__3175 (
            .O(N__21308),
            .I(N__21299));
    InMux I__3174 (
            .O(N__21307),
            .I(N__21299));
    Odrv4 I__3173 (
            .O(N__21304),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    LocalMux I__3172 (
            .O(N__21299),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    InMux I__3171 (
            .O(N__21294),
            .I(N__21291));
    LocalMux I__3170 (
            .O(N__21291),
            .I(N__21288));
    Span4Mux_v I__3169 (
            .O(N__21288),
            .I(N__21285));
    Odrv4 I__3168 (
            .O(N__21285),
            .I(\b2v_inst200.curr_state_3_1 ));
    InMux I__3167 (
            .O(N__21282),
            .I(\b2v_inst20.counter_1_cry_1 ));
    InMux I__3166 (
            .O(N__21279),
            .I(\b2v_inst20.counter_1_cry_2 ));
    InMux I__3165 (
            .O(N__21276),
            .I(\b2v_inst20.counter_1_cry_3 ));
    InMux I__3164 (
            .O(N__21273),
            .I(\b2v_inst20.counter_1_cry_4 ));
    InMux I__3163 (
            .O(N__21270),
            .I(\b2v_inst20.counter_1_cry_5 ));
    InMux I__3162 (
            .O(N__21267),
            .I(\b2v_inst20.counter_1_cry_6 ));
    InMux I__3161 (
            .O(N__21264),
            .I(N__21258));
    InMux I__3160 (
            .O(N__21263),
            .I(N__21258));
    LocalMux I__3159 (
            .O(N__21258),
            .I(\b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ));
    InMux I__3158 (
            .O(N__21255),
            .I(\b2v_inst11.un3_count_off_1_cry_13 ));
    InMux I__3157 (
            .O(N__21252),
            .I(N__21248));
    InMux I__3156 (
            .O(N__21251),
            .I(N__21245));
    LocalMux I__3155 (
            .O(N__21248),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    LocalMux I__3154 (
            .O(N__21245),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    InMux I__3153 (
            .O(N__21240),
            .I(\b2v_inst11.un3_count_off_1_cry_14 ));
    CascadeMux I__3152 (
            .O(N__21237),
            .I(N__21233));
    InMux I__3151 (
            .O(N__21236),
            .I(N__21228));
    InMux I__3150 (
            .O(N__21233),
            .I(N__21228));
    LocalMux I__3149 (
            .O(N__21228),
            .I(\b2v_inst11.count_offZ0Z_12 ));
    CascadeMux I__3148 (
            .O(N__21225),
            .I(N__21221));
    InMux I__3147 (
            .O(N__21224),
            .I(N__21216));
    InMux I__3146 (
            .O(N__21221),
            .I(N__21216));
    LocalMux I__3145 (
            .O(N__21216),
            .I(\b2v_inst11.count_offZ0Z_11 ));
    CascadeMux I__3144 (
            .O(N__21213),
            .I(N__21209));
    CascadeMux I__3143 (
            .O(N__21212),
            .I(N__21206));
    InMux I__3142 (
            .O(N__21209),
            .I(N__21201));
    InMux I__3141 (
            .O(N__21206),
            .I(N__21201));
    LocalMux I__3140 (
            .O(N__21201),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    CascadeMux I__3139 (
            .O(N__21198),
            .I(N__21194));
    InMux I__3138 (
            .O(N__21197),
            .I(N__21189));
    InMux I__3137 (
            .O(N__21194),
            .I(N__21189));
    LocalMux I__3136 (
            .O(N__21189),
            .I(\b2v_inst11.count_offZ0Z_9 ));
    CascadeMux I__3135 (
            .O(N__21186),
            .I(\b2v_inst200.curr_state_i_2_cascade_ ));
    InMux I__3134 (
            .O(N__21183),
            .I(N__21180));
    LocalMux I__3133 (
            .O(N__21180),
            .I(\b2v_inst200.i4_mux ));
    InMux I__3132 (
            .O(N__21177),
            .I(N__21173));
    InMux I__3131 (
            .O(N__21176),
            .I(N__21170));
    LocalMux I__3130 (
            .O(N__21173),
            .I(N__21167));
    LocalMux I__3129 (
            .O(N__21170),
            .I(\b2v_inst200.N_2989_i ));
    Odrv12 I__3128 (
            .O(N__21167),
            .I(\b2v_inst200.N_2989_i ));
    CascadeMux I__3127 (
            .O(N__21162),
            .I(\b2v_inst200.N_205_cascade_ ));
    InMux I__3126 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__3125 (
            .O(N__21156),
            .I(\b2v_inst200.curr_stateZ0Z_2 ));
    InMux I__3124 (
            .O(N__21153),
            .I(\b2v_inst11.un3_count_off_1_cry_5 ));
    InMux I__3123 (
            .O(N__21150),
            .I(\b2v_inst11.un3_count_off_1_cry_6 ));
    InMux I__3122 (
            .O(N__21147),
            .I(\b2v_inst11.un3_count_off_1_cry_7 ));
    InMux I__3121 (
            .O(N__21144),
            .I(bfn_5_7_0_));
    InMux I__3120 (
            .O(N__21141),
            .I(N__21137));
    InMux I__3119 (
            .O(N__21140),
            .I(N__21134));
    LocalMux I__3118 (
            .O(N__21137),
            .I(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ));
    LocalMux I__3117 (
            .O(N__21134),
            .I(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ));
    InMux I__3116 (
            .O(N__21129),
            .I(\b2v_inst11.un3_count_off_1_cry_9 ));
    InMux I__3115 (
            .O(N__21126),
            .I(N__21120));
    InMux I__3114 (
            .O(N__21125),
            .I(N__21120));
    LocalMux I__3113 (
            .O(N__21120),
            .I(\b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ));
    InMux I__3112 (
            .O(N__21117),
            .I(\b2v_inst11.un3_count_off_1_cry_10 ));
    CascadeMux I__3111 (
            .O(N__21114),
            .I(N__21111));
    InMux I__3110 (
            .O(N__21111),
            .I(N__21105));
    InMux I__3109 (
            .O(N__21110),
            .I(N__21105));
    LocalMux I__3108 (
            .O(N__21105),
            .I(\b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ));
    InMux I__3107 (
            .O(N__21102),
            .I(\b2v_inst11.un3_count_off_1_cry_11 ));
    CascadeMux I__3106 (
            .O(N__21099),
            .I(N__21095));
    InMux I__3105 (
            .O(N__21098),
            .I(N__21092));
    InMux I__3104 (
            .O(N__21095),
            .I(N__21089));
    LocalMux I__3103 (
            .O(N__21092),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    LocalMux I__3102 (
            .O(N__21089),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    InMux I__3101 (
            .O(N__21084),
            .I(N__21078));
    InMux I__3100 (
            .O(N__21083),
            .I(N__21078));
    LocalMux I__3099 (
            .O(N__21078),
            .I(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ));
    InMux I__3098 (
            .O(N__21075),
            .I(\b2v_inst11.un3_count_off_1_cry_12 ));
    CascadeMux I__3097 (
            .O(N__21072),
            .I(N__21069));
    InMux I__3096 (
            .O(N__21069),
            .I(N__21066));
    LocalMux I__3095 (
            .O(N__21066),
            .I(\b2v_inst11.count_offZ0Z_14 ));
    CascadeMux I__3094 (
            .O(N__21063),
            .I(\b2v_inst200.m6_i_0_cascade_ ));
    CascadeMux I__3093 (
            .O(N__21060),
            .I(\b2v_inst200.N_58_cascade_ ));
    CascadeMux I__3092 (
            .O(N__21057),
            .I(\b2v_inst200.curr_stateZ0Z_0_cascade_ ));
    InMux I__3091 (
            .O(N__21054),
            .I(N__21051));
    LocalMux I__3090 (
            .O(N__21051),
            .I(N__21046));
    InMux I__3089 (
            .O(N__21050),
            .I(N__21043));
    InMux I__3088 (
            .O(N__21049),
            .I(N__21040));
    Span4Mux_v I__3087 (
            .O(N__21046),
            .I(N__21037));
    LocalMux I__3086 (
            .O(N__21043),
            .I(N_411));
    LocalMux I__3085 (
            .O(N__21040),
            .I(N_411));
    Odrv4 I__3084 (
            .O(N__21037),
            .I(N_411));
    CascadeMux I__3083 (
            .O(N__21030),
            .I(N_411_cascade_));
    InMux I__3082 (
            .O(N__21027),
            .I(N__21024));
    LocalMux I__3081 (
            .O(N__21024),
            .I(\b2v_inst200.m6_i_0 ));
    InMux I__3080 (
            .O(N__21021),
            .I(N__21018));
    LocalMux I__3079 (
            .O(N__21018),
            .I(\b2v_inst200.curr_state_3_0 ));
    InMux I__3078 (
            .O(N__21015),
            .I(\b2v_inst11.un3_count_off_1_cry_1 ));
    CascadeMux I__3077 (
            .O(N__21012),
            .I(N__21008));
    InMux I__3076 (
            .O(N__21011),
            .I(N__21003));
    InMux I__3075 (
            .O(N__21008),
            .I(N__21003));
    LocalMux I__3074 (
            .O(N__21003),
            .I(N__21000));
    Odrv4 I__3073 (
            .O(N__21000),
            .I(\b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ));
    InMux I__3072 (
            .O(N__20997),
            .I(\b2v_inst11.un3_count_off_1_cry_2 ));
    InMux I__3071 (
            .O(N__20994),
            .I(\b2v_inst11.un3_count_off_1_cry_3 ));
    InMux I__3070 (
            .O(N__20991),
            .I(\b2v_inst11.un3_count_off_1_cry_4 ));
    InMux I__3069 (
            .O(N__20988),
            .I(\b2v_inst200.un2_count_1_cry_14 ));
    InMux I__3068 (
            .O(N__20985),
            .I(N__20982));
    LocalMux I__3067 (
            .O(N__20982),
            .I(N__20979));
    Odrv4 I__3066 (
            .O(N__20979),
            .I(\b2v_inst200.un2_count_1_axb_16 ));
    InMux I__3065 (
            .O(N__20976),
            .I(N__20967));
    InMux I__3064 (
            .O(N__20975),
            .I(N__20967));
    InMux I__3063 (
            .O(N__20974),
            .I(N__20967));
    LocalMux I__3062 (
            .O(N__20967),
            .I(N__20964));
    Span4Mux_s0_v I__3061 (
            .O(N__20964),
            .I(N__20961));
    Odrv4 I__3060 (
            .O(N__20961),
            .I(\b2v_inst200.count_1_16 ));
    InMux I__3059 (
            .O(N__20958),
            .I(\b2v_inst200.un2_count_1_cry_15 ));
    InMux I__3058 (
            .O(N__20955),
            .I(N__20951));
    CascadeMux I__3057 (
            .O(N__20954),
            .I(N__20948));
    LocalMux I__3056 (
            .O(N__20951),
            .I(N__20945));
    InMux I__3055 (
            .O(N__20948),
            .I(N__20942));
    Odrv4 I__3054 (
            .O(N__20945),
            .I(\b2v_inst200.countZ0Z_17 ));
    LocalMux I__3053 (
            .O(N__20942),
            .I(\b2v_inst200.countZ0Z_17 ));
    InMux I__3052 (
            .O(N__20937),
            .I(bfn_5_4_0_));
    InMux I__3051 (
            .O(N__20934),
            .I(N__20930));
    InMux I__3050 (
            .O(N__20933),
            .I(N__20927));
    LocalMux I__3049 (
            .O(N__20930),
            .I(N__20924));
    LocalMux I__3048 (
            .O(N__20927),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    Odrv4 I__3047 (
            .O(N__20924),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    InMux I__3046 (
            .O(N__20919),
            .I(N__20916));
    LocalMux I__3045 (
            .O(N__20916),
            .I(N__20913));
    Odrv4 I__3044 (
            .O(N__20913),
            .I(\b2v_inst200.count_0_17 ));
    CascadeMux I__3043 (
            .O(N__20910),
            .I(\b2v_inst200.N_56_cascade_ ));
    InMux I__3042 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__3041 (
            .O(N__20904),
            .I(N__20901));
    Span4Mux_v I__3040 (
            .O(N__20901),
            .I(N__20898));
    Span4Mux_h I__3039 (
            .O(N__20898),
            .I(N__20895));
    Odrv4 I__3038 (
            .O(N__20895),
            .I(gpio_fpga_soc_1));
    CascadeMux I__3037 (
            .O(N__20892),
            .I(\b2v_inst200.curr_stateZ0Z_1_cascade_ ));
    InMux I__3036 (
            .O(N__20889),
            .I(N__20885));
    InMux I__3035 (
            .O(N__20888),
            .I(N__20882));
    LocalMux I__3034 (
            .O(N__20885),
            .I(\b2v_inst200.countZ0Z_7 ));
    LocalMux I__3033 (
            .O(N__20882),
            .I(\b2v_inst200.countZ0Z_7 ));
    InMux I__3032 (
            .O(N__20877),
            .I(\b2v_inst200.un2_count_1_cry_6 ));
    InMux I__3031 (
            .O(N__20874),
            .I(\b2v_inst200.un2_count_1_cry_7 ));
    InMux I__3030 (
            .O(N__20871),
            .I(N__20868));
    LocalMux I__3029 (
            .O(N__20868),
            .I(\b2v_inst200.un2_count_1_axb_9 ));
    InMux I__3028 (
            .O(N__20865),
            .I(N__20856));
    InMux I__3027 (
            .O(N__20864),
            .I(N__20856));
    InMux I__3026 (
            .O(N__20863),
            .I(N__20856));
    LocalMux I__3025 (
            .O(N__20856),
            .I(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ));
    InMux I__3024 (
            .O(N__20853),
            .I(bfn_5_3_0_));
    InMux I__3023 (
            .O(N__20850),
            .I(\b2v_inst200.un2_count_1_cry_9 ));
    InMux I__3022 (
            .O(N__20847),
            .I(N__20844));
    LocalMux I__3021 (
            .O(N__20844),
            .I(N__20840));
    InMux I__3020 (
            .O(N__20843),
            .I(N__20837));
    Odrv4 I__3019 (
            .O(N__20840),
            .I(\b2v_inst200.countZ0Z_11 ));
    LocalMux I__3018 (
            .O(N__20837),
            .I(\b2v_inst200.countZ0Z_11 ));
    InMux I__3017 (
            .O(N__20832),
            .I(\b2v_inst200.un2_count_1_cry_10 ));
    InMux I__3016 (
            .O(N__20829),
            .I(N__20826));
    LocalMux I__3015 (
            .O(N__20826),
            .I(\b2v_inst200.countZ0Z_12 ));
    InMux I__3014 (
            .O(N__20823),
            .I(N__20817));
    InMux I__3013 (
            .O(N__20822),
            .I(N__20817));
    LocalMux I__3012 (
            .O(N__20817),
            .I(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ));
    InMux I__3011 (
            .O(N__20814),
            .I(\b2v_inst200.un2_count_1_cry_11 ));
    InMux I__3010 (
            .O(N__20811),
            .I(N__20808));
    LocalMux I__3009 (
            .O(N__20808),
            .I(\b2v_inst200.un2_count_1_axb_13 ));
    InMux I__3008 (
            .O(N__20805),
            .I(N__20796));
    InMux I__3007 (
            .O(N__20804),
            .I(N__20796));
    InMux I__3006 (
            .O(N__20803),
            .I(N__20796));
    LocalMux I__3005 (
            .O(N__20796),
            .I(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ));
    InMux I__3004 (
            .O(N__20793),
            .I(\b2v_inst200.un2_count_1_cry_12 ));
    InMux I__3003 (
            .O(N__20790),
            .I(N__20786));
    InMux I__3002 (
            .O(N__20789),
            .I(N__20783));
    LocalMux I__3001 (
            .O(N__20786),
            .I(N__20780));
    LocalMux I__3000 (
            .O(N__20783),
            .I(\b2v_inst200.countZ0Z_14 ));
    Odrv4 I__2999 (
            .O(N__20780),
            .I(\b2v_inst200.countZ0Z_14 ));
    InMux I__2998 (
            .O(N__20775),
            .I(\b2v_inst200.un2_count_1_cry_13 ));
    CascadeMux I__2997 (
            .O(N__20772),
            .I(\b2v_inst200.count_1_0_cascade_ ));
    CascadeMux I__2996 (
            .O(N__20769),
            .I(N__20765));
    InMux I__2995 (
            .O(N__20768),
            .I(N__20762));
    InMux I__2994 (
            .O(N__20765),
            .I(N__20759));
    LocalMux I__2993 (
            .O(N__20762),
            .I(\b2v_inst200.un2_count_1_axb_1 ));
    LocalMux I__2992 (
            .O(N__20759),
            .I(\b2v_inst200.un2_count_1_axb_1 ));
    InMux I__2991 (
            .O(N__20754),
            .I(N__20750));
    InMux I__2990 (
            .O(N__20753),
            .I(N__20747));
    LocalMux I__2989 (
            .O(N__20750),
            .I(N__20744));
    LocalMux I__2988 (
            .O(N__20747),
            .I(N__20741));
    Odrv12 I__2987 (
            .O(N__20744),
            .I(\b2v_inst200.countZ0Z_2 ));
    Odrv4 I__2986 (
            .O(N__20741),
            .I(\b2v_inst200.countZ0Z_2 ));
    InMux I__2985 (
            .O(N__20736),
            .I(\b2v_inst200.un2_count_1_cry_1 ));
    InMux I__2984 (
            .O(N__20733),
            .I(N__20730));
    LocalMux I__2983 (
            .O(N__20730),
            .I(\b2v_inst200.un2_count_1_axb_3 ));
    InMux I__2982 (
            .O(N__20727),
            .I(N__20720));
    InMux I__2981 (
            .O(N__20726),
            .I(N__20720));
    InMux I__2980 (
            .O(N__20725),
            .I(N__20717));
    LocalMux I__2979 (
            .O(N__20720),
            .I(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ));
    LocalMux I__2978 (
            .O(N__20717),
            .I(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ));
    InMux I__2977 (
            .O(N__20712),
            .I(\b2v_inst200.un2_count_1_cry_2 ));
    InMux I__2976 (
            .O(N__20709),
            .I(N__20705));
    InMux I__2975 (
            .O(N__20708),
            .I(N__20702));
    LocalMux I__2974 (
            .O(N__20705),
            .I(N__20697));
    LocalMux I__2973 (
            .O(N__20702),
            .I(N__20697));
    Odrv4 I__2972 (
            .O(N__20697),
            .I(\b2v_inst200.countZ0Z_4 ));
    InMux I__2971 (
            .O(N__20694),
            .I(\b2v_inst200.un2_count_1_cry_3 ));
    InMux I__2970 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__2969 (
            .O(N__20688),
            .I(\b2v_inst200.un2_count_1_axb_5 ));
    InMux I__2968 (
            .O(N__20685),
            .I(N__20680));
    InMux I__2967 (
            .O(N__20684),
            .I(N__20675));
    InMux I__2966 (
            .O(N__20683),
            .I(N__20675));
    LocalMux I__2965 (
            .O(N__20680),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    LocalMux I__2964 (
            .O(N__20675),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    InMux I__2963 (
            .O(N__20670),
            .I(\b2v_inst200.un2_count_1_cry_4 ));
    InMux I__2962 (
            .O(N__20667),
            .I(\b2v_inst200.un2_count_1_cry_5_cZ0 ));
    InMux I__2961 (
            .O(N__20664),
            .I(N__20661));
    LocalMux I__2960 (
            .O(N__20661),
            .I(\b2v_inst11.mult1_un124_sum_cry_5_s ));
    InMux I__2959 (
            .O(N__20658),
            .I(N__20655));
    LocalMux I__2958 (
            .O(N__20655),
            .I(N__20652));
    Odrv4 I__2957 (
            .O(N__20652),
            .I(\b2v_inst11.mult1_un131_sum_cry_6_s ));
    InMux I__2956 (
            .O(N__20649),
            .I(\b2v_inst11.mult1_un131_sum_cry_5 ));
    InMux I__2955 (
            .O(N__20646),
            .I(N__20643));
    LocalMux I__2954 (
            .O(N__20643),
            .I(\b2v_inst11.mult1_un124_sum_cry_6_s ));
    InMux I__2953 (
            .O(N__20640),
            .I(N__20637));
    LocalMux I__2952 (
            .O(N__20637),
            .I(N__20634));
    Odrv4 I__2951 (
            .O(N__20634),
            .I(\b2v_inst11.mult1_un138_sum_axb_8 ));
    InMux I__2950 (
            .O(N__20631),
            .I(\b2v_inst11.mult1_un131_sum_cry_6 ));
    CascadeMux I__2949 (
            .O(N__20628),
            .I(N__20625));
    InMux I__2948 (
            .O(N__20625),
            .I(N__20622));
    LocalMux I__2947 (
            .O(N__20622),
            .I(\b2v_inst11.mult1_un131_sum_axb_8 ));
    InMux I__2946 (
            .O(N__20619),
            .I(\b2v_inst11.mult1_un131_sum_cry_7 ));
    InMux I__2945 (
            .O(N__20616),
            .I(N__20612));
    CascadeMux I__2944 (
            .O(N__20615),
            .I(N__20609));
    LocalMux I__2943 (
            .O(N__20612),
            .I(N__20604));
    InMux I__2942 (
            .O(N__20609),
            .I(N__20596));
    InMux I__2941 (
            .O(N__20608),
            .I(N__20596));
    InMux I__2940 (
            .O(N__20607),
            .I(N__20596));
    Span4Mux_s3_h I__2939 (
            .O(N__20604),
            .I(N__20593));
    InMux I__2938 (
            .O(N__20603),
            .I(N__20590));
    LocalMux I__2937 (
            .O(N__20596),
            .I(N__20587));
    Odrv4 I__2936 (
            .O(N__20593),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__2935 (
            .O(N__20590),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    Odrv12 I__2934 (
            .O(N__20587),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    InMux I__2933 (
            .O(N__20580),
            .I(N__20577));
    LocalMux I__2932 (
            .O(N__20577),
            .I(N__20573));
    CascadeMux I__2931 (
            .O(N__20576),
            .I(N__20569));
    Span4Mux_s3_h I__2930 (
            .O(N__20573),
            .I(N__20564));
    InMux I__2929 (
            .O(N__20572),
            .I(N__20561));
    InMux I__2928 (
            .O(N__20569),
            .I(N__20554));
    InMux I__2927 (
            .O(N__20568),
            .I(N__20554));
    InMux I__2926 (
            .O(N__20567),
            .I(N__20554));
    Odrv4 I__2925 (
            .O(N__20564),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__2924 (
            .O(N__20561),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__2923 (
            .O(N__20554),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    CascadeMux I__2922 (
            .O(N__20547),
            .I(N__20543));
    CascadeMux I__2921 (
            .O(N__20546),
            .I(N__20539));
    InMux I__2920 (
            .O(N__20543),
            .I(N__20532));
    InMux I__2919 (
            .O(N__20542),
            .I(N__20532));
    InMux I__2918 (
            .O(N__20539),
            .I(N__20532));
    LocalMux I__2917 (
            .O(N__20532),
            .I(\b2v_inst11.mult1_un124_sum_i_0_8 ));
    InMux I__2916 (
            .O(N__20529),
            .I(N__20526));
    LocalMux I__2915 (
            .O(N__20526),
            .I(N__20523));
    Span4Mux_h I__2914 (
            .O(N__20523),
            .I(N__20520));
    Span4Mux_v I__2913 (
            .O(N__20520),
            .I(N__20516));
    InMux I__2912 (
            .O(N__20519),
            .I(N__20513));
    Odrv4 I__2911 (
            .O(N__20516),
            .I(\b2v_inst16.N_208_0 ));
    LocalMux I__2910 (
            .O(N__20513),
            .I(\b2v_inst16.N_208_0 ));
    InMux I__2909 (
            .O(N__20508),
            .I(N__20505));
    LocalMux I__2908 (
            .O(N__20505),
            .I(N__20502));
    Span12Mux_s8_h I__2907 (
            .O(N__20502),
            .I(N__20499));
    Odrv12 I__2906 (
            .O(N__20499),
            .I(\b2v_inst16.delayed_vddq_pwrgd_en ));
    CascadeMux I__2905 (
            .O(N__20496),
            .I(N__20493));
    InMux I__2904 (
            .O(N__20493),
            .I(N__20490));
    LocalMux I__2903 (
            .O(N__20490),
            .I(N__20487));
    Span4Mux_s0_v I__2902 (
            .O(N__20487),
            .I(N__20481));
    InMux I__2901 (
            .O(N__20486),
            .I(N__20478));
    InMux I__2900 (
            .O(N__20485),
            .I(N__20470));
    InMux I__2899 (
            .O(N__20484),
            .I(N__20470));
    Span4Mux_v I__2898 (
            .O(N__20481),
            .I(N__20465));
    LocalMux I__2897 (
            .O(N__20478),
            .I(N__20465));
    InMux I__2896 (
            .O(N__20477),
            .I(N__20462));
    InMux I__2895 (
            .O(N__20476),
            .I(N__20457));
    InMux I__2894 (
            .O(N__20475),
            .I(N__20457));
    LocalMux I__2893 (
            .O(N__20470),
            .I(N__20454));
    Span4Mux_h I__2892 (
            .O(N__20465),
            .I(N__20451));
    LocalMux I__2891 (
            .O(N__20462),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    LocalMux I__2890 (
            .O(N__20457),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    Odrv4 I__2889 (
            .O(N__20454),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    Odrv4 I__2888 (
            .O(N__20451),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    InMux I__2887 (
            .O(N__20442),
            .I(N__20439));
    LocalMux I__2886 (
            .O(N__20439),
            .I(N__20436));
    Span12Mux_s4_h I__2885 (
            .O(N__20436),
            .I(N__20432));
    InMux I__2884 (
            .O(N__20435),
            .I(N__20429));
    Odrv12 I__2883 (
            .O(N__20432),
            .I(\b2v_inst16.delayed_vddq_pwrgdZ0 ));
    LocalMux I__2882 (
            .O(N__20429),
            .I(\b2v_inst16.delayed_vddq_pwrgdZ0 ));
    InMux I__2881 (
            .O(N__20424),
            .I(N__20420));
    CascadeMux I__2880 (
            .O(N__20423),
            .I(N__20416));
    LocalMux I__2879 (
            .O(N__20420),
            .I(N__20412));
    InMux I__2878 (
            .O(N__20419),
            .I(N__20407));
    InMux I__2877 (
            .O(N__20416),
            .I(N__20407));
    InMux I__2876 (
            .O(N__20415),
            .I(N__20404));
    Odrv4 I__2875 (
            .O(N__20412),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__2874 (
            .O(N__20407),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__2873 (
            .O(N__20404),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    CascadeMux I__2872 (
            .O(N__20397),
            .I(N__20394));
    InMux I__2871 (
            .O(N__20394),
            .I(N__20391));
    LocalMux I__2870 (
            .O(N__20391),
            .I(\b2v_inst11.mult1_un117_sum_cry_5_s ));
    InMux I__2869 (
            .O(N__20388),
            .I(\b2v_inst11.mult1_un124_sum_cry_5 ));
    InMux I__2868 (
            .O(N__20385),
            .I(N__20382));
    LocalMux I__2867 (
            .O(N__20382),
            .I(\b2v_inst11.mult1_un117_sum_cry_6_s ));
    CascadeMux I__2866 (
            .O(N__20379),
            .I(N__20375));
    CascadeMux I__2865 (
            .O(N__20378),
            .I(N__20371));
    InMux I__2864 (
            .O(N__20375),
            .I(N__20364));
    InMux I__2863 (
            .O(N__20374),
            .I(N__20364));
    InMux I__2862 (
            .O(N__20371),
            .I(N__20364));
    LocalMux I__2861 (
            .O(N__20364),
            .I(\b2v_inst11.mult1_un117_sum_i_0_8 ));
    InMux I__2860 (
            .O(N__20361),
            .I(\b2v_inst11.mult1_un124_sum_cry_6 ));
    CascadeMux I__2859 (
            .O(N__20358),
            .I(N__20355));
    InMux I__2858 (
            .O(N__20355),
            .I(N__20352));
    LocalMux I__2857 (
            .O(N__20352),
            .I(\b2v_inst11.mult1_un124_sum_axb_8 ));
    InMux I__2856 (
            .O(N__20349),
            .I(\b2v_inst11.mult1_un124_sum_cry_7 ));
    InMux I__2855 (
            .O(N__20346),
            .I(N__20343));
    LocalMux I__2854 (
            .O(N__20343),
            .I(\b2v_inst11.mult1_un117_sum_i ));
    CascadeMux I__2853 (
            .O(N__20340),
            .I(N__20337));
    InMux I__2852 (
            .O(N__20337),
            .I(N__20334));
    LocalMux I__2851 (
            .O(N__20334),
            .I(N__20331));
    Odrv4 I__2850 (
            .O(N__20331),
            .I(\b2v_inst11.mult1_un131_sum_cry_3_s ));
    InMux I__2849 (
            .O(N__20328),
            .I(\b2v_inst11.mult1_un131_sum_cry_2 ));
    CascadeMux I__2848 (
            .O(N__20325),
            .I(N__20322));
    InMux I__2847 (
            .O(N__20322),
            .I(N__20319));
    LocalMux I__2846 (
            .O(N__20319),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    CascadeMux I__2845 (
            .O(N__20316),
            .I(N__20313));
    InMux I__2844 (
            .O(N__20313),
            .I(N__20310));
    LocalMux I__2843 (
            .O(N__20310),
            .I(N__20307));
    Odrv4 I__2842 (
            .O(N__20307),
            .I(\b2v_inst11.mult1_un131_sum_cry_4_s ));
    InMux I__2841 (
            .O(N__20304),
            .I(\b2v_inst11.mult1_un131_sum_cry_3 ));
    CascadeMux I__2840 (
            .O(N__20301),
            .I(N__20298));
    InMux I__2839 (
            .O(N__20298),
            .I(N__20295));
    LocalMux I__2838 (
            .O(N__20295),
            .I(\b2v_inst11.mult1_un124_sum_cry_4_s ));
    InMux I__2837 (
            .O(N__20292),
            .I(N__20289));
    LocalMux I__2836 (
            .O(N__20289),
            .I(N__20286));
    Odrv4 I__2835 (
            .O(N__20286),
            .I(\b2v_inst11.mult1_un131_sum_cry_5_s ));
    InMux I__2834 (
            .O(N__20283),
            .I(\b2v_inst11.mult1_un131_sum_cry_4 ));
    InMux I__2833 (
            .O(N__20280),
            .I(\b2v_inst11.mult1_un117_sum_cry_4 ));
    InMux I__2832 (
            .O(N__20277),
            .I(\b2v_inst11.mult1_un117_sum_cry_5 ));
    InMux I__2831 (
            .O(N__20274),
            .I(\b2v_inst11.mult1_un117_sum_cry_6 ));
    InMux I__2830 (
            .O(N__20271),
            .I(\b2v_inst11.mult1_un117_sum_cry_7 ));
    CascadeMux I__2829 (
            .O(N__20268),
            .I(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ));
    InMux I__2828 (
            .O(N__20265),
            .I(\b2v_inst11.mult1_un124_sum_cry_2 ));
    CascadeMux I__2827 (
            .O(N__20262),
            .I(N__20259));
    InMux I__2826 (
            .O(N__20259),
            .I(N__20256));
    LocalMux I__2825 (
            .O(N__20256),
            .I(\b2v_inst11.mult1_un117_sum_cry_3_s ));
    InMux I__2824 (
            .O(N__20253),
            .I(\b2v_inst11.mult1_un124_sum_cry_3 ));
    InMux I__2823 (
            .O(N__20250),
            .I(N__20247));
    LocalMux I__2822 (
            .O(N__20247),
            .I(\b2v_inst11.mult1_un117_sum_cry_4_s ));
    InMux I__2821 (
            .O(N__20244),
            .I(\b2v_inst11.mult1_un124_sum_cry_4 ));
    CascadeMux I__2820 (
            .O(N__20241),
            .I(N__20238));
    InMux I__2819 (
            .O(N__20238),
            .I(N__20235));
    LocalMux I__2818 (
            .O(N__20235),
            .I(\b2v_inst11.mult1_un138_sum_cry_4_s ));
    InMux I__2817 (
            .O(N__20232),
            .I(\b2v_inst11.mult1_un138_sum_cry_3 ));
    InMux I__2816 (
            .O(N__20229),
            .I(N__20226));
    LocalMux I__2815 (
            .O(N__20226),
            .I(\b2v_inst11.mult1_un138_sum_cry_5_s ));
    InMux I__2814 (
            .O(N__20223),
            .I(\b2v_inst11.mult1_un138_sum_cry_4 ));
    InMux I__2813 (
            .O(N__20220),
            .I(N__20217));
    LocalMux I__2812 (
            .O(N__20217),
            .I(\b2v_inst11.mult1_un138_sum_cry_6_s ));
    InMux I__2811 (
            .O(N__20214),
            .I(\b2v_inst11.mult1_un138_sum_cry_5 ));
    CascadeMux I__2810 (
            .O(N__20211),
            .I(N__20208));
    InMux I__2809 (
            .O(N__20208),
            .I(N__20205));
    LocalMux I__2808 (
            .O(N__20205),
            .I(\b2v_inst11.mult1_un145_sum_axb_8 ));
    InMux I__2807 (
            .O(N__20202),
            .I(\b2v_inst11.mult1_un138_sum_cry_6 ));
    InMux I__2806 (
            .O(N__20199),
            .I(\b2v_inst11.mult1_un138_sum_cry_7 ));
    InMux I__2805 (
            .O(N__20196),
            .I(N__20193));
    LocalMux I__2804 (
            .O(N__20193),
            .I(N__20189));
    CascadeMux I__2803 (
            .O(N__20192),
            .I(N__20185));
    Span4Mux_s3_h I__2802 (
            .O(N__20189),
            .I(N__20180));
    InMux I__2801 (
            .O(N__20188),
            .I(N__20177));
    InMux I__2800 (
            .O(N__20185),
            .I(N__20170));
    InMux I__2799 (
            .O(N__20184),
            .I(N__20170));
    InMux I__2798 (
            .O(N__20183),
            .I(N__20170));
    Odrv4 I__2797 (
            .O(N__20180),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__2796 (
            .O(N__20177),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__2795 (
            .O(N__20170),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    CascadeMux I__2794 (
            .O(N__20163),
            .I(N__20159));
    CascadeMux I__2793 (
            .O(N__20162),
            .I(N__20155));
    InMux I__2792 (
            .O(N__20159),
            .I(N__20148));
    InMux I__2791 (
            .O(N__20158),
            .I(N__20148));
    InMux I__2790 (
            .O(N__20155),
            .I(N__20148));
    LocalMux I__2789 (
            .O(N__20148),
            .I(\b2v_inst11.mult1_un131_sum_i_0_8 ));
    InMux I__2788 (
            .O(N__20145),
            .I(\b2v_inst11.mult1_un117_sum_cry_2 ));
    InMux I__2787 (
            .O(N__20142),
            .I(\b2v_inst11.mult1_un117_sum_cry_3 ));
    InMux I__2786 (
            .O(N__20139),
            .I(\b2v_inst11.mult1_un145_sum_cry_2 ));
    InMux I__2785 (
            .O(N__20136),
            .I(\b2v_inst11.mult1_un145_sum_cry_3 ));
    InMux I__2784 (
            .O(N__20133),
            .I(\b2v_inst11.mult1_un145_sum_cry_4 ));
    InMux I__2783 (
            .O(N__20130),
            .I(\b2v_inst11.mult1_un145_sum_cry_5 ));
    InMux I__2782 (
            .O(N__20127),
            .I(\b2v_inst11.mult1_un145_sum_cry_6 ));
    InMux I__2781 (
            .O(N__20124),
            .I(\b2v_inst11.mult1_un145_sum_cry_7 ));
    CascadeMux I__2780 (
            .O(N__20121),
            .I(N__20117));
    CascadeMux I__2779 (
            .O(N__20120),
            .I(N__20113));
    InMux I__2778 (
            .O(N__20117),
            .I(N__20106));
    InMux I__2777 (
            .O(N__20116),
            .I(N__20106));
    InMux I__2776 (
            .O(N__20113),
            .I(N__20106));
    LocalMux I__2775 (
            .O(N__20106),
            .I(\b2v_inst11.mult1_un138_sum_i_0_8 ));
    CascadeMux I__2774 (
            .O(N__20103),
            .I(N__20100));
    InMux I__2773 (
            .O(N__20100),
            .I(N__20097));
    LocalMux I__2772 (
            .O(N__20097),
            .I(\b2v_inst11.mult1_un138_sum_cry_3_s ));
    InMux I__2771 (
            .O(N__20094),
            .I(\b2v_inst11.mult1_un138_sum_cry_2 ));
    InMux I__2770 (
            .O(N__20091),
            .I(N__20088));
    LocalMux I__2769 (
            .O(N__20088),
            .I(N__20081));
    InMux I__2768 (
            .O(N__20087),
            .I(N__20074));
    InMux I__2767 (
            .O(N__20086),
            .I(N__20074));
    InMux I__2766 (
            .O(N__20085),
            .I(N__20074));
    InMux I__2765 (
            .O(N__20084),
            .I(N__20071));
    Odrv4 I__2764 (
            .O(N__20081),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__2763 (
            .O(N__20074),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__2762 (
            .O(N__20071),
            .I(\b2v_inst11.countZ0Z_0 ));
    InMux I__2761 (
            .O(N__20064),
            .I(N__20043));
    InMux I__2760 (
            .O(N__20063),
            .I(N__20043));
    InMux I__2759 (
            .O(N__20062),
            .I(N__20043));
    InMux I__2758 (
            .O(N__20061),
            .I(N__20034));
    InMux I__2757 (
            .O(N__20060),
            .I(N__20034));
    InMux I__2756 (
            .O(N__20059),
            .I(N__20034));
    InMux I__2755 (
            .O(N__20058),
            .I(N__20034));
    InMux I__2754 (
            .O(N__20057),
            .I(N__20031));
    InMux I__2753 (
            .O(N__20056),
            .I(N__20022));
    InMux I__2752 (
            .O(N__20055),
            .I(N__20022));
    InMux I__2751 (
            .O(N__20054),
            .I(N__20022));
    InMux I__2750 (
            .O(N__20053),
            .I(N__20022));
    InMux I__2749 (
            .O(N__20052),
            .I(N__20015));
    InMux I__2748 (
            .O(N__20051),
            .I(N__20015));
    InMux I__2747 (
            .O(N__20050),
            .I(N__20015));
    LocalMux I__2746 (
            .O(N__20043),
            .I(N__20007));
    LocalMux I__2745 (
            .O(N__20034),
            .I(N__20007));
    LocalMux I__2744 (
            .O(N__20031),
            .I(N__20004));
    LocalMux I__2743 (
            .O(N__20022),
            .I(N__19999));
    LocalMux I__2742 (
            .O(N__20015),
            .I(N__19999));
    InMux I__2741 (
            .O(N__20014),
            .I(N__19992));
    InMux I__2740 (
            .O(N__20013),
            .I(N__19992));
    InMux I__2739 (
            .O(N__20012),
            .I(N__19992));
    Span4Mux_v I__2738 (
            .O(N__20007),
            .I(N__19987));
    Span4Mux_h I__2737 (
            .O(N__20004),
            .I(N__19987));
    Odrv4 I__2736 (
            .O(N__19999),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    LocalMux I__2735 (
            .O(N__19992),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__2734 (
            .O(N__19987),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    InMux I__2733 (
            .O(N__19980),
            .I(N__19977));
    LocalMux I__2732 (
            .O(N__19977),
            .I(N__19974));
    Odrv4 I__2731 (
            .O(N__19974),
            .I(\b2v_inst11.count_1_0 ));
    CascadeMux I__2730 (
            .O(N__19971),
            .I(N__19967));
    CascadeMux I__2729 (
            .O(N__19970),
            .I(N__19963));
    InMux I__2728 (
            .O(N__19967),
            .I(N__19956));
    InMux I__2727 (
            .O(N__19966),
            .I(N__19956));
    InMux I__2726 (
            .O(N__19963),
            .I(N__19956));
    LocalMux I__2725 (
            .O(N__19956),
            .I(G_2848));
    InMux I__2724 (
            .O(N__19953),
            .I(\b2v_inst11.mult1_un166_sum_cry_5 ));
    InMux I__2723 (
            .O(N__19950),
            .I(N__19945));
    InMux I__2722 (
            .O(N__19949),
            .I(N__19942));
    InMux I__2721 (
            .O(N__19948),
            .I(N__19939));
    LocalMux I__2720 (
            .O(N__19945),
            .I(N__19936));
    LocalMux I__2719 (
            .O(N__19942),
            .I(N__19933));
    LocalMux I__2718 (
            .O(N__19939),
            .I(N__19930));
    Span4Mux_s3_h I__2717 (
            .O(N__19936),
            .I(N__19925));
    Span4Mux_s3_h I__2716 (
            .O(N__19933),
            .I(N__19925));
    Odrv4 I__2715 (
            .O(N__19930),
            .I(\b2v_inst11.mult1_un166_sum_s_6 ));
    Odrv4 I__2714 (
            .O(N__19925),
            .I(\b2v_inst11.mult1_un166_sum_s_6 ));
    SRMux I__2713 (
            .O(N__19920),
            .I(N__19917));
    LocalMux I__2712 (
            .O(N__19917),
            .I(N__19914));
    Span4Mux_h I__2711 (
            .O(N__19914),
            .I(N__19911));
    Odrv4 I__2710 (
            .O(N__19911),
            .I(\b2v_inst11.g0_0_0_rep1_1 ));
    InMux I__2709 (
            .O(N__19908),
            .I(N__19902));
    InMux I__2708 (
            .O(N__19907),
            .I(N__19902));
    LocalMux I__2707 (
            .O(N__19902),
            .I(\b2v_inst11.pwm_outZ0 ));
    CascadeMux I__2706 (
            .O(N__19899),
            .I(N__19896));
    InMux I__2705 (
            .O(N__19896),
            .I(N__19890));
    InMux I__2704 (
            .O(N__19895),
            .I(N__19890));
    LocalMux I__2703 (
            .O(N__19890),
            .I(N__19887));
    Odrv4 I__2702 (
            .O(N__19887),
            .I(\b2v_inst11.g0_i_a3_0_1 ));
    InMux I__2701 (
            .O(N__19884),
            .I(N__19881));
    LocalMux I__2700 (
            .O(N__19881),
            .I(\b2v_inst11.N_6 ));
    IoInMux I__2699 (
            .O(N__19878),
            .I(N__19875));
    LocalMux I__2698 (
            .O(N__19875),
            .I(N__19872));
    IoSpan4Mux I__2697 (
            .O(N__19872),
            .I(N__19869));
    IoSpan4Mux I__2696 (
            .O(N__19869),
            .I(N__19866));
    Span4Mux_s2_h I__2695 (
            .O(N__19866),
            .I(N__19863));
    Odrv4 I__2694 (
            .O(N__19863),
            .I(pwrbtn_led));
    IoInMux I__2693 (
            .O(N__19860),
            .I(N__19857));
    LocalMux I__2692 (
            .O(N__19857),
            .I(N__19854));
    Odrv12 I__2691 (
            .O(N__19854),
            .I(\b2v_inst200.count_enZ0 ));
    CascadeMux I__2690 (
            .O(N__19851),
            .I(\b2v_inst16.delayed_vddq_pwrgd_en_cascade_ ));
    IoInMux I__2689 (
            .O(N__19848),
            .I(N__19845));
    LocalMux I__2688 (
            .O(N__19845),
            .I(N__19842));
    Span4Mux_s1_h I__2687 (
            .O(N__19842),
            .I(N__19839));
    Span4Mux_v I__2686 (
            .O(N__19839),
            .I(N__19836));
    Sp12to4 I__2685 (
            .O(N__19836),
            .I(N__19833));
    Odrv12 I__2684 (
            .O(N__19833),
            .I(vpp_en));
    InMux I__2683 (
            .O(N__19830),
            .I(N__19826));
    InMux I__2682 (
            .O(N__19829),
            .I(N__19823));
    LocalMux I__2681 (
            .O(N__19826),
            .I(N__19820));
    LocalMux I__2680 (
            .O(N__19823),
            .I(\b2v_inst16.curr_state_RNIBO6I1Z0Z_0 ));
    Odrv4 I__2679 (
            .O(N__19820),
            .I(\b2v_inst16.curr_state_RNIBO6I1Z0Z_0 ));
    InMux I__2678 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__2677 (
            .O(N__19812),
            .I(\b2v_inst16.N_268 ));
    CascadeMux I__2676 (
            .O(N__19809),
            .I(\b2v_inst16.N_268_cascade_ ));
    CascadeMux I__2675 (
            .O(N__19806),
            .I(N__19799));
    InMux I__2674 (
            .O(N__19805),
            .I(N__19786));
    InMux I__2673 (
            .O(N__19804),
            .I(N__19786));
    InMux I__2672 (
            .O(N__19803),
            .I(N__19786));
    InMux I__2671 (
            .O(N__19802),
            .I(N__19786));
    InMux I__2670 (
            .O(N__19799),
            .I(N__19786));
    InMux I__2669 (
            .O(N__19798),
            .I(N__19783));
    InMux I__2668 (
            .O(N__19797),
            .I(N__19759));
    LocalMux I__2667 (
            .O(N__19786),
            .I(N__19754));
    LocalMux I__2666 (
            .O(N__19783),
            .I(N__19754));
    InMux I__2665 (
            .O(N__19782),
            .I(N__19749));
    InMux I__2664 (
            .O(N__19781),
            .I(N__19749));
    InMux I__2663 (
            .O(N__19780),
            .I(N__19746));
    InMux I__2662 (
            .O(N__19779),
            .I(N__19735));
    InMux I__2661 (
            .O(N__19778),
            .I(N__19735));
    InMux I__2660 (
            .O(N__19777),
            .I(N__19735));
    InMux I__2659 (
            .O(N__19776),
            .I(N__19735));
    InMux I__2658 (
            .O(N__19775),
            .I(N__19735));
    InMux I__2657 (
            .O(N__19774),
            .I(N__19726));
    InMux I__2656 (
            .O(N__19773),
            .I(N__19726));
    InMux I__2655 (
            .O(N__19772),
            .I(N__19726));
    InMux I__2654 (
            .O(N__19771),
            .I(N__19726));
    InMux I__2653 (
            .O(N__19770),
            .I(N__19715));
    InMux I__2652 (
            .O(N__19769),
            .I(N__19715));
    InMux I__2651 (
            .O(N__19768),
            .I(N__19715));
    InMux I__2650 (
            .O(N__19767),
            .I(N__19715));
    InMux I__2649 (
            .O(N__19766),
            .I(N__19715));
    InMux I__2648 (
            .O(N__19765),
            .I(N__19706));
    InMux I__2647 (
            .O(N__19764),
            .I(N__19706));
    InMux I__2646 (
            .O(N__19763),
            .I(N__19706));
    InMux I__2645 (
            .O(N__19762),
            .I(N__19706));
    LocalMux I__2644 (
            .O(N__19759),
            .I(N__19701));
    Span4Mux_s2_h I__2643 (
            .O(N__19754),
            .I(N__19701));
    LocalMux I__2642 (
            .O(N__19749),
            .I(N__19698));
    LocalMux I__2641 (
            .O(N__19746),
            .I(N__19695));
    LocalMux I__2640 (
            .O(N__19735),
            .I(N__19692));
    LocalMux I__2639 (
            .O(N__19726),
            .I(N__19689));
    LocalMux I__2638 (
            .O(N__19715),
            .I(N__19684));
    LocalMux I__2637 (
            .O(N__19706),
            .I(N__19684));
    Span4Mux_v I__2636 (
            .O(N__19701),
            .I(N__19681));
    Span4Mux_s3_h I__2635 (
            .O(N__19698),
            .I(N__19676));
    Span4Mux_s3_h I__2634 (
            .O(N__19695),
            .I(N__19676));
    Span4Mux_s3_h I__2633 (
            .O(N__19692),
            .I(N__19671));
    Span4Mux_s3_h I__2632 (
            .O(N__19689),
            .I(N__19671));
    Span4Mux_s3_h I__2631 (
            .O(N__19684),
            .I(N__19668));
    Odrv4 I__2630 (
            .O(N__19681),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2629 (
            .O(N__19676),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2628 (
            .O(N__19671),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__2627 (
            .O(N__19668),
            .I(\b2v_inst16.N_26 ));
    InMux I__2626 (
            .O(N__19659),
            .I(N__19656));
    LocalMux I__2625 (
            .O(N__19656),
            .I(\b2v_inst11.count_off_0_3 ));
    InMux I__2624 (
            .O(N__19653),
            .I(N__19650));
    LocalMux I__2623 (
            .O(N__19650),
            .I(N__19647));
    Odrv4 I__2622 (
            .O(N__19647),
            .I(\b2v_inst11.count_off_0_14 ));
    CascadeMux I__2621 (
            .O(N__19644),
            .I(\b2v_inst11.count_offZ0Z_14_cascade_ ));
    InMux I__2620 (
            .O(N__19641),
            .I(N__19638));
    LocalMux I__2619 (
            .O(N__19638),
            .I(\b2v_inst11.count_off_0_13 ));
    InMux I__2618 (
            .O(N__19635),
            .I(N__19632));
    LocalMux I__2617 (
            .O(N__19632),
            .I(N__19629));
    Odrv4 I__2616 (
            .O(N__19629),
            .I(\b2v_inst11.g0_i_o3_0 ));
    CascadeMux I__2615 (
            .O(N__19626),
            .I(N__19621));
    CascadeMux I__2614 (
            .O(N__19625),
            .I(N__19618));
    InMux I__2613 (
            .O(N__19624),
            .I(N__19613));
    InMux I__2612 (
            .O(N__19621),
            .I(N__19613));
    InMux I__2611 (
            .O(N__19618),
            .I(N__19610));
    LocalMux I__2610 (
            .O(N__19613),
            .I(N__19605));
    LocalMux I__2609 (
            .O(N__19610),
            .I(N__19605));
    Span4Mux_h I__2608 (
            .O(N__19605),
            .I(N__19602));
    Span4Mux_v I__2607 (
            .O(N__19602),
            .I(N__19599));
    Odrv4 I__2606 (
            .O(N__19599),
            .I(\b2v_inst11.un85_clk_100khz1_THRU_CO ));
    InMux I__2605 (
            .O(N__19596),
            .I(N__19591));
    InMux I__2604 (
            .O(N__19595),
            .I(N__19586));
    InMux I__2603 (
            .O(N__19594),
            .I(N__19586));
    LocalMux I__2602 (
            .O(N__19591),
            .I(N__19583));
    LocalMux I__2601 (
            .O(N__19586),
            .I(N__19580));
    Span4Mux_v I__2600 (
            .O(N__19583),
            .I(N__19577));
    Span4Mux_v I__2599 (
            .O(N__19580),
            .I(N__19574));
    Span4Mux_h I__2598 (
            .O(N__19577),
            .I(N__19571));
    Odrv4 I__2597 (
            .O(N__19574),
            .I(\b2v_inst11.un85_clk_100khz0_THRU_CO ));
    Odrv4 I__2596 (
            .O(N__19571),
            .I(\b2v_inst11.un85_clk_100khz0_THRU_CO ));
    CascadeMux I__2595 (
            .O(N__19566),
            .I(\b2v_inst11.N_6_cascade_ ));
    CascadeMux I__2594 (
            .O(N__19563),
            .I(\b2v_inst36.curr_stateZ0Z_0_cascade_ ));
    InMux I__2593 (
            .O(N__19560),
            .I(N__19550));
    InMux I__2592 (
            .O(N__19559),
            .I(N__19550));
    SRMux I__2591 (
            .O(N__19558),
            .I(N__19550));
    SRMux I__2590 (
            .O(N__19557),
            .I(N__19544));
    LocalMux I__2589 (
            .O(N__19550),
            .I(N__19538));
    InMux I__2588 (
            .O(N__19549),
            .I(N__19531));
    InMux I__2587 (
            .O(N__19548),
            .I(N__19531));
    SRMux I__2586 (
            .O(N__19547),
            .I(N__19531));
    LocalMux I__2585 (
            .O(N__19544),
            .I(N__19527));
    CascadeMux I__2584 (
            .O(N__19543),
            .I(N__19521));
    SRMux I__2583 (
            .O(N__19542),
            .I(N__19518));
    SRMux I__2582 (
            .O(N__19541),
            .I(N__19515));
    Span4Mux_v I__2581 (
            .O(N__19538),
            .I(N__19510));
    LocalMux I__2580 (
            .O(N__19531),
            .I(N__19510));
    SRMux I__2579 (
            .O(N__19530),
            .I(N__19502));
    Span4Mux_s1_h I__2578 (
            .O(N__19527),
            .I(N__19499));
    InMux I__2577 (
            .O(N__19526),
            .I(N__19492));
    InMux I__2576 (
            .O(N__19525),
            .I(N__19492));
    InMux I__2575 (
            .O(N__19524),
            .I(N__19492));
    InMux I__2574 (
            .O(N__19521),
            .I(N__19489));
    LocalMux I__2573 (
            .O(N__19518),
            .I(N__19486));
    LocalMux I__2572 (
            .O(N__19515),
            .I(N__19481));
    Span4Mux_s1_v I__2571 (
            .O(N__19510),
            .I(N__19481));
    InMux I__2570 (
            .O(N__19509),
            .I(N__19472));
    InMux I__2569 (
            .O(N__19508),
            .I(N__19472));
    InMux I__2568 (
            .O(N__19507),
            .I(N__19472));
    InMux I__2567 (
            .O(N__19506),
            .I(N__19472));
    SRMux I__2566 (
            .O(N__19505),
            .I(N__19464));
    LocalMux I__2565 (
            .O(N__19502),
            .I(N__19453));
    IoSpan4Mux I__2564 (
            .O(N__19499),
            .I(N__19446));
    LocalMux I__2563 (
            .O(N__19492),
            .I(N__19446));
    LocalMux I__2562 (
            .O(N__19489),
            .I(N__19446));
    Span4Mux_v I__2561 (
            .O(N__19486),
            .I(N__19437));
    Span4Mux_s1_h I__2560 (
            .O(N__19481),
            .I(N__19437));
    LocalMux I__2559 (
            .O(N__19472),
            .I(N__19437));
    InMux I__2558 (
            .O(N__19471),
            .I(N__19434));
    InMux I__2557 (
            .O(N__19470),
            .I(N__19427));
    InMux I__2556 (
            .O(N__19469),
            .I(N__19427));
    InMux I__2555 (
            .O(N__19468),
            .I(N__19427));
    InMux I__2554 (
            .O(N__19467),
            .I(N__19424));
    LocalMux I__2553 (
            .O(N__19464),
            .I(N__19421));
    InMux I__2552 (
            .O(N__19463),
            .I(N__19416));
    InMux I__2551 (
            .O(N__19462),
            .I(N__19416));
    InMux I__2550 (
            .O(N__19461),
            .I(N__19409));
    InMux I__2549 (
            .O(N__19460),
            .I(N__19409));
    InMux I__2548 (
            .O(N__19459),
            .I(N__19409));
    InMux I__2547 (
            .O(N__19458),
            .I(N__19402));
    InMux I__2546 (
            .O(N__19457),
            .I(N__19402));
    InMux I__2545 (
            .O(N__19456),
            .I(N__19402));
    Span4Mux_v I__2544 (
            .O(N__19453),
            .I(N__19397));
    Span4Mux_s2_v I__2543 (
            .O(N__19446),
            .I(N__19397));
    InMux I__2542 (
            .O(N__19445),
            .I(N__19392));
    InMux I__2541 (
            .O(N__19444),
            .I(N__19392));
    Sp12to4 I__2540 (
            .O(N__19437),
            .I(N__19385));
    LocalMux I__2539 (
            .O(N__19434),
            .I(N__19385));
    LocalMux I__2538 (
            .O(N__19427),
            .I(N__19385));
    LocalMux I__2537 (
            .O(N__19424),
            .I(N__19382));
    IoSpan4Mux I__2536 (
            .O(N__19421),
            .I(N__19377));
    LocalMux I__2535 (
            .O(N__19416),
            .I(N__19377));
    LocalMux I__2534 (
            .O(N__19409),
            .I(N__19368));
    LocalMux I__2533 (
            .O(N__19402),
            .I(N__19368));
    IoSpan4Mux I__2532 (
            .O(N__19397),
            .I(N__19368));
    LocalMux I__2531 (
            .O(N__19392),
            .I(N__19368));
    Span12Mux_s5_v I__2530 (
            .O(N__19385),
            .I(N__19365));
    Span4Mux_s3_h I__2529 (
            .O(N__19382),
            .I(N__19362));
    Span4Mux_s3_h I__2528 (
            .O(N__19377),
            .I(N__19357));
    Span4Mux_s3_h I__2527 (
            .O(N__19368),
            .I(N__19357));
    Odrv12 I__2526 (
            .O(N__19365),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__2525 (
            .O(N__19362),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__2524 (
            .O(N__19357),
            .I(\b2v_inst36.count_0_sqmuxa ));
    InMux I__2523 (
            .O(N__19350),
            .I(N__19347));
    LocalMux I__2522 (
            .O(N__19347),
            .I(\b2v_inst11.count_off_0_11 ));
    InMux I__2521 (
            .O(N__19344),
            .I(N__19341));
    LocalMux I__2520 (
            .O(N__19341),
            .I(\b2v_inst11.count_off_0_10 ));
    InMux I__2519 (
            .O(N__19338),
            .I(N__19335));
    LocalMux I__2518 (
            .O(N__19335),
            .I(\b2v_inst11.count_off_0_12 ));
    InMux I__2517 (
            .O(N__19332),
            .I(N__19329));
    LocalMux I__2516 (
            .O(N__19329),
            .I(N__19326));
    Span4Mux_v I__2515 (
            .O(N__19326),
            .I(N__19322));
    InMux I__2514 (
            .O(N__19325),
            .I(N__19319));
    Odrv4 I__2513 (
            .O(N__19322),
            .I(\b2v_inst16.count_rst_7 ));
    LocalMux I__2512 (
            .O(N__19319),
            .I(\b2v_inst16.count_rst_7 ));
    InMux I__2511 (
            .O(N__19314),
            .I(N__19311));
    LocalMux I__2510 (
            .O(N__19311),
            .I(N__19308));
    Odrv4 I__2509 (
            .O(N__19308),
            .I(\b2v_inst16.count_4_2 ));
    InMux I__2508 (
            .O(N__19305),
            .I(N__19301));
    InMux I__2507 (
            .O(N__19304),
            .I(N__19298));
    LocalMux I__2506 (
            .O(N__19301),
            .I(N__19293));
    LocalMux I__2505 (
            .O(N__19298),
            .I(N__19293));
    Span4Mux_h I__2504 (
            .O(N__19293),
            .I(N__19290));
    Odrv4 I__2503 (
            .O(N__19290),
            .I(\b2v_inst16.count_rst_11 ));
    InMux I__2502 (
            .O(N__19287),
            .I(N__19284));
    LocalMux I__2501 (
            .O(N__19284),
            .I(N__19281));
    Odrv12 I__2500 (
            .O(N__19281),
            .I(\b2v_inst16.count_4_6 ));
    InMux I__2499 (
            .O(N__19278),
            .I(N__19266));
    CEMux I__2498 (
            .O(N__19277),
            .I(N__19266));
    CEMux I__2497 (
            .O(N__19276),
            .I(N__19263));
    InMux I__2496 (
            .O(N__19275),
            .I(N__19258));
    CEMux I__2495 (
            .O(N__19274),
            .I(N__19258));
    CEMux I__2494 (
            .O(N__19273),
            .I(N__19253));
    InMux I__2493 (
            .O(N__19272),
            .I(N__19248));
    InMux I__2492 (
            .O(N__19271),
            .I(N__19248));
    LocalMux I__2491 (
            .O(N__19266),
            .I(N__19237));
    LocalMux I__2490 (
            .O(N__19263),
            .I(N__19234));
    LocalMux I__2489 (
            .O(N__19258),
            .I(N__19231));
    CEMux I__2488 (
            .O(N__19257),
            .I(N__19228));
    CEMux I__2487 (
            .O(N__19256),
            .I(N__19225));
    LocalMux I__2486 (
            .O(N__19253),
            .I(N__19218));
    LocalMux I__2485 (
            .O(N__19248),
            .I(N__19215));
    InMux I__2484 (
            .O(N__19247),
            .I(N__19210));
    InMux I__2483 (
            .O(N__19246),
            .I(N__19210));
    InMux I__2482 (
            .O(N__19245),
            .I(N__19207));
    InMux I__2481 (
            .O(N__19244),
            .I(N__19200));
    InMux I__2480 (
            .O(N__19243),
            .I(N__19200));
    InMux I__2479 (
            .O(N__19242),
            .I(N__19200));
    InMux I__2478 (
            .O(N__19241),
            .I(N__19195));
    InMux I__2477 (
            .O(N__19240),
            .I(N__19195));
    Span4Mux_h I__2476 (
            .O(N__19237),
            .I(N__19190));
    Span4Mux_s2_h I__2475 (
            .O(N__19234),
            .I(N__19190));
    Span4Mux_v I__2474 (
            .O(N__19231),
            .I(N__19185));
    LocalMux I__2473 (
            .O(N__19228),
            .I(N__19185));
    LocalMux I__2472 (
            .O(N__19225),
            .I(N__19182));
    InMux I__2471 (
            .O(N__19224),
            .I(N__19179));
    InMux I__2470 (
            .O(N__19223),
            .I(N__19172));
    InMux I__2469 (
            .O(N__19222),
            .I(N__19172));
    InMux I__2468 (
            .O(N__19221),
            .I(N__19172));
    Span4Mux_s1_h I__2467 (
            .O(N__19218),
            .I(N__19159));
    Span4Mux_h I__2466 (
            .O(N__19215),
            .I(N__19159));
    LocalMux I__2465 (
            .O(N__19210),
            .I(N__19159));
    LocalMux I__2464 (
            .O(N__19207),
            .I(N__19159));
    LocalMux I__2463 (
            .O(N__19200),
            .I(N__19159));
    LocalMux I__2462 (
            .O(N__19195),
            .I(N__19159));
    Odrv4 I__2461 (
            .O(N__19190),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__2460 (
            .O(N__19185),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__2459 (
            .O(N__19182),
            .I(\b2v_inst16.count_en ));
    LocalMux I__2458 (
            .O(N__19179),
            .I(\b2v_inst16.count_en ));
    LocalMux I__2457 (
            .O(N__19172),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__2456 (
            .O(N__19159),
            .I(\b2v_inst16.count_en ));
    SRMux I__2455 (
            .O(N__19146),
            .I(N__19142));
    SRMux I__2454 (
            .O(N__19145),
            .I(N__19138));
    LocalMux I__2453 (
            .O(N__19142),
            .I(N__19134));
    SRMux I__2452 (
            .O(N__19141),
            .I(N__19131));
    LocalMux I__2451 (
            .O(N__19138),
            .I(N__19127));
    SRMux I__2450 (
            .O(N__19137),
            .I(N__19124));
    Span4Mux_h I__2449 (
            .O(N__19134),
            .I(N__19120));
    LocalMux I__2448 (
            .O(N__19131),
            .I(N__19117));
    SRMux I__2447 (
            .O(N__19130),
            .I(N__19114));
    Span4Mux_v I__2446 (
            .O(N__19127),
            .I(N__19109));
    LocalMux I__2445 (
            .O(N__19124),
            .I(N__19109));
    SRMux I__2444 (
            .O(N__19123),
            .I(N__19106));
    Odrv4 I__2443 (
            .O(N__19120),
            .I(\b2v_inst16.N_3037_i ));
    Odrv4 I__2442 (
            .O(N__19117),
            .I(\b2v_inst16.N_3037_i ));
    LocalMux I__2441 (
            .O(N__19114),
            .I(\b2v_inst16.N_3037_i ));
    Odrv4 I__2440 (
            .O(N__19109),
            .I(\b2v_inst16.N_3037_i ));
    LocalMux I__2439 (
            .O(N__19106),
            .I(\b2v_inst16.N_3037_i ));
    InMux I__2438 (
            .O(N__19095),
            .I(N__19092));
    LocalMux I__2437 (
            .O(N__19092),
            .I(\b2v_inst36.curr_state_0_1 ));
    CascadeMux I__2436 (
            .O(N__19089),
            .I(\b2v_inst36.curr_state_7_1_cascade_ ));
    CascadeMux I__2435 (
            .O(N__19086),
            .I(\b2v_inst36.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__2434 (
            .O(N__19083),
            .I(N__19077));
    CascadeMux I__2433 (
            .O(N__19082),
            .I(N__19074));
    CascadeMux I__2432 (
            .O(N__19081),
            .I(N__19065));
    InMux I__2431 (
            .O(N__19080),
            .I(N__19057));
    InMux I__2430 (
            .O(N__19077),
            .I(N__19054));
    InMux I__2429 (
            .O(N__19074),
            .I(N__19049));
    InMux I__2428 (
            .O(N__19073),
            .I(N__19049));
    InMux I__2427 (
            .O(N__19072),
            .I(N__19044));
    InMux I__2426 (
            .O(N__19071),
            .I(N__19044));
    InMux I__2425 (
            .O(N__19070),
            .I(N__19037));
    InMux I__2424 (
            .O(N__19069),
            .I(N__19037));
    InMux I__2423 (
            .O(N__19068),
            .I(N__19037));
    InMux I__2422 (
            .O(N__19065),
            .I(N__19026));
    InMux I__2421 (
            .O(N__19064),
            .I(N__19026));
    InMux I__2420 (
            .O(N__19063),
            .I(N__19026));
    InMux I__2419 (
            .O(N__19062),
            .I(N__19026));
    InMux I__2418 (
            .O(N__19061),
            .I(N__19026));
    CascadeMux I__2417 (
            .O(N__19060),
            .I(N__19022));
    LocalMux I__2416 (
            .O(N__19057),
            .I(N__19014));
    LocalMux I__2415 (
            .O(N__19054),
            .I(N__19014));
    LocalMux I__2414 (
            .O(N__19049),
            .I(N__19009));
    LocalMux I__2413 (
            .O(N__19044),
            .I(N__19009));
    LocalMux I__2412 (
            .O(N__19037),
            .I(N__19004));
    LocalMux I__2411 (
            .O(N__19026),
            .I(N__19004));
    InMux I__2410 (
            .O(N__19025),
            .I(N__18993));
    InMux I__2409 (
            .O(N__19022),
            .I(N__18993));
    InMux I__2408 (
            .O(N__19021),
            .I(N__18993));
    InMux I__2407 (
            .O(N__19020),
            .I(N__18993));
    InMux I__2406 (
            .O(N__19019),
            .I(N__18993));
    Span4Mux_s1_v I__2405 (
            .O(N__19014),
            .I(N__18988));
    Span4Mux_h I__2404 (
            .O(N__19009),
            .I(N__18988));
    Odrv4 I__2403 (
            .O(N__19004),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__2402 (
            .O(N__18993),
            .I(\b2v_inst36.N_1_i ));
    Odrv4 I__2401 (
            .O(N__18988),
            .I(\b2v_inst36.N_1_i ));
    InMux I__2400 (
            .O(N__18981),
            .I(N__18978));
    LocalMux I__2399 (
            .O(N__18978),
            .I(\b2v_inst36.curr_state_0_0 ));
    CascadeMux I__2398 (
            .O(N__18975),
            .I(\b2v_inst36.curr_state_7_0_cascade_ ));
    CascadeMux I__2397 (
            .O(N__18972),
            .I(N__18969));
    InMux I__2396 (
            .O(N__18969),
            .I(N__18965));
    InMux I__2395 (
            .O(N__18968),
            .I(N__18962));
    LocalMux I__2394 (
            .O(N__18965),
            .I(\b2v_inst200.count_3_5 ));
    LocalMux I__2393 (
            .O(N__18962),
            .I(\b2v_inst200.count_3_5 ));
    CascadeMux I__2392 (
            .O(N__18957),
            .I(N__18953));
    InMux I__2391 (
            .O(N__18956),
            .I(N__18950));
    InMux I__2390 (
            .O(N__18953),
            .I(N__18947));
    LocalMux I__2389 (
            .O(N__18950),
            .I(N__18942));
    LocalMux I__2388 (
            .O(N__18947),
            .I(N__18942));
    Span4Mux_v I__2387 (
            .O(N__18942),
            .I(N__18939));
    Odrv4 I__2386 (
            .O(N__18939),
            .I(\b2v_inst16.countZ0Z_15 ));
    InMux I__2385 (
            .O(N__18936),
            .I(N__18930));
    InMux I__2384 (
            .O(N__18935),
            .I(N__18930));
    LocalMux I__2383 (
            .O(N__18930),
            .I(N__18927));
    Span4Mux_h I__2382 (
            .O(N__18927),
            .I(N__18924));
    Odrv4 I__2381 (
            .O(N__18924),
            .I(\b2v_inst16.count_rst_4 ));
    InMux I__2380 (
            .O(N__18921),
            .I(N__18918));
    LocalMux I__2379 (
            .O(N__18918),
            .I(\b2v_inst16.count_4_15 ));
    InMux I__2378 (
            .O(N__18915),
            .I(N__18912));
    LocalMux I__2377 (
            .O(N__18912),
            .I(N__18908));
    InMux I__2376 (
            .O(N__18911),
            .I(N__18905));
    Span4Mux_v I__2375 (
            .O(N__18908),
            .I(N__18900));
    LocalMux I__2374 (
            .O(N__18905),
            .I(N__18900));
    Span4Mux_h I__2373 (
            .O(N__18900),
            .I(N__18897));
    Odrv4 I__2372 (
            .O(N__18897),
            .I(\b2v_inst16.countZ0Z_13 ));
    InMux I__2371 (
            .O(N__18894),
            .I(N__18888));
    InMux I__2370 (
            .O(N__18893),
            .I(N__18888));
    LocalMux I__2369 (
            .O(N__18888),
            .I(N__18885));
    Span4Mux_v I__2368 (
            .O(N__18885),
            .I(N__18882));
    Sp12to4 I__2367 (
            .O(N__18882),
            .I(N__18879));
    Odrv12 I__2366 (
            .O(N__18879),
            .I(\b2v_inst16.count_rst_2 ));
    InMux I__2365 (
            .O(N__18876),
            .I(N__18873));
    LocalMux I__2364 (
            .O(N__18873),
            .I(\b2v_inst16.count_4_13 ));
    CascadeMux I__2363 (
            .O(N__18870),
            .I(N__18867));
    InMux I__2362 (
            .O(N__18867),
            .I(N__18863));
    InMux I__2361 (
            .O(N__18866),
            .I(N__18860));
    LocalMux I__2360 (
            .O(N__18863),
            .I(N__18857));
    LocalMux I__2359 (
            .O(N__18860),
            .I(N__18854));
    Span4Mux_v I__2358 (
            .O(N__18857),
            .I(N__18851));
    Span4Mux_s3_h I__2357 (
            .O(N__18854),
            .I(N__18848));
    Odrv4 I__2356 (
            .O(N__18851),
            .I(\b2v_inst16.countZ0Z_14 ));
    Odrv4 I__2355 (
            .O(N__18848),
            .I(\b2v_inst16.countZ0Z_14 ));
    InMux I__2354 (
            .O(N__18843),
            .I(N__18837));
    InMux I__2353 (
            .O(N__18842),
            .I(N__18837));
    LocalMux I__2352 (
            .O(N__18837),
            .I(N__18834));
    Span4Mux_v I__2351 (
            .O(N__18834),
            .I(N__18831));
    Odrv4 I__2350 (
            .O(N__18831),
            .I(\b2v_inst16.count_rst_3 ));
    InMux I__2349 (
            .O(N__18828),
            .I(N__18825));
    LocalMux I__2348 (
            .O(N__18825),
            .I(\b2v_inst16.count_4_14 ));
    CascadeMux I__2347 (
            .O(N__18822),
            .I(N__18819));
    InMux I__2346 (
            .O(N__18819),
            .I(N__18813));
    InMux I__2345 (
            .O(N__18818),
            .I(N__18813));
    LocalMux I__2344 (
            .O(N__18813),
            .I(\b2v_inst200.count_3_3 ));
    InMux I__2343 (
            .O(N__18810),
            .I(N__18807));
    LocalMux I__2342 (
            .O(N__18807),
            .I(\b2v_inst200.un25_clk_100khz_2 ));
    CascadeMux I__2341 (
            .O(N__18804),
            .I(N__18801));
    InMux I__2340 (
            .O(N__18801),
            .I(N__18795));
    InMux I__2339 (
            .O(N__18800),
            .I(N__18795));
    LocalMux I__2338 (
            .O(N__18795),
            .I(\b2v_inst200.count_3_13 ));
    InMux I__2337 (
            .O(N__18792),
            .I(N__18789));
    LocalMux I__2336 (
            .O(N__18789),
            .I(\b2v_inst200.un25_clk_100khz_5 ));
    InMux I__2335 (
            .O(N__18786),
            .I(N__18783));
    LocalMux I__2334 (
            .O(N__18783),
            .I(\b2v_inst200.count_3_12 ));
    InMux I__2333 (
            .O(N__18780),
            .I(N__18774));
    InMux I__2332 (
            .O(N__18779),
            .I(N__18774));
    LocalMux I__2331 (
            .O(N__18774),
            .I(\b2v_inst200.count_3_9 ));
    CascadeMux I__2330 (
            .O(N__18771),
            .I(\b2v_inst200.countZ0Z_12_cascade_ ));
    InMux I__2329 (
            .O(N__18768),
            .I(N__18765));
    LocalMux I__2328 (
            .O(N__18765),
            .I(\b2v_inst200.un25_clk_100khz_4 ));
    CascadeMux I__2327 (
            .O(N__18762),
            .I(\b2v_inst200.un25_clk_100khz_1_cascade_ ));
    CascadeMux I__2326 (
            .O(N__18759),
            .I(\b2v_inst200.un2_count_1_axb_1_cascade_ ));
    InMux I__2325 (
            .O(N__18756),
            .I(N__18752));
    InMux I__2324 (
            .O(N__18755),
            .I(N__18749));
    LocalMux I__2323 (
            .O(N__18752),
            .I(\b2v_inst200.count_RNIZ0Z_1 ));
    LocalMux I__2322 (
            .O(N__18749),
            .I(\b2v_inst200.count_RNIZ0Z_1 ));
    InMux I__2321 (
            .O(N__18744),
            .I(N__18738));
    InMux I__2320 (
            .O(N__18743),
            .I(N__18738));
    LocalMux I__2319 (
            .O(N__18738),
            .I(\b2v_inst200.countZ0Z_16 ));
    InMux I__2318 (
            .O(N__18735),
            .I(N__18732));
    LocalMux I__2317 (
            .O(N__18732),
            .I(\b2v_inst200.un25_clk_100khz_0 ));
    CascadeMux I__2316 (
            .O(N__18729),
            .I(N__18726));
    InMux I__2315 (
            .O(N__18726),
            .I(N__18720));
    InMux I__2314 (
            .O(N__18725),
            .I(N__18720));
    LocalMux I__2313 (
            .O(N__18720),
            .I(\b2v_inst200.count_3_1 ));
    CascadeMux I__2312 (
            .O(N__18717),
            .I(\b2v_inst200.un25_clk_100khz_3_cascade_ ));
    InMux I__2311 (
            .O(N__18714),
            .I(\b2v_inst11.mult1_un103_sum_cry_3 ));
    InMux I__2310 (
            .O(N__18711),
            .I(\b2v_inst11.mult1_un103_sum_cry_4 ));
    InMux I__2309 (
            .O(N__18708),
            .I(\b2v_inst11.mult1_un103_sum_cry_5 ));
    InMux I__2308 (
            .O(N__18705),
            .I(\b2v_inst11.mult1_un103_sum_cry_6 ));
    InMux I__2307 (
            .O(N__18702),
            .I(\b2v_inst11.mult1_un103_sum_cry_7 ));
    CascadeMux I__2306 (
            .O(N__18699),
            .I(N__18695));
    CascadeMux I__2305 (
            .O(N__18698),
            .I(N__18691));
    InMux I__2304 (
            .O(N__18695),
            .I(N__18684));
    InMux I__2303 (
            .O(N__18694),
            .I(N__18684));
    InMux I__2302 (
            .O(N__18691),
            .I(N__18684));
    LocalMux I__2301 (
            .O(N__18684),
            .I(\b2v_inst11.mult1_un96_sum_i_0_8 ));
    InMux I__2300 (
            .O(N__18681),
            .I(N__18677));
    InMux I__2299 (
            .O(N__18680),
            .I(N__18674));
    LocalMux I__2298 (
            .O(N__18677),
            .I(\b2v_inst11.N_5862_i ));
    LocalMux I__2297 (
            .O(N__18674),
            .I(\b2v_inst11.N_5862_i ));
    CascadeMux I__2296 (
            .O(N__18669),
            .I(N__18665));
    CascadeMux I__2295 (
            .O(N__18668),
            .I(N__18662));
    InMux I__2294 (
            .O(N__18665),
            .I(N__18659));
    InMux I__2293 (
            .O(N__18662),
            .I(N__18656));
    LocalMux I__2292 (
            .O(N__18659),
            .I(N__18653));
    LocalMux I__2291 (
            .O(N__18656),
            .I(\b2v_inst11.un85_clk_100khz_1_8 ));
    Odrv4 I__2290 (
            .O(N__18653),
            .I(\b2v_inst11.un85_clk_100khz_1_8 ));
    CascadeMux I__2289 (
            .O(N__18648),
            .I(N__18645));
    InMux I__2288 (
            .O(N__18645),
            .I(N__18641));
    InMux I__2287 (
            .O(N__18644),
            .I(N__18638));
    LocalMux I__2286 (
            .O(N__18641),
            .I(\b2v_inst11.N_5863_i ));
    LocalMux I__2285 (
            .O(N__18638),
            .I(\b2v_inst11.N_5863_i ));
    CascadeMux I__2284 (
            .O(N__18633),
            .I(N__18630));
    InMux I__2283 (
            .O(N__18630),
            .I(N__18626));
    InMux I__2282 (
            .O(N__18629),
            .I(N__18623));
    LocalMux I__2281 (
            .O(N__18626),
            .I(N__18620));
    LocalMux I__2280 (
            .O(N__18623),
            .I(\b2v_inst11.un85_clk_100khz_1_9 ));
    Odrv4 I__2279 (
            .O(N__18620),
            .I(\b2v_inst11.un85_clk_100khz_1_9 ));
    CascadeMux I__2278 (
            .O(N__18615),
            .I(N__18612));
    InMux I__2277 (
            .O(N__18612),
            .I(N__18608));
    InMux I__2276 (
            .O(N__18611),
            .I(N__18605));
    LocalMux I__2275 (
            .O(N__18608),
            .I(\b2v_inst11.N_5864_i ));
    LocalMux I__2274 (
            .O(N__18605),
            .I(\b2v_inst11.N_5864_i ));
    CascadeMux I__2273 (
            .O(N__18600),
            .I(N__18596));
    InMux I__2272 (
            .O(N__18599),
            .I(N__18593));
    InMux I__2271 (
            .O(N__18596),
            .I(N__18590));
    LocalMux I__2270 (
            .O(N__18593),
            .I(\b2v_inst11.un85_clk_100khz_1_10 ));
    LocalMux I__2269 (
            .O(N__18590),
            .I(\b2v_inst11.un85_clk_100khz_1_10 ));
    CascadeMux I__2268 (
            .O(N__18585),
            .I(N__18581));
    CascadeMux I__2267 (
            .O(N__18584),
            .I(N__18578));
    InMux I__2266 (
            .O(N__18581),
            .I(N__18575));
    InMux I__2265 (
            .O(N__18578),
            .I(N__18572));
    LocalMux I__2264 (
            .O(N__18575),
            .I(\b2v_inst11.N_5865_i ));
    LocalMux I__2263 (
            .O(N__18572),
            .I(\b2v_inst11.N_5865_i ));
    InMux I__2262 (
            .O(N__18567),
            .I(N__18563));
    InMux I__2261 (
            .O(N__18566),
            .I(N__18560));
    LocalMux I__2260 (
            .O(N__18563),
            .I(N__18557));
    LocalMux I__2259 (
            .O(N__18560),
            .I(\b2v_inst11.un85_clk_100khz_1_11 ));
    Odrv4 I__2258 (
            .O(N__18557),
            .I(\b2v_inst11.un85_clk_100khz_1_11 ));
    CascadeMux I__2257 (
            .O(N__18552),
            .I(N__18548));
    InMux I__2256 (
            .O(N__18551),
            .I(N__18545));
    InMux I__2255 (
            .O(N__18548),
            .I(N__18542));
    LocalMux I__2254 (
            .O(N__18545),
            .I(\b2v_inst11.N_5866_i ));
    LocalMux I__2253 (
            .O(N__18542),
            .I(\b2v_inst11.N_5866_i ));
    CascadeMux I__2252 (
            .O(N__18537),
            .I(N__18534));
    InMux I__2251 (
            .O(N__18534),
            .I(N__18530));
    InMux I__2250 (
            .O(N__18533),
            .I(N__18527));
    LocalMux I__2249 (
            .O(N__18530),
            .I(\b2v_inst11.un85_clk_100khz_1_12 ));
    LocalMux I__2248 (
            .O(N__18527),
            .I(\b2v_inst11.un85_clk_100khz_1_12 ));
    CascadeMux I__2247 (
            .O(N__18522),
            .I(N__18518));
    CascadeMux I__2246 (
            .O(N__18521),
            .I(N__18515));
    InMux I__2245 (
            .O(N__18518),
            .I(N__18512));
    InMux I__2244 (
            .O(N__18515),
            .I(N__18509));
    LocalMux I__2243 (
            .O(N__18512),
            .I(\b2v_inst11.N_5867_i ));
    LocalMux I__2242 (
            .O(N__18509),
            .I(\b2v_inst11.N_5867_i ));
    InMux I__2241 (
            .O(N__18504),
            .I(N__18500));
    InMux I__2240 (
            .O(N__18503),
            .I(N__18497));
    LocalMux I__2239 (
            .O(N__18500),
            .I(\b2v_inst11.un85_clk_100khz_1_13 ));
    LocalMux I__2238 (
            .O(N__18497),
            .I(\b2v_inst11.un85_clk_100khz_1_13 ));
    InMux I__2237 (
            .O(N__18492),
            .I(\b2v_inst11.un85_clk_100khz1 ));
    InMux I__2236 (
            .O(N__18489),
            .I(\b2v_inst11.mult1_un103_sum_cry_2 ));
    InMux I__2235 (
            .O(N__18486),
            .I(N__18482));
    InMux I__2234 (
            .O(N__18485),
            .I(N__18479));
    LocalMux I__2233 (
            .O(N__18482),
            .I(\b2v_inst11.N_5855_i ));
    LocalMux I__2232 (
            .O(N__18479),
            .I(\b2v_inst11.N_5855_i ));
    CascadeMux I__2231 (
            .O(N__18474),
            .I(N__18470));
    CascadeMux I__2230 (
            .O(N__18473),
            .I(N__18467));
    InMux I__2229 (
            .O(N__18470),
            .I(N__18464));
    InMux I__2228 (
            .O(N__18467),
            .I(N__18461));
    LocalMux I__2227 (
            .O(N__18464),
            .I(\b2v_inst11.un85_clk_100khz_0_1 ));
    LocalMux I__2226 (
            .O(N__18461),
            .I(\b2v_inst11.un85_clk_100khz_0_1 ));
    CascadeMux I__2225 (
            .O(N__18456),
            .I(N__18452));
    InMux I__2224 (
            .O(N__18455),
            .I(N__18449));
    InMux I__2223 (
            .O(N__18452),
            .I(N__18446));
    LocalMux I__2222 (
            .O(N__18449),
            .I(\b2v_inst11.N_5856_i ));
    LocalMux I__2221 (
            .O(N__18446),
            .I(\b2v_inst11.N_5856_i ));
    CascadeMux I__2220 (
            .O(N__18441),
            .I(N__18438));
    InMux I__2219 (
            .O(N__18438),
            .I(N__18434));
    InMux I__2218 (
            .O(N__18437),
            .I(N__18431));
    LocalMux I__2217 (
            .O(N__18434),
            .I(\b2v_inst11.un85_clk_100khz_0_2 ));
    LocalMux I__2216 (
            .O(N__18431),
            .I(\b2v_inst11.un85_clk_100khz_0_2 ));
    InMux I__2215 (
            .O(N__18426),
            .I(N__18422));
    InMux I__2214 (
            .O(N__18425),
            .I(N__18419));
    LocalMux I__2213 (
            .O(N__18422),
            .I(\b2v_inst11.N_5857_i ));
    LocalMux I__2212 (
            .O(N__18419),
            .I(\b2v_inst11.N_5857_i ));
    CascadeMux I__2211 (
            .O(N__18414),
            .I(N__18410));
    CascadeMux I__2210 (
            .O(N__18413),
            .I(N__18407));
    InMux I__2209 (
            .O(N__18410),
            .I(N__18404));
    InMux I__2208 (
            .O(N__18407),
            .I(N__18401));
    LocalMux I__2207 (
            .O(N__18404),
            .I(N__18398));
    LocalMux I__2206 (
            .O(N__18401),
            .I(\b2v_inst11.un85_clk_100khz_0_3 ));
    Odrv4 I__2205 (
            .O(N__18398),
            .I(\b2v_inst11.un85_clk_100khz_0_3 ));
    InMux I__2204 (
            .O(N__18393),
            .I(N__18389));
    InMux I__2203 (
            .O(N__18392),
            .I(N__18386));
    LocalMux I__2202 (
            .O(N__18389),
            .I(\b2v_inst11.N_5858_i ));
    LocalMux I__2201 (
            .O(N__18386),
            .I(\b2v_inst11.N_5858_i ));
    CascadeMux I__2200 (
            .O(N__18381),
            .I(N__18377));
    CascadeMux I__2199 (
            .O(N__18380),
            .I(N__18374));
    InMux I__2198 (
            .O(N__18377),
            .I(N__18371));
    InMux I__2197 (
            .O(N__18374),
            .I(N__18368));
    LocalMux I__2196 (
            .O(N__18371),
            .I(\b2v_inst11.un85_clk_100khz_0_4 ));
    LocalMux I__2195 (
            .O(N__18368),
            .I(\b2v_inst11.un85_clk_100khz_0_4 ));
    CascadeMux I__2194 (
            .O(N__18363),
            .I(N__18360));
    InMux I__2193 (
            .O(N__18360),
            .I(N__18356));
    InMux I__2192 (
            .O(N__18359),
            .I(N__18353));
    LocalMux I__2191 (
            .O(N__18356),
            .I(\b2v_inst11.N_5859_i ));
    LocalMux I__2190 (
            .O(N__18353),
            .I(\b2v_inst11.N_5859_i ));
    CascadeMux I__2189 (
            .O(N__18348),
            .I(N__18344));
    InMux I__2188 (
            .O(N__18347),
            .I(N__18341));
    InMux I__2187 (
            .O(N__18344),
            .I(N__18338));
    LocalMux I__2186 (
            .O(N__18341),
            .I(\b2v_inst11.un85_clk_100khz_0_5 ));
    LocalMux I__2185 (
            .O(N__18338),
            .I(\b2v_inst11.un85_clk_100khz_0_5 ));
    InMux I__2184 (
            .O(N__18333),
            .I(N__18329));
    InMux I__2183 (
            .O(N__18332),
            .I(N__18326));
    LocalMux I__2182 (
            .O(N__18329),
            .I(\b2v_inst11.N_5860_i ));
    LocalMux I__2181 (
            .O(N__18326),
            .I(\b2v_inst11.N_5860_i ));
    CascadeMux I__2180 (
            .O(N__18321),
            .I(N__18317));
    CascadeMux I__2179 (
            .O(N__18320),
            .I(N__18314));
    InMux I__2178 (
            .O(N__18317),
            .I(N__18311));
    InMux I__2177 (
            .O(N__18314),
            .I(N__18308));
    LocalMux I__2176 (
            .O(N__18311),
            .I(\b2v_inst11.un85_clk_100khz_0_6 ));
    LocalMux I__2175 (
            .O(N__18308),
            .I(\b2v_inst11.un85_clk_100khz_0_6 ));
    InMux I__2174 (
            .O(N__18303),
            .I(N__18299));
    InMux I__2173 (
            .O(N__18302),
            .I(N__18296));
    LocalMux I__2172 (
            .O(N__18299),
            .I(\b2v_inst11.N_5861_i ));
    LocalMux I__2171 (
            .O(N__18296),
            .I(\b2v_inst11.N_5861_i ));
    CascadeMux I__2170 (
            .O(N__18291),
            .I(N__18287));
    CascadeMux I__2169 (
            .O(N__18290),
            .I(N__18284));
    InMux I__2168 (
            .O(N__18287),
            .I(N__18281));
    InMux I__2167 (
            .O(N__18284),
            .I(N__18278));
    LocalMux I__2166 (
            .O(N__18281),
            .I(N__18275));
    LocalMux I__2165 (
            .O(N__18278),
            .I(\b2v_inst11.un85_clk_100khz_0_7 ));
    Odrv4 I__2164 (
            .O(N__18275),
            .I(\b2v_inst11.un85_clk_100khz_0_7 ));
    InMux I__2163 (
            .O(N__18270),
            .I(N__18266));
    InMux I__2162 (
            .O(N__18269),
            .I(N__18263));
    LocalMux I__2161 (
            .O(N__18266),
            .I(N__18259));
    LocalMux I__2160 (
            .O(N__18263),
            .I(N__18256));
    InMux I__2159 (
            .O(N__18262),
            .I(N__18253));
    Odrv4 I__2158 (
            .O(N__18259),
            .I(\b2v_inst11.countZ0Z_2 ));
    Odrv4 I__2157 (
            .O(N__18256),
            .I(\b2v_inst11.countZ0Z_2 ));
    LocalMux I__2156 (
            .O(N__18253),
            .I(\b2v_inst11.countZ0Z_2 ));
    InMux I__2155 (
            .O(N__18246),
            .I(N__18241));
    CascadeMux I__2154 (
            .O(N__18245),
            .I(N__18238));
    InMux I__2153 (
            .O(N__18244),
            .I(N__18235));
    LocalMux I__2152 (
            .O(N__18241),
            .I(N__18232));
    InMux I__2151 (
            .O(N__18238),
            .I(N__18229));
    LocalMux I__2150 (
            .O(N__18235),
            .I(\b2v_inst11.countZ0Z_3 ));
    Odrv4 I__2149 (
            .O(N__18232),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__2148 (
            .O(N__18229),
            .I(\b2v_inst11.countZ0Z_3 ));
    InMux I__2147 (
            .O(N__18222),
            .I(N__18217));
    CascadeMux I__2146 (
            .O(N__18221),
            .I(N__18214));
    InMux I__2145 (
            .O(N__18220),
            .I(N__18211));
    LocalMux I__2144 (
            .O(N__18217),
            .I(N__18208));
    InMux I__2143 (
            .O(N__18214),
            .I(N__18205));
    LocalMux I__2142 (
            .O(N__18211),
            .I(\b2v_inst11.countZ0Z_4 ));
    Odrv4 I__2141 (
            .O(N__18208),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__2140 (
            .O(N__18205),
            .I(\b2v_inst11.countZ0Z_4 ));
    InMux I__2139 (
            .O(N__18198),
            .I(N__18193));
    InMux I__2138 (
            .O(N__18197),
            .I(N__18190));
    CascadeMux I__2137 (
            .O(N__18196),
            .I(N__18187));
    LocalMux I__2136 (
            .O(N__18193),
            .I(N__18184));
    LocalMux I__2135 (
            .O(N__18190),
            .I(N__18181));
    InMux I__2134 (
            .O(N__18187),
            .I(N__18178));
    Span4Mux_v I__2133 (
            .O(N__18184),
            .I(N__18175));
    Span4Mux_v I__2132 (
            .O(N__18181),
            .I(N__18170));
    LocalMux I__2131 (
            .O(N__18178),
            .I(N__18170));
    Odrv4 I__2130 (
            .O(N__18175),
            .I(\b2v_inst11.countZ0Z_7 ));
    Odrv4 I__2129 (
            .O(N__18170),
            .I(\b2v_inst11.countZ0Z_7 ));
    CascadeMux I__2128 (
            .O(N__18165),
            .I(N__18162));
    InMux I__2127 (
            .O(N__18162),
            .I(N__18157));
    InMux I__2126 (
            .O(N__18161),
            .I(N__18154));
    InMux I__2125 (
            .O(N__18160),
            .I(N__18151));
    LocalMux I__2124 (
            .O(N__18157),
            .I(N__18148));
    LocalMux I__2123 (
            .O(N__18154),
            .I(\b2v_inst11.countZ0Z_6 ));
    LocalMux I__2122 (
            .O(N__18151),
            .I(\b2v_inst11.countZ0Z_6 ));
    Odrv4 I__2121 (
            .O(N__18148),
            .I(\b2v_inst11.countZ0Z_6 ));
    CascadeMux I__2120 (
            .O(N__18141),
            .I(\b2v_inst11.un79_clk_100khzlt6_cascade_ ));
    CascadeMux I__2119 (
            .O(N__18138),
            .I(N__18134));
    InMux I__2118 (
            .O(N__18137),
            .I(N__18131));
    InMux I__2117 (
            .O(N__18134),
            .I(N__18127));
    LocalMux I__2116 (
            .O(N__18131),
            .I(N__18124));
    InMux I__2115 (
            .O(N__18130),
            .I(N__18121));
    LocalMux I__2114 (
            .O(N__18127),
            .I(N__18118));
    Odrv4 I__2113 (
            .O(N__18124),
            .I(\b2v_inst11.countZ0Z_5 ));
    LocalMux I__2112 (
            .O(N__18121),
            .I(\b2v_inst11.countZ0Z_5 ));
    Odrv4 I__2111 (
            .O(N__18118),
            .I(\b2v_inst11.countZ0Z_5 ));
    InMux I__2110 (
            .O(N__18111),
            .I(N__18107));
    InMux I__2109 (
            .O(N__18110),
            .I(N__18103));
    LocalMux I__2108 (
            .O(N__18107),
            .I(N__18100));
    CascadeMux I__2107 (
            .O(N__18106),
            .I(N__18097));
    LocalMux I__2106 (
            .O(N__18103),
            .I(N__18094));
    Span4Mux_s2_v I__2105 (
            .O(N__18100),
            .I(N__18091));
    InMux I__2104 (
            .O(N__18097),
            .I(N__18088));
    Odrv12 I__2103 (
            .O(N__18094),
            .I(\b2v_inst11.countZ0Z_10 ));
    Odrv4 I__2102 (
            .O(N__18091),
            .I(\b2v_inst11.countZ0Z_10 ));
    LocalMux I__2101 (
            .O(N__18088),
            .I(\b2v_inst11.countZ0Z_10 ));
    InMux I__2100 (
            .O(N__18081),
            .I(N__18078));
    LocalMux I__2099 (
            .O(N__18078),
            .I(N__18073));
    CascadeMux I__2098 (
            .O(N__18077),
            .I(N__18070));
    InMux I__2097 (
            .O(N__18076),
            .I(N__18067));
    Span4Mux_s2_v I__2096 (
            .O(N__18073),
            .I(N__18064));
    InMux I__2095 (
            .O(N__18070),
            .I(N__18061));
    LocalMux I__2094 (
            .O(N__18067),
            .I(\b2v_inst11.countZ0Z_12 ));
    Odrv4 I__2093 (
            .O(N__18064),
            .I(\b2v_inst11.countZ0Z_12 ));
    LocalMux I__2092 (
            .O(N__18061),
            .I(\b2v_inst11.countZ0Z_12 ));
    CascadeMux I__2091 (
            .O(N__18054),
            .I(N__18050));
    InMux I__2090 (
            .O(N__18053),
            .I(N__18047));
    InMux I__2089 (
            .O(N__18050),
            .I(N__18043));
    LocalMux I__2088 (
            .O(N__18047),
            .I(N__18040));
    CascadeMux I__2087 (
            .O(N__18046),
            .I(N__18037));
    LocalMux I__2086 (
            .O(N__18043),
            .I(N__18032));
    Span4Mux_s2_v I__2085 (
            .O(N__18040),
            .I(N__18032));
    InMux I__2084 (
            .O(N__18037),
            .I(N__18029));
    Odrv4 I__2083 (
            .O(N__18032),
            .I(\b2v_inst11.countZ0Z_11 ));
    LocalMux I__2082 (
            .O(N__18029),
            .I(\b2v_inst11.countZ0Z_11 ));
    InMux I__2081 (
            .O(N__18024),
            .I(N__18019));
    InMux I__2080 (
            .O(N__18023),
            .I(N__18016));
    CascadeMux I__2079 (
            .O(N__18022),
            .I(N__18013));
    LocalMux I__2078 (
            .O(N__18019),
            .I(N__18008));
    LocalMux I__2077 (
            .O(N__18016),
            .I(N__18008));
    InMux I__2076 (
            .O(N__18013),
            .I(N__18005));
    Odrv4 I__2075 (
            .O(N__18008),
            .I(\b2v_inst11.countZ0Z_13 ));
    LocalMux I__2074 (
            .O(N__18005),
            .I(\b2v_inst11.countZ0Z_13 ));
    InMux I__2073 (
            .O(N__18000),
            .I(N__17995));
    CascadeMux I__2072 (
            .O(N__17999),
            .I(N__17992));
    InMux I__2071 (
            .O(N__17998),
            .I(N__17989));
    LocalMux I__2070 (
            .O(N__17995),
            .I(N__17986));
    InMux I__2069 (
            .O(N__17992),
            .I(N__17983));
    LocalMux I__2068 (
            .O(N__17989),
            .I(\b2v_inst11.countZ0Z_14 ));
    Odrv4 I__2067 (
            .O(N__17986),
            .I(\b2v_inst11.countZ0Z_14 ));
    LocalMux I__2066 (
            .O(N__17983),
            .I(\b2v_inst11.countZ0Z_14 ));
    CascadeMux I__2065 (
            .O(N__17976),
            .I(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ));
    InMux I__2064 (
            .O(N__17973),
            .I(N__17968));
    InMux I__2063 (
            .O(N__17972),
            .I(N__17965));
    InMux I__2062 (
            .O(N__17971),
            .I(N__17962));
    LocalMux I__2061 (
            .O(N__17968),
            .I(N__17959));
    LocalMux I__2060 (
            .O(N__17965),
            .I(\b2v_inst11.countZ0Z_15 ));
    LocalMux I__2059 (
            .O(N__17962),
            .I(\b2v_inst11.countZ0Z_15 ));
    Odrv4 I__2058 (
            .O(N__17959),
            .I(\b2v_inst11.countZ0Z_15 ));
    InMux I__2057 (
            .O(N__17952),
            .I(N__17949));
    LocalMux I__2056 (
            .O(N__17949),
            .I(\b2v_inst11.un79_clk_100khzlto15_3 ));
    InMux I__2055 (
            .O(N__17946),
            .I(N__17942));
    InMux I__2054 (
            .O(N__17945),
            .I(N__17938));
    LocalMux I__2053 (
            .O(N__17942),
            .I(N__17935));
    CascadeMux I__2052 (
            .O(N__17941),
            .I(N__17932));
    LocalMux I__2051 (
            .O(N__17938),
            .I(N__17927));
    Span4Mux_s3_v I__2050 (
            .O(N__17935),
            .I(N__17927));
    InMux I__2049 (
            .O(N__17932),
            .I(N__17924));
    Odrv4 I__2048 (
            .O(N__17927),
            .I(\b2v_inst11.countZ0Z_8 ));
    LocalMux I__2047 (
            .O(N__17924),
            .I(\b2v_inst11.countZ0Z_8 ));
    CascadeMux I__2046 (
            .O(N__17919),
            .I(\b2v_inst11.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__2045 (
            .O(N__17916),
            .I(N__17912));
    InMux I__2044 (
            .O(N__17915),
            .I(N__17908));
    LocalMux I__2043 (
            .O(N__17912),
            .I(N__17905));
    CascadeMux I__2042 (
            .O(N__17911),
            .I(N__17902));
    LocalMux I__2041 (
            .O(N__17908),
            .I(N__17899));
    Span4Mux_s3_v I__2040 (
            .O(N__17905),
            .I(N__17896));
    InMux I__2039 (
            .O(N__17902),
            .I(N__17893));
    Odrv4 I__2038 (
            .O(N__17899),
            .I(\b2v_inst11.countZ0Z_9 ));
    Odrv4 I__2037 (
            .O(N__17896),
            .I(\b2v_inst11.countZ0Z_9 ));
    LocalMux I__2036 (
            .O(N__17893),
            .I(\b2v_inst11.countZ0Z_9 ));
    CascadeMux I__2035 (
            .O(N__17886),
            .I(N__17881));
    InMux I__2034 (
            .O(N__17885),
            .I(N__17871));
    InMux I__2033 (
            .O(N__17884),
            .I(N__17871));
    InMux I__2032 (
            .O(N__17881),
            .I(N__17871));
    InMux I__2031 (
            .O(N__17880),
            .I(N__17871));
    LocalMux I__2030 (
            .O(N__17871),
            .I(N__17868));
    Odrv12 I__2029 (
            .O(N__17868),
            .I(\b2v_inst11.count_RNIZ0Z_8 ));
    InMux I__2028 (
            .O(N__17865),
            .I(N__17861));
    CascadeMux I__2027 (
            .O(N__17864),
            .I(N__17856));
    LocalMux I__2026 (
            .O(N__17861),
            .I(N__17851));
    InMux I__2025 (
            .O(N__17860),
            .I(N__17848));
    InMux I__2024 (
            .O(N__17859),
            .I(N__17839));
    InMux I__2023 (
            .O(N__17856),
            .I(N__17839));
    InMux I__2022 (
            .O(N__17855),
            .I(N__17839));
    InMux I__2021 (
            .O(N__17854),
            .I(N__17839));
    Span4Mux_v I__2020 (
            .O(N__17851),
            .I(N__17836));
    LocalMux I__2019 (
            .O(N__17848),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    LocalMux I__2018 (
            .O(N__17839),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    Odrv4 I__2017 (
            .O(N__17836),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    CascadeMux I__2016 (
            .O(N__17829),
            .I(\b2v_inst11.count_RNIZ0Z_8_cascade_ ));
    InMux I__2015 (
            .O(N__17826),
            .I(N__17823));
    LocalMux I__2014 (
            .O(N__17823),
            .I(N__17820));
    Odrv12 I__2013 (
            .O(N__17820),
            .I(\b2v_inst11.curr_state_3_i_m2_0_rep1_1 ));
    InMux I__2012 (
            .O(N__17817),
            .I(N__17813));
    InMux I__2011 (
            .O(N__17816),
            .I(N__17810));
    LocalMux I__2010 (
            .O(N__17813),
            .I(\b2v_inst11.N_5853_i ));
    LocalMux I__2009 (
            .O(N__17810),
            .I(\b2v_inst11.N_5853_i ));
    CascadeMux I__2008 (
            .O(N__17805),
            .I(N__17801));
    CascadeMux I__2007 (
            .O(N__17804),
            .I(N__17798));
    InMux I__2006 (
            .O(N__17801),
            .I(N__17795));
    InMux I__2005 (
            .O(N__17798),
            .I(N__17792));
    LocalMux I__2004 (
            .O(N__17795),
            .I(\b2v_inst11.un85_clk_100khz_0 ));
    LocalMux I__2003 (
            .O(N__17792),
            .I(\b2v_inst11.un85_clk_100khz_0 ));
    InMux I__2002 (
            .O(N__17787),
            .I(N__17783));
    InMux I__2001 (
            .O(N__17786),
            .I(N__17780));
    LocalMux I__2000 (
            .O(N__17783),
            .I(\b2v_inst11.N_5854_i ));
    LocalMux I__1999 (
            .O(N__17780),
            .I(\b2v_inst11.N_5854_i ));
    CascadeMux I__1998 (
            .O(N__17775),
            .I(N__17771));
    CascadeMux I__1997 (
            .O(N__17774),
            .I(N__17768));
    InMux I__1996 (
            .O(N__17771),
            .I(N__17765));
    InMux I__1995 (
            .O(N__17768),
            .I(N__17762));
    LocalMux I__1994 (
            .O(N__17765),
            .I(N__17759));
    LocalMux I__1993 (
            .O(N__17762),
            .I(\b2v_inst11.un85_clk_100khz_0_0 ));
    Odrv4 I__1992 (
            .O(N__17759),
            .I(\b2v_inst11.un85_clk_100khz_0_0 ));
    CascadeMux I__1991 (
            .O(N__17754),
            .I(N__17750));
    InMux I__1990 (
            .O(N__17753),
            .I(N__17745));
    InMux I__1989 (
            .O(N__17750),
            .I(N__17745));
    LocalMux I__1988 (
            .O(N__17745),
            .I(\b2v_inst11.count_1_2 ));
    InMux I__1987 (
            .O(N__17742),
            .I(N__17739));
    LocalMux I__1986 (
            .O(N__17739),
            .I(\b2v_inst11.count_0_2 ));
    CascadeMux I__1985 (
            .O(N__17736),
            .I(N__17733));
    InMux I__1984 (
            .O(N__17733),
            .I(N__17727));
    InMux I__1983 (
            .O(N__17732),
            .I(N__17727));
    LocalMux I__1982 (
            .O(N__17727),
            .I(\b2v_inst11.count_1_12 ));
    InMux I__1981 (
            .O(N__17724),
            .I(N__17721));
    LocalMux I__1980 (
            .O(N__17721),
            .I(\b2v_inst11.count_0_12 ));
    InMux I__1979 (
            .O(N__17718),
            .I(N__17712));
    InMux I__1978 (
            .O(N__17717),
            .I(N__17712));
    LocalMux I__1977 (
            .O(N__17712),
            .I(\b2v_inst11.count_1_3 ));
    CascadeMux I__1976 (
            .O(N__17709),
            .I(N__17706));
    InMux I__1975 (
            .O(N__17706),
            .I(N__17703));
    LocalMux I__1974 (
            .O(N__17703),
            .I(\b2v_inst11.count_0_3 ));
    CascadeMux I__1973 (
            .O(N__17700),
            .I(N__17697));
    InMux I__1972 (
            .O(N__17697),
            .I(N__17691));
    InMux I__1971 (
            .O(N__17696),
            .I(N__17691));
    LocalMux I__1970 (
            .O(N__17691),
            .I(\b2v_inst11.count_1_13 ));
    InMux I__1969 (
            .O(N__17688),
            .I(N__17685));
    LocalMux I__1968 (
            .O(N__17685),
            .I(\b2v_inst11.count_0_13 ));
    InMux I__1967 (
            .O(N__17682),
            .I(N__17676));
    InMux I__1966 (
            .O(N__17681),
            .I(N__17676));
    LocalMux I__1965 (
            .O(N__17676),
            .I(\b2v_inst11.count_1_4 ));
    InMux I__1964 (
            .O(N__17673),
            .I(N__17670));
    LocalMux I__1963 (
            .O(N__17670),
            .I(\b2v_inst11.count_0_4 ));
    InMux I__1962 (
            .O(N__17667),
            .I(N__17664));
    LocalMux I__1961 (
            .O(N__17664),
            .I(N__17658));
    CascadeMux I__1960 (
            .O(N__17663),
            .I(N__17655));
    InMux I__1959 (
            .O(N__17662),
            .I(N__17650));
    InMux I__1958 (
            .O(N__17661),
            .I(N__17650));
    Span4Mux_s3_v I__1957 (
            .O(N__17658),
            .I(N__17647));
    InMux I__1956 (
            .O(N__17655),
            .I(N__17644));
    LocalMux I__1955 (
            .O(N__17650),
            .I(\b2v_inst11.countZ0Z_1 ));
    Odrv4 I__1954 (
            .O(N__17647),
            .I(\b2v_inst11.countZ0Z_1 ));
    LocalMux I__1953 (
            .O(N__17644),
            .I(\b2v_inst11.countZ0Z_1 ));
    InMux I__1952 (
            .O(N__17637),
            .I(N__17634));
    LocalMux I__1951 (
            .O(N__17634),
            .I(\b2v_inst11.count_0_1 ));
    InMux I__1950 (
            .O(N__17631),
            .I(N__17628));
    LocalMux I__1949 (
            .O(N__17628),
            .I(N__17625));
    Odrv4 I__1948 (
            .O(N__17625),
            .I(\b2v_inst11.count_0_8 ));
    InMux I__1947 (
            .O(N__17622),
            .I(N__17618));
    InMux I__1946 (
            .O(N__17621),
            .I(N__17615));
    LocalMux I__1945 (
            .O(N__17618),
            .I(\b2v_inst11.count_1_8 ));
    LocalMux I__1944 (
            .O(N__17615),
            .I(\b2v_inst11.count_1_8 ));
    CascadeMux I__1943 (
            .O(N__17610),
            .I(N__17607));
    InMux I__1942 (
            .O(N__17607),
            .I(N__17601));
    InMux I__1941 (
            .O(N__17606),
            .I(N__17601));
    LocalMux I__1940 (
            .O(N__17601),
            .I(\b2v_inst11.count_1_9 ));
    InMux I__1939 (
            .O(N__17598),
            .I(N__17595));
    LocalMux I__1938 (
            .O(N__17595),
            .I(\b2v_inst11.count_0_9 ));
    CascadeMux I__1937 (
            .O(N__17592),
            .I(N__17589));
    InMux I__1936 (
            .O(N__17589),
            .I(N__17583));
    InMux I__1935 (
            .O(N__17588),
            .I(N__17583));
    LocalMux I__1934 (
            .O(N__17583),
            .I(\b2v_inst11.count_1_10 ));
    InMux I__1933 (
            .O(N__17580),
            .I(N__17577));
    LocalMux I__1932 (
            .O(N__17577),
            .I(\b2v_inst11.count_0_10 ));
    CascadeMux I__1931 (
            .O(N__17574),
            .I(N__17571));
    InMux I__1930 (
            .O(N__17571),
            .I(N__17565));
    InMux I__1929 (
            .O(N__17570),
            .I(N__17565));
    LocalMux I__1928 (
            .O(N__17565),
            .I(\b2v_inst11.count_1_11 ));
    InMux I__1927 (
            .O(N__17562),
            .I(N__17559));
    LocalMux I__1926 (
            .O(N__17559),
            .I(\b2v_inst11.count_0_11 ));
    InMux I__1925 (
            .O(N__17556),
            .I(N__17553));
    LocalMux I__1924 (
            .O(N__17553),
            .I(\b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJZ0Z62 ));
    InMux I__1923 (
            .O(N__17550),
            .I(N__17547));
    LocalMux I__1922 (
            .O(N__17547),
            .I(\b2v_inst11.curr_state_4_0 ));
    InMux I__1921 (
            .O(N__17544),
            .I(N__17541));
    LocalMux I__1920 (
            .O(N__17541),
            .I(\b2v_inst11.count_0_0 ));
    CascadeMux I__1919 (
            .O(N__17538),
            .I(\b2v_inst11.countZ0Z_0_cascade_ ));
    CascadeMux I__1918 (
            .O(N__17535),
            .I(\b2v_inst11.count_1_1_cascade_ ));
    CascadeMux I__1917 (
            .O(N__17532),
            .I(CONSTANT_ONE_NET_cascade_));
    InMux I__1916 (
            .O(N__17529),
            .I(N__17526));
    LocalMux I__1915 (
            .O(N__17526),
            .I(N__17522));
    InMux I__1914 (
            .O(N__17525),
            .I(N__17519));
    Span4Mux_v I__1913 (
            .O(N__17522),
            .I(N__17516));
    LocalMux I__1912 (
            .O(N__17519),
            .I(\b2v_inst11.N_5852_i ));
    Odrv4 I__1911 (
            .O(N__17516),
            .I(\b2v_inst11.N_5852_i ));
    InMux I__1910 (
            .O(N__17511),
            .I(N__17505));
    InMux I__1909 (
            .O(N__17510),
            .I(N__17505));
    LocalMux I__1908 (
            .O(N__17505),
            .I(\b2v_inst16.un4_count_1_cry_8_THRU_CO ));
    CascadeMux I__1907 (
            .O(N__17502),
            .I(\b2v_inst16.countZ0Z_9_cascade_ ));
    CascadeMux I__1906 (
            .O(N__17499),
            .I(N__17495));
    InMux I__1905 (
            .O(N__17498),
            .I(N__17480));
    InMux I__1904 (
            .O(N__17495),
            .I(N__17480));
    InMux I__1903 (
            .O(N__17494),
            .I(N__17480));
    InMux I__1902 (
            .O(N__17493),
            .I(N__17464));
    InMux I__1901 (
            .O(N__17492),
            .I(N__17464));
    InMux I__1900 (
            .O(N__17491),
            .I(N__17464));
    InMux I__1899 (
            .O(N__17490),
            .I(N__17464));
    InMux I__1898 (
            .O(N__17489),
            .I(N__17464));
    InMux I__1897 (
            .O(N__17488),
            .I(N__17459));
    InMux I__1896 (
            .O(N__17487),
            .I(N__17459));
    LocalMux I__1895 (
            .O(N__17480),
            .I(N__17456));
    InMux I__1894 (
            .O(N__17479),
            .I(N__17445));
    InMux I__1893 (
            .O(N__17478),
            .I(N__17445));
    InMux I__1892 (
            .O(N__17477),
            .I(N__17445));
    InMux I__1891 (
            .O(N__17476),
            .I(N__17445));
    InMux I__1890 (
            .O(N__17475),
            .I(N__17445));
    LocalMux I__1889 (
            .O(N__17464),
            .I(N__17440));
    LocalMux I__1888 (
            .O(N__17459),
            .I(N__17440));
    Odrv4 I__1887 (
            .O(N__17456),
            .I(\b2v_inst16.N_416 ));
    LocalMux I__1886 (
            .O(N__17445),
            .I(\b2v_inst16.N_416 ));
    Odrv4 I__1885 (
            .O(N__17440),
            .I(\b2v_inst16.N_416 ));
    InMux I__1884 (
            .O(N__17433),
            .I(N__17430));
    LocalMux I__1883 (
            .O(N__17430),
            .I(\b2v_inst16.count_4_9 ));
    InMux I__1882 (
            .O(N__17427),
            .I(N__17424));
    LocalMux I__1881 (
            .O(N__17424),
            .I(\b2v_inst16.count_4_10 ));
    InMux I__1880 (
            .O(N__17421),
            .I(N__17415));
    InMux I__1879 (
            .O(N__17420),
            .I(N__17415));
    LocalMux I__1878 (
            .O(N__17415),
            .I(\b2v_inst16.count_rst ));
    InMux I__1877 (
            .O(N__17412),
            .I(N__17409));
    LocalMux I__1876 (
            .O(N__17409),
            .I(N__17405));
    InMux I__1875 (
            .O(N__17408),
            .I(N__17402));
    Odrv4 I__1874 (
            .O(N__17405),
            .I(\b2v_inst16.countZ0Z_10 ));
    LocalMux I__1873 (
            .O(N__17402),
            .I(\b2v_inst16.countZ0Z_10 ));
    InMux I__1872 (
            .O(N__17397),
            .I(N__17393));
    InMux I__1871 (
            .O(N__17396),
            .I(N__17390));
    LocalMux I__1870 (
            .O(N__17393),
            .I(\b2v_inst16.count_rst_1 ));
    LocalMux I__1869 (
            .O(N__17390),
            .I(\b2v_inst16.count_rst_1 ));
    InMux I__1868 (
            .O(N__17385),
            .I(N__17382));
    LocalMux I__1867 (
            .O(N__17382),
            .I(\b2v_inst16.count_4_12 ));
    CascadeMux I__1866 (
            .O(N__17379),
            .I(\b2v_inst11.curr_state_3_0_cascade_ ));
    CascadeMux I__1865 (
            .O(N__17376),
            .I(\b2v_inst11.curr_stateZ0Z_0_cascade_ ));
    InMux I__1864 (
            .O(N__17373),
            .I(\b2v_inst16.un4_count_1_cry_10 ));
    InMux I__1863 (
            .O(N__17370),
            .I(\b2v_inst16.un4_count_1_cry_11 ));
    InMux I__1862 (
            .O(N__17367),
            .I(\b2v_inst16.un4_count_1_cry_12 ));
    InMux I__1861 (
            .O(N__17364),
            .I(\b2v_inst16.un4_count_1_cry_13 ));
    InMux I__1860 (
            .O(N__17361),
            .I(\b2v_inst16.un4_count_1_cry_14 ));
    InMux I__1859 (
            .O(N__17358),
            .I(N__17354));
    InMux I__1858 (
            .O(N__17357),
            .I(N__17351));
    LocalMux I__1857 (
            .O(N__17354),
            .I(\b2v_inst16.countZ0Z_12 ));
    LocalMux I__1856 (
            .O(N__17351),
            .I(\b2v_inst16.countZ0Z_12 ));
    InMux I__1855 (
            .O(N__17346),
            .I(N__17342));
    InMux I__1854 (
            .O(N__17345),
            .I(N__17339));
    LocalMux I__1853 (
            .O(N__17342),
            .I(N__17334));
    LocalMux I__1852 (
            .O(N__17339),
            .I(N__17334));
    Odrv4 I__1851 (
            .O(N__17334),
            .I(\b2v_inst16.un4_count_1_cry_7_THRU_CO ));
    CascadeMux I__1850 (
            .O(N__17331),
            .I(N__17328));
    InMux I__1849 (
            .O(N__17328),
            .I(N__17323));
    InMux I__1848 (
            .O(N__17327),
            .I(N__17320));
    InMux I__1847 (
            .O(N__17326),
            .I(N__17317));
    LocalMux I__1846 (
            .O(N__17323),
            .I(N__17314));
    LocalMux I__1845 (
            .O(N__17320),
            .I(N__17311));
    LocalMux I__1844 (
            .O(N__17317),
            .I(\b2v_inst16.countZ0Z_8 ));
    Odrv4 I__1843 (
            .O(N__17314),
            .I(\b2v_inst16.countZ0Z_8 ));
    Odrv4 I__1842 (
            .O(N__17311),
            .I(\b2v_inst16.countZ0Z_8 ));
    InMux I__1841 (
            .O(N__17304),
            .I(N__17301));
    LocalMux I__1840 (
            .O(N__17301),
            .I(\b2v_inst16.count_rst_13 ));
    CascadeMux I__1839 (
            .O(N__17298),
            .I(\b2v_inst16.count_rst_14_cascade_ ));
    InMux I__1838 (
            .O(N__17295),
            .I(N__17291));
    CascadeMux I__1837 (
            .O(N__17294),
            .I(N__17288));
    LocalMux I__1836 (
            .O(N__17291),
            .I(N__17284));
    InMux I__1835 (
            .O(N__17288),
            .I(N__17281));
    InMux I__1834 (
            .O(N__17287),
            .I(N__17278));
    Odrv4 I__1833 (
            .O(N__17284),
            .I(\b2v_inst16.countZ0Z_9 ));
    LocalMux I__1832 (
            .O(N__17281),
            .I(\b2v_inst16.countZ0Z_9 ));
    LocalMux I__1831 (
            .O(N__17278),
            .I(\b2v_inst16.countZ0Z_9 ));
    InMux I__1830 (
            .O(N__17271),
            .I(N__17264));
    InMux I__1829 (
            .O(N__17270),
            .I(N__17264));
    CascadeMux I__1828 (
            .O(N__17269),
            .I(N__17261));
    LocalMux I__1827 (
            .O(N__17264),
            .I(N__17258));
    InMux I__1826 (
            .O(N__17261),
            .I(N__17255));
    Odrv4 I__1825 (
            .O(N__17258),
            .I(\b2v_inst16.countZ0Z_3 ));
    LocalMux I__1824 (
            .O(N__17255),
            .I(\b2v_inst16.countZ0Z_3 ));
    InMux I__1823 (
            .O(N__17250),
            .I(N__17246));
    InMux I__1822 (
            .O(N__17249),
            .I(N__17243));
    LocalMux I__1821 (
            .O(N__17246),
            .I(\b2v_inst16.un4_count_1_cry_2_THRU_CO ));
    LocalMux I__1820 (
            .O(N__17243),
            .I(\b2v_inst16.un4_count_1_cry_2_THRU_CO ));
    InMux I__1819 (
            .O(N__17238),
            .I(\b2v_inst16.un4_count_1_cry_2 ));
    InMux I__1818 (
            .O(N__17235),
            .I(N__17230));
    InMux I__1817 (
            .O(N__17234),
            .I(N__17227));
    InMux I__1816 (
            .O(N__17233),
            .I(N__17224));
    LocalMux I__1815 (
            .O(N__17230),
            .I(\b2v_inst16.countZ0Z_4 ));
    LocalMux I__1814 (
            .O(N__17227),
            .I(\b2v_inst16.countZ0Z_4 ));
    LocalMux I__1813 (
            .O(N__17224),
            .I(\b2v_inst16.countZ0Z_4 ));
    CascadeMux I__1812 (
            .O(N__17217),
            .I(N__17213));
    InMux I__1811 (
            .O(N__17216),
            .I(N__17210));
    InMux I__1810 (
            .O(N__17213),
            .I(N__17207));
    LocalMux I__1809 (
            .O(N__17210),
            .I(\b2v_inst16.un4_count_1_cry_3_THRU_CO ));
    LocalMux I__1808 (
            .O(N__17207),
            .I(\b2v_inst16.un4_count_1_cry_3_THRU_CO ));
    InMux I__1807 (
            .O(N__17202),
            .I(\b2v_inst16.un4_count_1_cry_3 ));
    InMux I__1806 (
            .O(N__17199),
            .I(N__17196));
    LocalMux I__1805 (
            .O(N__17196),
            .I(N__17192));
    InMux I__1804 (
            .O(N__17195),
            .I(N__17189));
    Span4Mux_v I__1803 (
            .O(N__17192),
            .I(N__17185));
    LocalMux I__1802 (
            .O(N__17189),
            .I(N__17182));
    InMux I__1801 (
            .O(N__17188),
            .I(N__17179));
    Odrv4 I__1800 (
            .O(N__17185),
            .I(\b2v_inst16.countZ0Z_5 ));
    Odrv4 I__1799 (
            .O(N__17182),
            .I(\b2v_inst16.countZ0Z_5 ));
    LocalMux I__1798 (
            .O(N__17179),
            .I(\b2v_inst16.countZ0Z_5 ));
    CascadeMux I__1797 (
            .O(N__17172),
            .I(N__17168));
    InMux I__1796 (
            .O(N__17171),
            .I(N__17165));
    InMux I__1795 (
            .O(N__17168),
            .I(N__17162));
    LocalMux I__1794 (
            .O(N__17165),
            .I(N__17157));
    LocalMux I__1793 (
            .O(N__17162),
            .I(N__17157));
    Span4Mux_s1_h I__1792 (
            .O(N__17157),
            .I(N__17154));
    Odrv4 I__1791 (
            .O(N__17154),
            .I(\b2v_inst16.un4_count_1_cry_4_THRU_CO ));
    InMux I__1790 (
            .O(N__17151),
            .I(\b2v_inst16.un4_count_1_cry_4 ));
    InMux I__1789 (
            .O(N__17148),
            .I(N__17144));
    InMux I__1788 (
            .O(N__17147),
            .I(N__17141));
    LocalMux I__1787 (
            .O(N__17144),
            .I(\b2v_inst16.countZ0Z_6 ));
    LocalMux I__1786 (
            .O(N__17141),
            .I(\b2v_inst16.countZ0Z_6 ));
    InMux I__1785 (
            .O(N__17136),
            .I(\b2v_inst16.un4_count_1_cry_5 ));
    CascadeMux I__1784 (
            .O(N__17133),
            .I(N__17129));
    InMux I__1783 (
            .O(N__17132),
            .I(N__17126));
    InMux I__1782 (
            .O(N__17129),
            .I(N__17123));
    LocalMux I__1781 (
            .O(N__17126),
            .I(N__17119));
    LocalMux I__1780 (
            .O(N__17123),
            .I(N__17116));
    CascadeMux I__1779 (
            .O(N__17122),
            .I(N__17113));
    Span4Mux_v I__1778 (
            .O(N__17119),
            .I(N__17110));
    Span4Mux_v I__1777 (
            .O(N__17116),
            .I(N__17107));
    InMux I__1776 (
            .O(N__17113),
            .I(N__17104));
    Odrv4 I__1775 (
            .O(N__17110),
            .I(\b2v_inst16.countZ0Z_7 ));
    Odrv4 I__1774 (
            .O(N__17107),
            .I(\b2v_inst16.countZ0Z_7 ));
    LocalMux I__1773 (
            .O(N__17104),
            .I(\b2v_inst16.countZ0Z_7 ));
    InMux I__1772 (
            .O(N__17097),
            .I(N__17091));
    InMux I__1771 (
            .O(N__17096),
            .I(N__17091));
    LocalMux I__1770 (
            .O(N__17091),
            .I(N__17088));
    Span4Mux_s1_h I__1769 (
            .O(N__17088),
            .I(N__17085));
    Odrv4 I__1768 (
            .O(N__17085),
            .I(\b2v_inst16.un4_count_1_cry_6_THRU_CO ));
    InMux I__1767 (
            .O(N__17082),
            .I(\b2v_inst16.un4_count_1_cry_6 ));
    InMux I__1766 (
            .O(N__17079),
            .I(\b2v_inst16.un4_count_1_cry_7 ));
    InMux I__1765 (
            .O(N__17076),
            .I(bfn_2_7_0_));
    InMux I__1764 (
            .O(N__17073),
            .I(\b2v_inst16.un4_count_1_cry_9 ));
    InMux I__1763 (
            .O(N__17070),
            .I(N__17066));
    InMux I__1762 (
            .O(N__17069),
            .I(N__17063));
    LocalMux I__1761 (
            .O(N__17066),
            .I(N__17059));
    LocalMux I__1760 (
            .O(N__17063),
            .I(N__17056));
    InMux I__1759 (
            .O(N__17062),
            .I(N__17053));
    Odrv4 I__1758 (
            .O(N__17059),
            .I(\b2v_inst16.countZ0Z_11 ));
    Odrv4 I__1757 (
            .O(N__17056),
            .I(\b2v_inst16.countZ0Z_11 ));
    LocalMux I__1756 (
            .O(N__17053),
            .I(\b2v_inst16.countZ0Z_11 ));
    InMux I__1755 (
            .O(N__17046),
            .I(N__17040));
    InMux I__1754 (
            .O(N__17045),
            .I(N__17040));
    LocalMux I__1753 (
            .O(N__17040),
            .I(N__17037));
    Odrv4 I__1752 (
            .O(N__17037),
            .I(\b2v_inst16.un4_count_1_cry_10_THRU_CO ));
    InMux I__1751 (
            .O(N__17034),
            .I(N__17031));
    LocalMux I__1750 (
            .O(N__17031),
            .I(N__17027));
    InMux I__1749 (
            .O(N__17030),
            .I(N__17024));
    Odrv4 I__1748 (
            .O(N__17027),
            .I(\b2v_inst36.count_rst_0 ));
    LocalMux I__1747 (
            .O(N__17024),
            .I(\b2v_inst36.count_rst_0 ));
    InMux I__1746 (
            .O(N__17019),
            .I(N__17016));
    LocalMux I__1745 (
            .O(N__17016),
            .I(\b2v_inst36.count_2_14 ));
    CEMux I__1744 (
            .O(N__17013),
            .I(N__17008));
    CEMux I__1743 (
            .O(N__17012),
            .I(N__17005));
    CEMux I__1742 (
            .O(N__17011),
            .I(N__17002));
    LocalMux I__1741 (
            .O(N__17008),
            .I(N__16994));
    LocalMux I__1740 (
            .O(N__17005),
            .I(N__16994));
    LocalMux I__1739 (
            .O(N__17002),
            .I(N__16994));
    CEMux I__1738 (
            .O(N__17001),
            .I(N__16979));
    Span4Mux_s2_v I__1737 (
            .O(N__16994),
            .I(N__16976));
    InMux I__1736 (
            .O(N__16993),
            .I(N__16973));
    InMux I__1735 (
            .O(N__16992),
            .I(N__16968));
    InMux I__1734 (
            .O(N__16991),
            .I(N__16968));
    InMux I__1733 (
            .O(N__16990),
            .I(N__16959));
    InMux I__1732 (
            .O(N__16989),
            .I(N__16959));
    InMux I__1731 (
            .O(N__16988),
            .I(N__16959));
    InMux I__1730 (
            .O(N__16987),
            .I(N__16959));
    InMux I__1729 (
            .O(N__16986),
            .I(N__16948));
    InMux I__1728 (
            .O(N__16985),
            .I(N__16948));
    InMux I__1727 (
            .O(N__16984),
            .I(N__16948));
    InMux I__1726 (
            .O(N__16983),
            .I(N__16948));
    InMux I__1725 (
            .O(N__16982),
            .I(N__16948));
    LocalMux I__1724 (
            .O(N__16979),
            .I(N__16939));
    Span4Mux_s1_h I__1723 (
            .O(N__16976),
            .I(N__16924));
    LocalMux I__1722 (
            .O(N__16973),
            .I(N__16924));
    LocalMux I__1721 (
            .O(N__16968),
            .I(N__16924));
    LocalMux I__1720 (
            .O(N__16959),
            .I(N__16924));
    LocalMux I__1719 (
            .O(N__16948),
            .I(N__16924));
    InMux I__1718 (
            .O(N__16947),
            .I(N__16917));
    InMux I__1717 (
            .O(N__16946),
            .I(N__16917));
    InMux I__1716 (
            .O(N__16945),
            .I(N__16917));
    CEMux I__1715 (
            .O(N__16944),
            .I(N__16911));
    CEMux I__1714 (
            .O(N__16943),
            .I(N__16908));
    CEMux I__1713 (
            .O(N__16942),
            .I(N__16905));
    Span4Mux_s2_h I__1712 (
            .O(N__16939),
            .I(N__16902));
    InMux I__1711 (
            .O(N__16938),
            .I(N__16893));
    InMux I__1710 (
            .O(N__16937),
            .I(N__16893));
    InMux I__1709 (
            .O(N__16936),
            .I(N__16893));
    InMux I__1708 (
            .O(N__16935),
            .I(N__16893));
    Sp12to4 I__1707 (
            .O(N__16924),
            .I(N__16888));
    LocalMux I__1706 (
            .O(N__16917),
            .I(N__16888));
    InMux I__1705 (
            .O(N__16916),
            .I(N__16881));
    InMux I__1704 (
            .O(N__16915),
            .I(N__16881));
    InMux I__1703 (
            .O(N__16914),
            .I(N__16881));
    LocalMux I__1702 (
            .O(N__16911),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    LocalMux I__1701 (
            .O(N__16908),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    LocalMux I__1700 (
            .O(N__16905),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    Odrv4 I__1699 (
            .O(N__16902),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    LocalMux I__1698 (
            .O(N__16893),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    Odrv12 I__1697 (
            .O(N__16888),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    LocalMux I__1696 (
            .O(N__16881),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ));
    InMux I__1695 (
            .O(N__16866),
            .I(N__16860));
    InMux I__1694 (
            .O(N__16865),
            .I(N__16860));
    LocalMux I__1693 (
            .O(N__16860),
            .I(N__16857));
    Odrv4 I__1692 (
            .O(N__16857),
            .I(\b2v_inst36.count_rst ));
    CascadeMux I__1691 (
            .O(N__16854),
            .I(\b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_ ));
    InMux I__1690 (
            .O(N__16851),
            .I(N__16848));
    LocalMux I__1689 (
            .O(N__16848),
            .I(\b2v_inst36.count_2_15 ));
    InMux I__1688 (
            .O(N__16845),
            .I(N__16841));
    InMux I__1687 (
            .O(N__16844),
            .I(N__16838));
    LocalMux I__1686 (
            .O(N__16841),
            .I(N__16833));
    LocalMux I__1685 (
            .O(N__16838),
            .I(N__16833));
    Odrv4 I__1684 (
            .O(N__16833),
            .I(\b2v_inst36.countZ0Z_15 ));
    CascadeMux I__1683 (
            .O(N__16830),
            .I(\b2v_inst16.count_en_cascade_ ));
    InMux I__1682 (
            .O(N__16827),
            .I(N__16823));
    InMux I__1681 (
            .O(N__16826),
            .I(N__16820));
    LocalMux I__1680 (
            .O(N__16823),
            .I(\b2v_inst16.un4_count_1_axb_1 ));
    LocalMux I__1679 (
            .O(N__16820),
            .I(\b2v_inst16.un4_count_1_axb_1 ));
    CascadeMux I__1678 (
            .O(N__16815),
            .I(N__16812));
    InMux I__1677 (
            .O(N__16812),
            .I(N__16806));
    InMux I__1676 (
            .O(N__16811),
            .I(N__16801));
    InMux I__1675 (
            .O(N__16810),
            .I(N__16801));
    InMux I__1674 (
            .O(N__16809),
            .I(N__16798));
    LocalMux I__1673 (
            .O(N__16806),
            .I(\b2v_inst16.countZ0Z_0 ));
    LocalMux I__1672 (
            .O(N__16801),
            .I(\b2v_inst16.countZ0Z_0 ));
    LocalMux I__1671 (
            .O(N__16798),
            .I(\b2v_inst16.countZ0Z_0 ));
    InMux I__1670 (
            .O(N__16791),
            .I(N__16787));
    InMux I__1669 (
            .O(N__16790),
            .I(N__16784));
    LocalMux I__1668 (
            .O(N__16787),
            .I(\b2v_inst16.countZ0Z_2 ));
    LocalMux I__1667 (
            .O(N__16784),
            .I(\b2v_inst16.countZ0Z_2 ));
    InMux I__1666 (
            .O(N__16779),
            .I(\b2v_inst16.un4_count_1_cry_1 ));
    InMux I__1665 (
            .O(N__16776),
            .I(N__16773));
    LocalMux I__1664 (
            .O(N__16773),
            .I(\b2v_inst36.count_2_12 ));
    InMux I__1663 (
            .O(N__16770),
            .I(N__16764));
    InMux I__1662 (
            .O(N__16769),
            .I(N__16764));
    LocalMux I__1661 (
            .O(N__16764),
            .I(\b2v_inst36.count_rst_2 ));
    InMux I__1660 (
            .O(N__16761),
            .I(N__16758));
    LocalMux I__1659 (
            .O(N__16758),
            .I(\b2v_inst36.countZ0Z_12 ));
    InMux I__1658 (
            .O(N__16755),
            .I(N__16748));
    InMux I__1657 (
            .O(N__16754),
            .I(N__16748));
    InMux I__1656 (
            .O(N__16753),
            .I(N__16745));
    LocalMux I__1655 (
            .O(N__16748),
            .I(\b2v_inst36.count_rst_5 ));
    LocalMux I__1654 (
            .O(N__16745),
            .I(\b2v_inst36.count_rst_5 ));
    CascadeMux I__1653 (
            .O(N__16740),
            .I(\b2v_inst36.countZ0Z_12_cascade_ ));
    InMux I__1652 (
            .O(N__16737),
            .I(N__16734));
    LocalMux I__1651 (
            .O(N__16734),
            .I(N__16730));
    InMux I__1650 (
            .O(N__16733),
            .I(N__16727));
    Odrv4 I__1649 (
            .O(N__16730),
            .I(\b2v_inst36.count_2_9 ));
    LocalMux I__1648 (
            .O(N__16727),
            .I(\b2v_inst36.count_2_9 ));
    InMux I__1647 (
            .O(N__16722),
            .I(N__16719));
    LocalMux I__1646 (
            .O(N__16719),
            .I(\b2v_inst36.un12_clk_100khz_6 ));
    InMux I__1645 (
            .O(N__16716),
            .I(N__16713));
    LocalMux I__1644 (
            .O(N__16713),
            .I(\b2v_inst36.countZ0Z_14 ));
    CascadeMux I__1643 (
            .O(N__16710),
            .I(\b2v_inst36.countZ0Z_14_cascade_ ));
    InMux I__1642 (
            .O(N__16707),
            .I(N__16702));
    InMux I__1641 (
            .O(N__16706),
            .I(N__16697));
    InMux I__1640 (
            .O(N__16705),
            .I(N__16694));
    LocalMux I__1639 (
            .O(N__16702),
            .I(N__16691));
    InMux I__1638 (
            .O(N__16701),
            .I(N__16686));
    InMux I__1637 (
            .O(N__16700),
            .I(N__16686));
    LocalMux I__1636 (
            .O(N__16697),
            .I(\b2v_inst36.countZ0Z_0 ));
    LocalMux I__1635 (
            .O(N__16694),
            .I(\b2v_inst36.countZ0Z_0 ));
    Odrv4 I__1634 (
            .O(N__16691),
            .I(\b2v_inst36.countZ0Z_0 ));
    LocalMux I__1633 (
            .O(N__16686),
            .I(\b2v_inst36.countZ0Z_0 ));
    InMux I__1632 (
            .O(N__16677),
            .I(N__16674));
    LocalMux I__1631 (
            .O(N__16674),
            .I(\b2v_inst36.un12_clk_100khz_10 ));
    InMux I__1630 (
            .O(N__16671),
            .I(N__16668));
    LocalMux I__1629 (
            .O(N__16668),
            .I(\b2v_inst36.count_2_13 ));
    InMux I__1628 (
            .O(N__16665),
            .I(N__16659));
    InMux I__1627 (
            .O(N__16664),
            .I(N__16659));
    LocalMux I__1626 (
            .O(N__16659),
            .I(\b2v_inst36.count_rst_1 ));
    InMux I__1625 (
            .O(N__16656),
            .I(N__16652));
    InMux I__1624 (
            .O(N__16655),
            .I(N__16649));
    LocalMux I__1623 (
            .O(N__16652),
            .I(\b2v_inst36.countZ0Z_13 ));
    LocalMux I__1622 (
            .O(N__16649),
            .I(\b2v_inst36.countZ0Z_13 ));
    InMux I__1621 (
            .O(N__16644),
            .I(N__16641));
    LocalMux I__1620 (
            .O(N__16641),
            .I(N__16637));
    InMux I__1619 (
            .O(N__16640),
            .I(N__16634));
    Odrv4 I__1618 (
            .O(N__16637),
            .I(\b2v_inst36.un2_count_1_axb_8 ));
    LocalMux I__1617 (
            .O(N__16634),
            .I(\b2v_inst36.un2_count_1_axb_8 ));
    CascadeMux I__1616 (
            .O(N__16629),
            .I(N__16625));
    InMux I__1615 (
            .O(N__16628),
            .I(N__16620));
    InMux I__1614 (
            .O(N__16625),
            .I(N__16620));
    LocalMux I__1613 (
            .O(N__16620),
            .I(\b2v_inst36.un2_count_1_cry_7_THRU_CO ));
    InMux I__1612 (
            .O(N__16617),
            .I(\b2v_inst36.un2_count_1_cry_7 ));
    InMux I__1611 (
            .O(N__16614),
            .I(bfn_2_3_0_));
    CascadeMux I__1610 (
            .O(N__16611),
            .I(N__16607));
    InMux I__1609 (
            .O(N__16610),
            .I(N__16603));
    InMux I__1608 (
            .O(N__16607),
            .I(N__16600));
    InMux I__1607 (
            .O(N__16606),
            .I(N__16597));
    LocalMux I__1606 (
            .O(N__16603),
            .I(N__16592));
    LocalMux I__1605 (
            .O(N__16600),
            .I(N__16592));
    LocalMux I__1604 (
            .O(N__16597),
            .I(N__16589));
    Odrv12 I__1603 (
            .O(N__16592),
            .I(\b2v_inst36.countZ0Z_10 ));
    Odrv4 I__1602 (
            .O(N__16589),
            .I(\b2v_inst36.countZ0Z_10 ));
    InMux I__1601 (
            .O(N__16584),
            .I(N__16580));
    CascadeMux I__1600 (
            .O(N__16583),
            .I(N__16577));
    LocalMux I__1599 (
            .O(N__16580),
            .I(N__16574));
    InMux I__1598 (
            .O(N__16577),
            .I(N__16571));
    Span4Mux_s2_v I__1597 (
            .O(N__16574),
            .I(N__16566));
    LocalMux I__1596 (
            .O(N__16571),
            .I(N__16566));
    Odrv4 I__1595 (
            .O(N__16566),
            .I(\b2v_inst36.un2_count_1_cry_9_THRU_CO ));
    InMux I__1594 (
            .O(N__16563),
            .I(\b2v_inst36.un2_count_1_cry_9 ));
    InMux I__1593 (
            .O(N__16560),
            .I(N__16556));
    InMux I__1592 (
            .O(N__16559),
            .I(N__16552));
    LocalMux I__1591 (
            .O(N__16556),
            .I(N__16549));
    InMux I__1590 (
            .O(N__16555),
            .I(N__16546));
    LocalMux I__1589 (
            .O(N__16552),
            .I(\b2v_inst36.countZ0Z_11 ));
    Odrv4 I__1588 (
            .O(N__16549),
            .I(\b2v_inst36.countZ0Z_11 ));
    LocalMux I__1587 (
            .O(N__16546),
            .I(\b2v_inst36.countZ0Z_11 ));
    InMux I__1586 (
            .O(N__16539),
            .I(N__16535));
    InMux I__1585 (
            .O(N__16538),
            .I(N__16532));
    LocalMux I__1584 (
            .O(N__16535),
            .I(\b2v_inst36.un2_count_1_cry_10_THRU_CO ));
    LocalMux I__1583 (
            .O(N__16532),
            .I(\b2v_inst36.un2_count_1_cry_10_THRU_CO ));
    InMux I__1582 (
            .O(N__16527),
            .I(\b2v_inst36.un2_count_1_cry_10 ));
    InMux I__1581 (
            .O(N__16524),
            .I(\b2v_inst36.un2_count_1_cry_11 ));
    InMux I__1580 (
            .O(N__16521),
            .I(\b2v_inst36.un2_count_1_cry_12 ));
    InMux I__1579 (
            .O(N__16518),
            .I(\b2v_inst36.un2_count_1_cry_13 ));
    InMux I__1578 (
            .O(N__16515),
            .I(\b2v_inst36.un2_count_1_cry_14 ));
    InMux I__1577 (
            .O(N__16512),
            .I(N__16509));
    LocalMux I__1576 (
            .O(N__16509),
            .I(\b2v_inst36.un2_count_1_axb_9 ));
    InMux I__1575 (
            .O(N__16506),
            .I(N__16503));
    LocalMux I__1574 (
            .O(N__16503),
            .I(\b2v_inst36.count_2_7 ));
    CascadeMux I__1573 (
            .O(N__16500),
            .I(N__16497));
    InMux I__1572 (
            .O(N__16497),
            .I(N__16492));
    InMux I__1571 (
            .O(N__16496),
            .I(N__16487));
    InMux I__1570 (
            .O(N__16495),
            .I(N__16487));
    LocalMux I__1569 (
            .O(N__16492),
            .I(N__16484));
    LocalMux I__1568 (
            .O(N__16487),
            .I(\b2v_inst36.un2_count_1_axb_1 ));
    Odrv4 I__1567 (
            .O(N__16484),
            .I(\b2v_inst36.un2_count_1_axb_1 ));
    CascadeMux I__1566 (
            .O(N__16479),
            .I(N__16475));
    InMux I__1565 (
            .O(N__16478),
            .I(N__16469));
    InMux I__1564 (
            .O(N__16475),
            .I(N__16469));
    InMux I__1563 (
            .O(N__16474),
            .I(N__16466));
    LocalMux I__1562 (
            .O(N__16469),
            .I(\b2v_inst36.un2_count_1_axb_2 ));
    LocalMux I__1561 (
            .O(N__16466),
            .I(\b2v_inst36.un2_count_1_axb_2 ));
    CascadeMux I__1560 (
            .O(N__16461),
            .I(N__16458));
    InMux I__1559 (
            .O(N__16458),
            .I(N__16452));
    InMux I__1558 (
            .O(N__16457),
            .I(N__16452));
    LocalMux I__1557 (
            .O(N__16452),
            .I(\b2v_inst36.un2_count_1_cry_1_THRU_CO ));
    InMux I__1556 (
            .O(N__16449),
            .I(\b2v_inst36.un2_count_1_cry_1 ));
    InMux I__1555 (
            .O(N__16446),
            .I(N__16439));
    InMux I__1554 (
            .O(N__16445),
            .I(N__16439));
    InMux I__1553 (
            .O(N__16444),
            .I(N__16436));
    LocalMux I__1552 (
            .O(N__16439),
            .I(\b2v_inst36.countZ0Z_3 ));
    LocalMux I__1551 (
            .O(N__16436),
            .I(\b2v_inst36.countZ0Z_3 ));
    CascadeMux I__1550 (
            .O(N__16431),
            .I(N__16427));
    CascadeMux I__1549 (
            .O(N__16430),
            .I(N__16424));
    InMux I__1548 (
            .O(N__16427),
            .I(N__16419));
    InMux I__1547 (
            .O(N__16424),
            .I(N__16419));
    LocalMux I__1546 (
            .O(N__16419),
            .I(\b2v_inst36.un2_count_1_cry_2_THRU_CO ));
    InMux I__1545 (
            .O(N__16416),
            .I(\b2v_inst36.un2_count_1_cry_2 ));
    CascadeMux I__1544 (
            .O(N__16413),
            .I(N__16410));
    InMux I__1543 (
            .O(N__16410),
            .I(N__16407));
    LocalMux I__1542 (
            .O(N__16407),
            .I(\b2v_inst36.un2_count_1_axb_4 ));
    InMux I__1541 (
            .O(N__16404),
            .I(N__16397));
    InMux I__1540 (
            .O(N__16403),
            .I(N__16397));
    InMux I__1539 (
            .O(N__16402),
            .I(N__16394));
    LocalMux I__1538 (
            .O(N__16397),
            .I(\b2v_inst36.count_rst_10 ));
    LocalMux I__1537 (
            .O(N__16394),
            .I(\b2v_inst36.count_rst_10 ));
    InMux I__1536 (
            .O(N__16389),
            .I(\b2v_inst36.un2_count_1_cry_3 ));
    InMux I__1535 (
            .O(N__16386),
            .I(N__16382));
    InMux I__1534 (
            .O(N__16385),
            .I(N__16379));
    LocalMux I__1533 (
            .O(N__16382),
            .I(\b2v_inst36.un2_count_1_axb_5 ));
    LocalMux I__1532 (
            .O(N__16379),
            .I(\b2v_inst36.un2_count_1_axb_5 ));
    InMux I__1531 (
            .O(N__16374),
            .I(N__16368));
    InMux I__1530 (
            .O(N__16373),
            .I(N__16368));
    LocalMux I__1529 (
            .O(N__16368),
            .I(\b2v_inst36.un2_count_1_cry_4_THRU_CO ));
    InMux I__1528 (
            .O(N__16365),
            .I(\b2v_inst36.un2_count_1_cry_4 ));
    InMux I__1527 (
            .O(N__16362),
            .I(N__16359));
    LocalMux I__1526 (
            .O(N__16359),
            .I(\b2v_inst36.un2_count_1_axb_6 ));
    InMux I__1525 (
            .O(N__16356),
            .I(N__16347));
    InMux I__1524 (
            .O(N__16355),
            .I(N__16347));
    InMux I__1523 (
            .O(N__16354),
            .I(N__16347));
    LocalMux I__1522 (
            .O(N__16347),
            .I(\b2v_inst36.un2_count_1_cry_5_c_RNIE2FZ0Z8 ));
    InMux I__1521 (
            .O(N__16344),
            .I(\b2v_inst36.un2_count_1_cry_5 ));
    CascadeMux I__1520 (
            .O(N__16341),
            .I(N__16338));
    InMux I__1519 (
            .O(N__16338),
            .I(N__16333));
    InMux I__1518 (
            .O(N__16337),
            .I(N__16329));
    InMux I__1517 (
            .O(N__16336),
            .I(N__16326));
    LocalMux I__1516 (
            .O(N__16333),
            .I(N__16323));
    InMux I__1515 (
            .O(N__16332),
            .I(N__16320));
    LocalMux I__1514 (
            .O(N__16329),
            .I(\b2v_inst36.countZ0Z_7 ));
    LocalMux I__1513 (
            .O(N__16326),
            .I(\b2v_inst36.countZ0Z_7 ));
    Odrv4 I__1512 (
            .O(N__16323),
            .I(\b2v_inst36.countZ0Z_7 ));
    LocalMux I__1511 (
            .O(N__16320),
            .I(\b2v_inst36.countZ0Z_7 ));
    InMux I__1510 (
            .O(N__16311),
            .I(N__16307));
    InMux I__1509 (
            .O(N__16310),
            .I(N__16304));
    LocalMux I__1508 (
            .O(N__16307),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    LocalMux I__1507 (
            .O(N__16304),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    InMux I__1506 (
            .O(N__16299),
            .I(\b2v_inst36.un2_count_1_cry_6 ));
    InMux I__1505 (
            .O(N__16296),
            .I(bfn_1_16_0_));
    CascadeMux I__1504 (
            .O(N__16293),
            .I(\b2v_inst36.count_rst_12_cascade_ ));
    InMux I__1503 (
            .O(N__16290),
            .I(N__16287));
    LocalMux I__1502 (
            .O(N__16287),
            .I(\b2v_inst36.count_rst_12 ));
    CascadeMux I__1501 (
            .O(N__16284),
            .I(\b2v_inst36.countZ0Z_3_cascade_ ));
    InMux I__1500 (
            .O(N__16281),
            .I(N__16278));
    LocalMux I__1499 (
            .O(N__16278),
            .I(N__16275));
    Span4Mux_s1_h I__1498 (
            .O(N__16275),
            .I(N__16272));
    Odrv4 I__1497 (
            .O(N__16272),
            .I(\b2v_inst36.un12_clk_100khz_3 ));
    InMux I__1496 (
            .O(N__16269),
            .I(N__16266));
    LocalMux I__1495 (
            .O(N__16266),
            .I(\b2v_inst36.count_rst_11 ));
    InMux I__1494 (
            .O(N__16263),
            .I(N__16257));
    InMux I__1493 (
            .O(N__16262),
            .I(N__16257));
    LocalMux I__1492 (
            .O(N__16257),
            .I(\b2v_inst36.count_2_2 ));
    InMux I__1491 (
            .O(N__16254),
            .I(N__16251));
    LocalMux I__1490 (
            .O(N__16251),
            .I(\b2v_inst36.count_2_3 ));
    InMux I__1489 (
            .O(N__16248),
            .I(N__16242));
    InMux I__1488 (
            .O(N__16247),
            .I(N__16242));
    LocalMux I__1487 (
            .O(N__16242),
            .I(N__16239));
    Odrv4 I__1486 (
            .O(N__16239),
            .I(\b2v_inst11.count_1_6 ));
    InMux I__1485 (
            .O(N__16236),
            .I(N__16233));
    LocalMux I__1484 (
            .O(N__16233),
            .I(\b2v_inst11.count_0_6 ));
    CascadeMux I__1483 (
            .O(N__16230),
            .I(N__16227));
    InMux I__1482 (
            .O(N__16227),
            .I(N__16221));
    InMux I__1481 (
            .O(N__16226),
            .I(N__16221));
    LocalMux I__1480 (
            .O(N__16221),
            .I(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ));
    InMux I__1479 (
            .O(N__16218),
            .I(N__16215));
    LocalMux I__1478 (
            .O(N__16215),
            .I(\b2v_inst11.count_0_15 ));
    InMux I__1477 (
            .O(N__16212),
            .I(\b2v_inst11.un1_count_cry_11 ));
    InMux I__1476 (
            .O(N__16209),
            .I(\b2v_inst11.un1_count_cry_12 ));
    InMux I__1475 (
            .O(N__16206),
            .I(\b2v_inst11.un1_count_cry_13 ));
    InMux I__1474 (
            .O(N__16203),
            .I(\b2v_inst11.un1_count_cry_14 ));
    InMux I__1473 (
            .O(N__16200),
            .I(N__16194));
    InMux I__1472 (
            .O(N__16199),
            .I(N__16194));
    LocalMux I__1471 (
            .O(N__16194),
            .I(N__16191));
    Odrv4 I__1470 (
            .O(N__16191),
            .I(\b2v_inst11.count_1_5 ));
    InMux I__1469 (
            .O(N__16188),
            .I(N__16185));
    LocalMux I__1468 (
            .O(N__16185),
            .I(\b2v_inst11.count_0_5 ));
    InMux I__1467 (
            .O(N__16182),
            .I(N__16178));
    InMux I__1466 (
            .O(N__16181),
            .I(N__16175));
    LocalMux I__1465 (
            .O(N__16178),
            .I(\b2v_inst11.count_1_14 ));
    LocalMux I__1464 (
            .O(N__16175),
            .I(\b2v_inst11.count_1_14 ));
    InMux I__1463 (
            .O(N__16170),
            .I(N__16167));
    LocalMux I__1462 (
            .O(N__16167),
            .I(\b2v_inst11.count_0_14 ));
    InMux I__1461 (
            .O(N__16164),
            .I(\b2v_inst11.un1_count_cry_2_cZ0 ));
    InMux I__1460 (
            .O(N__16161),
            .I(\b2v_inst11.un1_count_cry_3 ));
    InMux I__1459 (
            .O(N__16158),
            .I(\b2v_inst11.un1_count_cry_4 ));
    InMux I__1458 (
            .O(N__16155),
            .I(\b2v_inst11.un1_count_cry_5 ));
    InMux I__1457 (
            .O(N__16152),
            .I(N__16148));
    InMux I__1456 (
            .O(N__16151),
            .I(N__16145));
    LocalMux I__1455 (
            .O(N__16148),
            .I(N__16142));
    LocalMux I__1454 (
            .O(N__16145),
            .I(\b2v_inst11.count_1_7 ));
    Odrv4 I__1453 (
            .O(N__16142),
            .I(\b2v_inst11.count_1_7 ));
    InMux I__1452 (
            .O(N__16137),
            .I(\b2v_inst11.un1_count_cry_6 ));
    InMux I__1451 (
            .O(N__16134),
            .I(\b2v_inst11.un1_count_cry_7 ));
    InMux I__1450 (
            .O(N__16131),
            .I(bfn_1_12_0_));
    InMux I__1449 (
            .O(N__16128),
            .I(\b2v_inst11.un1_count_cry_9 ));
    InMux I__1448 (
            .O(N__16125),
            .I(\b2v_inst11.un1_count_cry_10 ));
    CascadeMux I__1447 (
            .O(N__16122),
            .I(\b2v_inst16.curr_state_7_0_1_cascade_ ));
    InMux I__1446 (
            .O(N__16119),
            .I(N__16116));
    LocalMux I__1445 (
            .O(N__16116),
            .I(N__16113));
    Span4Mux_v I__1444 (
            .O(N__16113),
            .I(N__16110));
    Span4Mux_v I__1443 (
            .O(N__16110),
            .I(N__16107));
    Sp12to4 I__1442 (
            .O(N__16107),
            .I(N__16104));
    Odrv12 I__1441 (
            .O(N__16104),
            .I(vddq_ok));
    CascadeMux I__1440 (
            .O(N__16101),
            .I(\b2v_inst16.N_208_0_cascade_ ));
    CascadeMux I__1439 (
            .O(N__16098),
            .I(\b2v_inst16.curr_state_RNIBO6I1Z0Z_0_cascade_ ));
    InMux I__1438 (
            .O(N__16095),
            .I(N__16092));
    LocalMux I__1437 (
            .O(N__16092),
            .I(\b2v_inst16.curr_state_2_1 ));
    InMux I__1436 (
            .O(N__16089),
            .I(N__16086));
    LocalMux I__1435 (
            .O(N__16086),
            .I(\b2v_inst16.curr_state_2_0 ));
    CascadeMux I__1434 (
            .O(N__16083),
            .I(N__16080));
    InMux I__1433 (
            .O(N__16080),
            .I(N__16077));
    LocalMux I__1432 (
            .O(N__16077),
            .I(\b2v_inst11.count_0_7 ));
    InMux I__1431 (
            .O(N__16074),
            .I(\b2v_inst11.un1_count_cry_1_cZ0 ));
    CascadeMux I__1430 (
            .O(N__16071),
            .I(\b2v_inst16.countZ0Z_7_cascade_ ));
    InMux I__1429 (
            .O(N__16068),
            .I(N__16065));
    LocalMux I__1428 (
            .O(N__16065),
            .I(\b2v_inst16.count_4_7 ));
    CascadeMux I__1427 (
            .O(N__16062),
            .I(\b2v_inst16.count_rst_10_cascade_ ));
    CascadeMux I__1426 (
            .O(N__16059),
            .I(\b2v_inst16.countZ0Z_5_cascade_ ));
    InMux I__1425 (
            .O(N__16056),
            .I(N__16053));
    LocalMux I__1424 (
            .O(N__16053),
            .I(\b2v_inst16.count_4_5 ));
    CascadeMux I__1423 (
            .O(N__16050),
            .I(\b2v_inst16.countZ0Z_8_cascade_ ));
    InMux I__1422 (
            .O(N__16047),
            .I(N__16044));
    LocalMux I__1421 (
            .O(N__16044),
            .I(\b2v_inst16.count_4_8 ));
    InMux I__1420 (
            .O(N__16041),
            .I(N__16038));
    LocalMux I__1419 (
            .O(N__16038),
            .I(\b2v_inst16.count_rst_12 ));
    CascadeMux I__1418 (
            .O(N__16035),
            .I(\b2v_inst16.N_416_cascade_ ));
    InMux I__1417 (
            .O(N__16032),
            .I(N__16029));
    LocalMux I__1416 (
            .O(N__16029),
            .I(\b2v_inst16.count_rst_8 ));
    CascadeMux I__1415 (
            .O(N__16026),
            .I(\b2v_inst16.count_RNIE4RF_2Z0Z_1_cascade_ ));
    CascadeMux I__1414 (
            .O(N__16023),
            .I(\b2v_inst16.count_rst_5_cascade_ ));
    InMux I__1413 (
            .O(N__16020),
            .I(N__16014));
    InMux I__1412 (
            .O(N__16019),
            .I(N__16014));
    LocalMux I__1411 (
            .O(N__16014),
            .I(\b2v_inst16.N_414 ));
    CascadeMux I__1410 (
            .O(N__16011),
            .I(\b2v_inst16.countZ0Z_0_cascade_ ));
    InMux I__1409 (
            .O(N__16008),
            .I(N__16005));
    LocalMux I__1408 (
            .O(N__16005),
            .I(\b2v_inst16.count_4_0 ));
    InMux I__1407 (
            .O(N__16002),
            .I(N__15999));
    LocalMux I__1406 (
            .O(N__15999),
            .I(\b2v_inst16.countZ0Z_1 ));
    InMux I__1405 (
            .O(N__15996),
            .I(N__15993));
    LocalMux I__1404 (
            .O(N__15993),
            .I(\b2v_inst16.count_4_i_a3_7_0 ));
    InMux I__1403 (
            .O(N__15990),
            .I(N__15984));
    InMux I__1402 (
            .O(N__15989),
            .I(N__15984));
    LocalMux I__1401 (
            .O(N__15984),
            .I(\b2v_inst16.count_RNIE4RF_2Z0Z_1 ));
    CascadeMux I__1400 (
            .O(N__15981),
            .I(N__15977));
    InMux I__1399 (
            .O(N__15980),
            .I(N__15972));
    InMux I__1398 (
            .O(N__15977),
            .I(N__15972));
    LocalMux I__1397 (
            .O(N__15972),
            .I(\b2v_inst16.count_4_1 ));
    CascadeMux I__1396 (
            .O(N__15969),
            .I(\b2v_inst16.count_rst_9_cascade_ ));
    CascadeMux I__1395 (
            .O(N__15966),
            .I(\b2v_inst16.countZ0Z_4_cascade_ ));
    InMux I__1394 (
            .O(N__15963),
            .I(N__15960));
    LocalMux I__1393 (
            .O(N__15960),
            .I(\b2v_inst16.count_4_4 ));
    CascadeMux I__1392 (
            .O(N__15957),
            .I(\b2v_inst16.countZ0Z_3_cascade_ ));
    InMux I__1391 (
            .O(N__15954),
            .I(N__15951));
    LocalMux I__1390 (
            .O(N__15951),
            .I(\b2v_inst16.count_4_3 ));
    InMux I__1389 (
            .O(N__15948),
            .I(N__15945));
    LocalMux I__1388 (
            .O(N__15945),
            .I(\b2v_inst16.count_4_i_a3_9_0 ));
    CascadeMux I__1387 (
            .O(N__15942),
            .I(\b2v_inst16.count_4_i_a3_8_0_cascade_ ));
    InMux I__1386 (
            .O(N__15939),
            .I(N__15936));
    LocalMux I__1385 (
            .O(N__15936),
            .I(\b2v_inst16.count_4_i_a3_10_0 ));
    CascadeMux I__1384 (
            .O(N__15933),
            .I(\b2v_inst16.N_414_cascade_ ));
    InMux I__1383 (
            .O(N__15930),
            .I(N__15927));
    LocalMux I__1382 (
            .O(N__15927),
            .I(\b2v_inst36.un12_clk_100khz_1 ));
    CascadeMux I__1381 (
            .O(N__15924),
            .I(\b2v_inst36.un12_clk_100khz_0_cascade_ ));
    InMux I__1380 (
            .O(N__15921),
            .I(N__15918));
    LocalMux I__1379 (
            .O(N__15918),
            .I(N__15915));
    Odrv12 I__1378 (
            .O(N__15915),
            .I(\b2v_inst36.un12_clk_100khz_2 ));
    InMux I__1377 (
            .O(N__15912),
            .I(N__15909));
    LocalMux I__1376 (
            .O(N__15909),
            .I(N__15906));
    Odrv12 I__1375 (
            .O(N__15906),
            .I(\b2v_inst36.un12_clk_100khz_7 ));
    CascadeMux I__1374 (
            .O(N__15903),
            .I(\b2v_inst36.un12_clk_100khz_12_cascade_ ));
    CascadeMux I__1373 (
            .O(N__15900),
            .I(\b2v_inst36.N_1_i_cascade_ ));
    InMux I__1372 (
            .O(N__15897),
            .I(N__15894));
    LocalMux I__1371 (
            .O(N__15894),
            .I(\b2v_inst36.count_2_0 ));
    InMux I__1370 (
            .O(N__15891),
            .I(N__15888));
    LocalMux I__1369 (
            .O(N__15888),
            .I(\b2v_inst36.count_rst_14 ));
    CascadeMux I__1368 (
            .O(N__15885),
            .I(\b2v_inst36.countZ0Z_0_cascade_ ));
    InMux I__1367 (
            .O(N__15882),
            .I(N__15876));
    InMux I__1366 (
            .O(N__15881),
            .I(N__15876));
    LocalMux I__1365 (
            .O(N__15876),
            .I(\b2v_inst36.count_2_1 ));
    CascadeMux I__1364 (
            .O(N__15873),
            .I(\b2v_inst16.count_rst_0_cascade_ ));
    CascadeMux I__1363 (
            .O(N__15870),
            .I(\b2v_inst16.countZ0Z_11_cascade_ ));
    InMux I__1362 (
            .O(N__15867),
            .I(N__15864));
    LocalMux I__1361 (
            .O(N__15864),
            .I(N__15861));
    Odrv4 I__1360 (
            .O(N__15861),
            .I(\b2v_inst16.count_4_11 ));
    InMux I__1359 (
            .O(N__15858),
            .I(N__15855));
    LocalMux I__1358 (
            .O(N__15855),
            .I(\b2v_inst36.count_rst_6 ));
    CascadeMux I__1357 (
            .O(N__15852),
            .I(\b2v_inst36.count_rst_6_cascade_ ));
    CascadeMux I__1356 (
            .O(N__15849),
            .I(\b2v_inst36.un2_count_1_axb_8_cascade_ ));
    InMux I__1355 (
            .O(N__15846),
            .I(N__15840));
    InMux I__1354 (
            .O(N__15845),
            .I(N__15840));
    LocalMux I__1353 (
            .O(N__15840),
            .I(\b2v_inst36.count_2_8 ));
    InMux I__1352 (
            .O(N__15837),
            .I(N__15834));
    LocalMux I__1351 (
            .O(N__15834),
            .I(N__15831));
    Odrv4 I__1350 (
            .O(N__15831),
            .I(\b2v_inst36.count_rst_4 ));
    InMux I__1349 (
            .O(N__15828),
            .I(N__15825));
    LocalMux I__1348 (
            .O(N__15825),
            .I(\b2v_inst36.count_rst_3 ));
    InMux I__1347 (
            .O(N__15822),
            .I(N__15819));
    LocalMux I__1346 (
            .O(N__15819),
            .I(\b2v_inst36.count_rst_13 ));
    CascadeMux I__1345 (
            .O(N__15816),
            .I(\b2v_inst36.count_rst_13_cascade_ ));
    CascadeMux I__1344 (
            .O(N__15813),
            .I(\b2v_inst36.count_rst_7_cascade_ ));
    CascadeMux I__1343 (
            .O(N__15810),
            .I(\b2v_inst36.countZ0Z_6_cascade_ ));
    InMux I__1342 (
            .O(N__15807),
            .I(N__15801));
    InMux I__1341 (
            .O(N__15806),
            .I(N__15801));
    LocalMux I__1340 (
            .O(N__15801),
            .I(\b2v_inst36.count_2_4 ));
    CascadeMux I__1339 (
            .O(N__15798),
            .I(\b2v_inst36.countZ0Z_11_cascade_ ));
    InMux I__1338 (
            .O(N__15795),
            .I(N__15792));
    LocalMux I__1337 (
            .O(N__15792),
            .I(\b2v_inst36.count_2_11 ));
    CascadeMux I__1336 (
            .O(N__15789),
            .I(N__15785));
    CascadeMux I__1335 (
            .O(N__15788),
            .I(N__15782));
    InMux I__1334 (
            .O(N__15785),
            .I(N__15777));
    InMux I__1333 (
            .O(N__15782),
            .I(N__15777));
    LocalMux I__1332 (
            .O(N__15777),
            .I(\b2v_inst36.count_2_6 ));
    CascadeMux I__1331 (
            .O(N__15774),
            .I(\b2v_inst36.countZ0Z_10_cascade_ ));
    InMux I__1330 (
            .O(N__15771),
            .I(N__15768));
    LocalMux I__1329 (
            .O(N__15768),
            .I(\b2v_inst36.count_2_10 ));
    InMux I__1328 (
            .O(N__15765),
            .I(N__15762));
    LocalMux I__1327 (
            .O(N__15762),
            .I(\b2v_inst36.count_rst_9 ));
    CascadeMux I__1326 (
            .O(N__15759),
            .I(\b2v_inst36.count_rst_9_cascade_ ));
    CascadeMux I__1325 (
            .O(N__15756),
            .I(\b2v_inst36.un2_count_1_axb_5_cascade_ ));
    InMux I__1324 (
            .O(N__15753),
            .I(N__15747));
    InMux I__1323 (
            .O(N__15752),
            .I(N__15747));
    LocalMux I__1322 (
            .O(N__15747),
            .I(\b2v_inst36.count_2_5 ));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(\b2v_inst6.un2_count_1_cry_8 ),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\b2v_inst5.un2_count_1_cry_7 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(\b2v_inst36.un2_count_1_cry_8 ),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_8 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_16 ),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(b2v_inst20_un4_counter_7),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_8 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_16 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_24 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(\b2v_inst16.un4_count_1_cry_8 ),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_0_cry_7 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz0 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(\b2v_inst11.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_16_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_94_cry_7_s1 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_94_cry_7_s0 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\b2v_inst11.un1_count_cry_8 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\b2v_inst11.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_1_cry_8 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_12_0_));
    ICE_GB \b2v_inst200.count_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__19860),
            .GLOBALBUFFEROUTPUT(\b2v_inst200.count_en_g ));
    ICE_GB N_607_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__35828),
            .GLOBALBUFFEROUTPUT(N_607_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \b2v_inst36.count_RNIJKUH1_0_5_LC_1_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJKUH1_0_5_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJKUH1_0_5_LC_1_1_0 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \b2v_inst36.count_RNIJKUH1_0_5_LC_1_1_0  (
            .in0(N__15765),
            .in1(N__15753),
            .in2(N__16341),
            .in3(N__16990),
            .lcout(\b2v_inst36.un12_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI4VQN1_10_LC_1_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI4VQN1_10_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI4VQN1_10_LC_1_1_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNI4VQN1_10_LC_1_1_1  (
            .in0(N__16989),
            .in1(N__15771),
            .in2(_gnd_net_),
            .in3(N__15837),
            .lcout(\b2v_inst36.countZ0Z_10 ),
            .ltout(\b2v_inst36.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_10_LC_1_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_10_LC_1_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_10_LC_1_1_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_10_LC_1_1_2  (
            .in0(N__19525),
            .in1(N__16584),
            .in2(N__15774),
            .in3(N__19070),
            .lcout(\b2v_inst36.count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36942),
            .ce(N__17012),
            .sr(N__19557));
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_1_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_1_1_3 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_1_1_3  (
            .in0(N__19068),
            .in1(N__16386),
            .in2(N__19543),
            .in3(N__16373),
            .lcout(\b2v_inst36.count_rst_9 ),
            .ltout(\b2v_inst36.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIJKUH1_5_LC_1_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJKUH1_5_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJKUH1_5_LC_1_1_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIJKUH1_5_LC_1_1_4  (
            .in0(_gnd_net_),
            .in1(N__15752),
            .in2(N__15759),
            .in3(N__16987),
            .lcout(\b2v_inst36.un2_count_1_axb_5 ),
            .ltout(\b2v_inst36.un2_count_1_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_5_LC_1_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_5_LC_1_1_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_5_LC_1_1_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_5_LC_1_1_5  (
            .in0(N__19069),
            .in1(N__16374),
            .in2(N__15756),
            .in3(N__19526),
            .lcout(\b2v_inst36.count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36942),
            .ce(N__17012),
            .sr(N__19557));
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_1_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_1_1_6 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_1_1_6  (
            .in0(N__19524),
            .in1(N__16310),
            .in2(N__19083),
            .in3(N__16337),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNINQ0I1_7_LC_1_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNINQ0I1_7_LC_1_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNINQ0I1_7_LC_1_1_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNINQ0I1_7_LC_1_1_7  (
            .in0(N__16988),
            .in1(_gnd_net_),
            .in2(N__15813),
            .in3(N__16506),
            .lcout(\b2v_inst36.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_6_LC_1_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_6_LC_1_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_6_LC_1_2_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst36.count_6_LC_1_2_0  (
            .in0(N__16356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19509),
            .lcout(\b2v_inst36.count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36898),
            .ce(N__17001),
            .sr(N__19541));
    defparam \b2v_inst36.count_RNIHHTH1_4_LC_1_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIHHTH1_4_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIHHTH1_4_LC_1_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIHHTH1_4_LC_1_2_1  (
            .in0(N__15806),
            .in1(N__16982),
            .in2(_gnd_net_),
            .in3(N__16402),
            .lcout(\b2v_inst36.un2_count_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_4_LC_1_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_4_LC_1_2_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_4_LC_1_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_4_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16404),
            .lcout(\b2v_inst36.count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36898),
            .ce(N__17001),
            .sr(N__19541));
    defparam \b2v_inst36.count_RNILNVH1_6_LC_1_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNILNVH1_6_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNILNVH1_6_LC_1_2_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst36.count_RNILNVH1_6_LC_1_2_3  (
            .in0(N__19507),
            .in1(N__16985),
            .in2(N__15789),
            .in3(N__16355),
            .lcout(),
            .ltout(\b2v_inst36.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI69T33_4_LC_1_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI69T33_4_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI69T33_4_LC_1_2_4 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst36.count_RNI69T33_4_LC_1_2_4  (
            .in0(N__16986),
            .in1(N__16403),
            .in2(N__15810),
            .in3(N__15807),
            .lcout(\b2v_inst36.un12_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIDPQG1_11_LC_1_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIDPQG1_11_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIDPQG1_11_LC_1_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIDPQG1_11_LC_1_2_5  (
            .in0(N__15795),
            .in1(N__16984),
            .in2(_gnd_net_),
            .in3(N__15828),
            .lcout(\b2v_inst36.countZ0Z_11 ),
            .ltout(\b2v_inst36.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_11_LC_1_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_11_LC_1_2_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_11_LC_1_2_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst36.count_11_LC_1_2_6  (
            .in0(N__19080),
            .in1(N__19508),
            .in2(N__15798),
            .in3(N__16539),
            .lcout(\b2v_inst36.count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36898),
            .ce(N__17001),
            .sr(N__19541));
    defparam \b2v_inst36.count_RNILNVH1_0_6_LC_1_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNILNVH1_0_6_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNILNVH1_0_6_LC_1_2_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst36.count_RNILNVH1_0_6_LC_1_2_7  (
            .in0(N__19506),
            .in1(N__16983),
            .in2(N__15788),
            .in3(N__16354),
            .lcout(\b2v_inst36.un2_count_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIPT1I1_0_8_LC_1_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPT1I1_0_8_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPT1I1_0_8_LC_1_3_0 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \b2v_inst36.count_RNIPT1I1_0_8_LC_1_3_0  (
            .in0(N__15858),
            .in1(N__15846),
            .in2(N__16611),
            .in3(N__16992),
            .lcout(\b2v_inst36.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_1_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_1_3_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_1_3_1  (
            .in0(N__19456),
            .in1(N__16644),
            .in2(N__16629),
            .in3(N__19020),
            .lcout(\b2v_inst36.count_rst_6 ),
            .ltout(\b2v_inst36.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIPT1I1_8_LC_1_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPT1I1_8_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPT1I1_8_LC_1_3_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIPT1I1_8_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__15845),
            .in2(N__15852),
            .in3(N__16991),
            .lcout(\b2v_inst36.un2_count_1_axb_8 ),
            .ltout(\b2v_inst36.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_8_LC_1_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_8_LC_1_3_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_8_LC_1_3_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst36.count_8_LC_1_3_3  (
            .in0(N__16628),
            .in1(N__19445),
            .in2(N__15849),
            .in3(N__19025),
            .lcout(\b2v_inst36.count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36889),
            .ce(N__17013),
            .sr(N__19505));
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_1_3_4 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_1_3_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_1_3_4  (
            .in0(N__19021),
            .in1(N__16610),
            .in2(N__16583),
            .in3(N__19457),
            .lcout(\b2v_inst36.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIRQCA_0_LC_1_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIRQCA_0_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIRQCA_0_LC_1_3_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst36.count_RNIRQCA_0_LC_1_3_5  (
            .in0(N__16705),
            .in1(N__19444),
            .in2(_gnd_net_),
            .in3(N__19019),
            .lcout(\b2v_inst36.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_1_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_1_3_6 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_1_3_6  (
            .in0(N__16559),
            .in1(N__19458),
            .in2(N__19060),
            .in3(N__16538),
            .lcout(\b2v_inst36.count_rst_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI2GG91_1_LC_1_4_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI2GG91_1_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI2GG91_1_LC_1_4_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNI2GG91_1_LC_1_4_0  (
            .in0(N__15881),
            .in1(N__16915),
            .in2(_gnd_net_),
            .in3(N__15822),
            .lcout(\b2v_inst36.un2_count_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIRQCA_1_LC_1_4_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIRQCA_1_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIRQCA_1_LC_1_4_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst36.count_RNIRQCA_1_LC_1_4_1  (
            .in0(N__16495),
            .in1(N__16700),
            .in2(_gnd_net_),
            .in3(N__19467),
            .lcout(\b2v_inst36.count_rst_13 ),
            .ltout(\b2v_inst36.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI2GG91_0_1_LC_1_4_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI2GG91_0_1_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI2GG91_0_1_LC_1_4_2 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \b2v_inst36.count_RNI2GG91_0_1_LC_1_4_2  (
            .in0(N__15882),
            .in1(N__16916),
            .in2(N__15816),
            .in3(N__16560),
            .lcout(),
            .ltout(\b2v_inst36.un12_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIRDCV5_1_LC_1_4_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIRDCV5_1_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIRDCV5_1_LC_1_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNIRDCV5_1_LC_1_4_3  (
            .in0(N__16281),
            .in1(N__15930),
            .in2(N__15924),
            .in3(N__15921),
            .lcout(),
            .ltout(\b2v_inst36.un12_clk_100khz_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNISNCLA_4_LC_1_4_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNISNCLA_4_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNISNCLA_4_LC_1_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNISNCLA_4_LC_1_4_4  (
            .in0(N__15912),
            .in1(N__16722),
            .in2(N__15903),
            .in3(N__16677),
            .lcout(\b2v_inst36.N_1_i ),
            .ltout(\b2v_inst36.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_0_LC_1_4_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_0_LC_1_4_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_0_LC_1_4_5 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst36.count_0_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(N__16701),
            .in2(N__15900),
            .in3(N__19559),
            .lcout(\b2v_inst36.count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37101),
            .ce(N__16944),
            .sr(N__19558));
    defparam \b2v_inst36.count_RNI1FG91_0_LC_1_4_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI1FG91_0_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI1FG91_0_LC_1_4_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNI1FG91_0_LC_1_4_6  (
            .in0(N__15897),
            .in1(N__16914),
            .in2(_gnd_net_),
            .in3(N__15891),
            .lcout(\b2v_inst36.countZ0Z_0 ),
            .ltout(\b2v_inst36.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_1_LC_1_4_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_1_LC_1_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_1_LC_1_4_7 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \b2v_inst36.count_1_LC_1_4_7  (
            .in0(N__16496),
            .in1(_gnd_net_),
            .in2(N__15885),
            .in3(N__19560),
            .lcout(\b2v_inst36.count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37101),
            .ce(N__16944),
            .sr(N__19558));
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_5_0 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_5_0 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_5_0  (
            .in0(N__17062),
            .in1(N__17045),
            .in2(N__19806),
            .in3(N__17476),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIV7UA_11_LC_1_5_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIV7UA_11_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIV7UA_11_LC_1_5_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst16.count_RNIV7UA_11_LC_1_5_1  (
            .in0(N__19222),
            .in1(_gnd_net_),
            .in2(N__15873),
            .in3(N__15867),
            .lcout(\b2v_inst16.countZ0Z_11 ),
            .ltout(\b2v_inst16.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_11_LC_1_5_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_11_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_11_LC_1_5_2 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst16.count_11_LC_1_5_2  (
            .in0(N__19803),
            .in1(N__17046),
            .in2(N__15870),
            .in3(N__17479),
            .lcout(\b2v_inst16.count_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37108),
            .ce(N__19256),
            .sr(N__19141));
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_5_3 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_5_3 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_5_3  (
            .in0(N__17475),
            .in1(N__19802),
            .in2(N__17217),
            .in3(N__17233),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNITRJU_4_LC_1_5_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNITRJU_4_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNITRJU_4_LC_1_5_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst16.count_RNITRJU_4_LC_1_5_4  (
            .in0(N__15963),
            .in1(_gnd_net_),
            .in2(N__15969),
            .in3(N__19221),
            .lcout(\b2v_inst16.countZ0Z_4 ),
            .ltout(\b2v_inst16.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_4_LC_1_5_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_4_LC_1_5_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_4_LC_1_5_5 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_4_LC_1_5_5  (
            .in0(N__17478),
            .in1(N__19805),
            .in2(N__15966),
            .in3(N__17216),
            .lcout(\b2v_inst16.count_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37108),
            .ce(N__19256),
            .sr(N__19141));
    defparam \b2v_inst16.count_RNIROIU_3_LC_1_5_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIROIU_3_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIROIU_3_LC_1_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIROIU_3_LC_1_5_6  (
            .in0(N__15954),
            .in1(N__16032),
            .in2(_gnd_net_),
            .in3(N__19223),
            .lcout(\b2v_inst16.countZ0Z_3 ),
            .ltout(\b2v_inst16.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_3_LC_1_5_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_3_LC_1_5_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_3_LC_1_5_7 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_3_LC_1_5_7  (
            .in0(N__17477),
            .in1(N__19804),
            .in2(N__15957),
            .in3(N__17249),
            .lcout(\b2v_inst16.count_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37108),
            .ce(N__19256),
            .sr(N__19141));
    defparam \b2v_inst16.count_RNI_10_LC_1_6_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_10_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_10_LC_1_6_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst16.count_RNI_10_LC_1_6_0  (
            .in0(N__17412),
            .in1(N__18915),
            .in2(N__18870),
            .in3(N__17327),
            .lcout(\b2v_inst16.count_4_i_a3_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_15_LC_1_6_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_15_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_15_LC_1_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst16.count_RNI_15_LC_1_6_1  (
            .in0(N__17358),
            .in1(N__16791),
            .in2(N__18957),
            .in3(N__17148),
            .lcout(\b2v_inst16.count_4_i_a3_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_3_LC_1_6_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_3_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_3_LC_1_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst16.count_RNI_3_LC_1_6_2  (
            .in0(N__17270),
            .in1(N__17195),
            .in2(N__17133),
            .in3(N__17234),
            .lcout(),
            .ltout(\b2v_inst16.count_4_i_a3_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIE4RF_3_1_LC_1_6_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIE4RF_3_1_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIE4RF_3_1_LC_1_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst16.count_RNIE4RF_3_1_LC_1_6_3  (
            .in0(N__15996),
            .in1(N__15948),
            .in2(N__15942),
            .in3(N__15939),
            .lcout(\b2v_inst16.N_414 ),
            .ltout(\b2v_inst16.N_414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_0_LC_1_6_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_LC_1_6_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst16.count_RNI_0_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15933),
            .in3(N__16809),
            .lcout(\b2v_inst16.N_416 ),
            .ltout(\b2v_inst16.N_416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_6_5 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_6_5 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_6_5  (
            .in0(N__19780),
            .in1(N__17271),
            .in2(N__16035),
            .in3(N__17250),
            .lcout(\b2v_inst16.count_rst_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIE4RF_2_1_LC_1_7_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIE4RF_2_1_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIE4RF_2_1_LC_1_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst16.count_RNIE4RF_2_1_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__16810),
            .in2(_gnd_net_),
            .in3(N__16827),
            .lcout(\b2v_inst16.count_RNIE4RF_2Z0Z_1 ),
            .ltout(\b2v_inst16.count_RNIE4RF_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIE4RF_1_LC_1_7_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIE4RF_1_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIE4RF_1_LC_1_7_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \b2v_inst16.count_RNIE4RF_1_LC_1_7_1  (
            .in0(N__19779),
            .in1(N__15980),
            .in2(N__16026),
            .in3(N__19275),
            .lcout(\b2v_inst16.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_0_0_LC_1_7_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_0_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_0_LC_1_7_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst16.count_RNI_0_0_LC_1_7_2  (
            .in0(N__16019),
            .in1(N__19775),
            .in2(_gnd_net_),
            .in3(N__16811),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNID3RF_0_LC_1_7_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNID3RF_0_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNID3RF_0_LC_1_7_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst16.count_RNID3RF_0_LC_1_7_3  (
            .in0(N__19241),
            .in1(_gnd_net_),
            .in2(N__16023),
            .in3(N__16008),
            .lcout(\b2v_inst16.countZ0Z_0 ),
            .ltout(\b2v_inst16.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_0_LC_1_7_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_0_LC_1_7_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_0_LC_1_7_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst16.count_0_LC_1_7_4  (
            .in0(N__16020),
            .in1(_gnd_net_),
            .in2(N__16011),
            .in3(N__19778),
            .lcout(\b2v_inst16.count_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37109),
            .ce(N__19274),
            .sr(N__19130));
    defparam \b2v_inst16.count_RNIE4RF_1_1_LC_1_7_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIE4RF_1_1_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIE4RF_1_1_LC_1_7_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst16.count_RNIE4RF_1_1_LC_1_7_5  (
            .in0(N__17295),
            .in1(N__16002),
            .in2(_gnd_net_),
            .in3(N__17069),
            .lcout(\b2v_inst16.count_4_i_a3_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIE4RF_0_1_LC_1_7_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIE4RF_0_1_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIE4RF_0_1_LC_1_7_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst16.count_RNIE4RF_0_1_LC_1_7_6  (
            .in0(N__15989),
            .in1(N__19776),
            .in2(N__15981),
            .in3(N__19240),
            .lcout(\b2v_inst16.un4_count_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_1_LC_1_7_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_1_LC_1_7_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_1_LC_1_7_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \b2v_inst16.count_1_LC_1_7_7  (
            .in0(N__19777),
            .in1(N__15990),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37109),
            .ce(N__19274),
            .sr(N__19130));
    defparam \b2v_inst16.count_RNI35NU_7_LC_1_8_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI35NU_7_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI35NU_7_LC_1_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNI35NU_7_LC_1_8_0  (
            .in0(N__19242),
            .in1(N__16068),
            .in2(_gnd_net_),
            .in3(N__16041),
            .lcout(\b2v_inst16.countZ0Z_7 ),
            .ltout(\b2v_inst16.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_7_LC_1_8_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_7_LC_1_8_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_7_LC_1_8_1 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst16.count_7_LC_1_8_1  (
            .in0(N__19768),
            .in1(N__17493),
            .in2(N__16071),
            .in3(N__17097),
            .lcout(\b2v_inst16.count_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37139),
            .ce(N__19273),
            .sr(N__19137));
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_8_2 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_8_2 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_8_2  (
            .in0(N__17490),
            .in1(N__17188),
            .in2(N__17172),
            .in3(N__19767),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIVUKU_5_LC_1_8_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIVUKU_5_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIVUKU_5_LC_1_8_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIVUKU_5_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__16056),
            .in2(N__16062),
            .in3(N__19243),
            .lcout(\b2v_inst16.countZ0Z_5 ),
            .ltout(\b2v_inst16.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_5_LC_1_8_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_5_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_5_LC_1_8_4 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst16.count_5_LC_1_8_4  (
            .in0(N__17491),
            .in1(N__17171),
            .in2(N__16059),
            .in3(N__19770),
            .lcout(\b2v_inst16.count_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37139),
            .ce(N__19273),
            .sr(N__19137));
    defparam \b2v_inst16.count_RNI58OU_8_LC_1_8_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI58OU_8_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI58OU_8_LC_1_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNI58OU_8_LC_1_8_5  (
            .in0(N__16047),
            .in1(N__17304),
            .in2(_gnd_net_),
            .in3(N__19244),
            .lcout(\b2v_inst16.countZ0Z_8 ),
            .ltout(\b2v_inst16.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_8_LC_1_8_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_8_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_8_LC_1_8_6 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_8_LC_1_8_6  (
            .in0(N__17492),
            .in1(N__19769),
            .in2(N__16050),
            .in3(N__17346),
            .lcout(\b2v_inst16.count_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37139),
            .ce(N__19273),
            .sr(N__19137));
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_8_7 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_8_7 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_8_7  (
            .in0(N__19766),
            .in1(N__17489),
            .in2(N__17122),
            .in3(N__17096),
            .lcout(\b2v_inst16.count_rst_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIBO6I1_1_0_LC_1_9_0 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIBO6I1_1_0_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIBO6I1_1_0_LC_1_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.curr_state_RNIBO6I1_1_0_LC_1_9_0  (
            .in0(N__20477),
            .in1(N__19829),
            .in2(_gnd_net_),
            .in3(N__17487),
            .lcout(),
            .ltout(\b2v_inst16.curr_state_7_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI4KJ02_1_LC_1_9_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI4KJ02_1_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI4KJ02_1_LC_1_9_1 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \b2v_inst16.curr_state_RNI4KJ02_1_LC_1_9_1  (
            .in0(N__28397),
            .in1(_gnd_net_),
            .in2(N__16122),
            .in3(N__16095),
            .lcout(\b2v_inst16.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_1_9_2 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_1_9_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_1_9_2  (
            .in0(N__38529),
            .in1(N__16119),
            .in2(_gnd_net_),
            .in3(N__34833),
            .lcout(\b2v_inst16.N_208_0 ),
            .ltout(\b2v_inst16.N_208_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIBO6I1_0_LC_1_9_3 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIBO6I1_0_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIBO6I1_0_LC_1_9_3 .LUT_INIT=16'b1010111111111111;
    LogicCell40 \b2v_inst16.curr_state_RNIBO6I1_0_LC_1_9_3  (
            .in0(N__28395),
            .in1(_gnd_net_),
            .in2(N__16101),
            .in3(N__16089),
            .lcout(\b2v_inst16.curr_state_RNIBO6I1Z0Z_0 ),
            .ltout(\b2v_inst16.curr_state_RNIBO6I1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_1_LC_1_9_4 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_LC_1_9_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_1_LC_1_9_4 .LUT_INIT=16'b0000001111001111;
    LogicCell40 \b2v_inst16.curr_state_1_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__20475),
            .in2(N__16098),
            .in3(N__17488),
            .lcout(\b2v_inst16.curr_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37125),
            .ce(N__27542),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIU6GN_7_LC_1_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_1_9_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst11.count_RNIU6GN_7_LC_1_9_5  (
            .in0(N__28396),
            .in1(_gnd_net_),
            .in2(N__16083),
            .in3(N__16152),
            .lcout(\b2v_inst11.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_0_LC_1_9_7 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_0_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_0_LC_1_9_7 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \b2v_inst16.curr_state_0_LC_1_9_7  (
            .in0(N__20476),
            .in1(N__20519),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37125),
            .ce(N__27542),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_8_LC_1_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_8_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_8_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_8_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17622),
            .lcout(\b2v_inst11.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37141),
            .ce(N__27540),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_7_LC_1_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_7_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_7_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_7_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16151),
            .lcout(\b2v_inst11.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37141),
            .ce(N__27540),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_LC_1_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__20084),
            .in2(N__17663),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\b2v_inst11.un1_count_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_11_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_11_1  (
            .in0(N__20058),
            .in1(N__18262),
            .in2(_gnd_net_),
            .in3(N__16074),
            .lcout(\b2v_inst11.count_1_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_1_cZ0 ),
            .carryout(\b2v_inst11.un1_count_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_11_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_11_2  (
            .in0(N__20050),
            .in1(_gnd_net_),
            .in2(N__18245),
            .in3(N__16164),
            .lcout(\b2v_inst11.count_1_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_2_cZ0 ),
            .carryout(\b2v_inst11.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_11_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_11_3  (
            .in0(N__20059),
            .in1(_gnd_net_),
            .in2(N__18221),
            .in3(N__16161),
            .lcout(\b2v_inst11.count_1_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_3 ),
            .carryout(\b2v_inst11.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_11_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_11_4  (
            .in0(N__20051),
            .in1(_gnd_net_),
            .in2(N__18138),
            .in3(N__16158),
            .lcout(\b2v_inst11.count_1_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_4 ),
            .carryout(\b2v_inst11.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_11_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_11_5  (
            .in0(N__20060),
            .in1(_gnd_net_),
            .in2(N__18165),
            .in3(N__16155),
            .lcout(\b2v_inst11.count_1_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_5 ),
            .carryout(\b2v_inst11.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_11_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_11_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_11_6  (
            .in0(N__20052),
            .in1(_gnd_net_),
            .in2(N__18196),
            .in3(N__16137),
            .lcout(\b2v_inst11.count_1_7 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_6 ),
            .carryout(\b2v_inst11.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_11_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_11_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_11_7  (
            .in0(N__20061),
            .in1(_gnd_net_),
            .in2(N__17941),
            .in3(N__16134),
            .lcout(\b2v_inst11.count_1_8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_7 ),
            .carryout(\b2v_inst11.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_12_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_12_0  (
            .in0(N__20053),
            .in1(_gnd_net_),
            .in2(N__17911),
            .in3(N__16131),
            .lcout(\b2v_inst11.count_1_9 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\b2v_inst11.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_12_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_12_1  (
            .in0(N__20062),
            .in1(_gnd_net_),
            .in2(N__18106),
            .in3(N__16128),
            .lcout(\b2v_inst11.count_1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_9 ),
            .carryout(\b2v_inst11.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_12_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_12_2  (
            .in0(N__20054),
            .in1(_gnd_net_),
            .in2(N__18046),
            .in3(N__16125),
            .lcout(\b2v_inst11.count_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_10 ),
            .carryout(\b2v_inst11.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_12_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_12_3  (
            .in0(N__20063),
            .in1(_gnd_net_),
            .in2(N__18077),
            .in3(N__16212),
            .lcout(\b2v_inst11.count_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_11 ),
            .carryout(\b2v_inst11.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_12_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_12_4  (
            .in0(N__20055),
            .in1(_gnd_net_),
            .in2(N__18022),
            .in3(N__16209),
            .lcout(\b2v_inst11.count_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_12 ),
            .carryout(\b2v_inst11.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_12_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_12_5  (
            .in0(N__20064),
            .in1(_gnd_net_),
            .in2(N__17999),
            .in3(N__16206),
            .lcout(\b2v_inst11.count_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_13 ),
            .carryout(\b2v_inst11.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_12_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_12_6  (
            .in0(N__20056),
            .in1(N__17972),
            .in2(_gnd_net_),
            .in3(N__16203),
            .lcout(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQF4M_14_LC_1_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_1_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIQF4M_14_LC_1_12_7  (
            .in0(N__16170),
            .in1(N__28409),
            .in2(_gnd_net_),
            .in3(N__16181),
            .lcout(\b2v_inst11.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_1_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_1_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIQ0EN_5_LC_1_13_0  (
            .in0(N__28406),
            .in1(N__16188),
            .in2(_gnd_net_),
            .in3(N__16199),
            .lcout(\b2v_inst11.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_5_LC_1_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_5_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_5_LC_1_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_5_LC_1_13_1  (
            .in0(N__16200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37148),
            .ce(N__27533),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_14_LC_1_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_14_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_14_LC_1_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_14_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16182),
            .lcout(\b2v_inst11.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37148),
            .ce(N__27533),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIS3FN_6_LC_1_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_1_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIS3FN_6_LC_1_13_4  (
            .in0(N__28407),
            .in1(N__16236),
            .in2(_gnd_net_),
            .in3(N__16247),
            .lcout(\b2v_inst11.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_6_LC_1_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_6_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_6_LC_1_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_6_LC_1_13_5  (
            .in0(N__16248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37148),
            .ce(N__27533),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNISI5M_15_LC_1_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNISI5M_15_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNISI5M_15_LC_1_13_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNISI5M_15_LC_1_13_6  (
            .in0(N__28408),
            .in1(N__16218),
            .in2(_gnd_net_),
            .in3(N__16226),
            .lcout(\b2v_inst11.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_15_LC_1_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_15_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_15_LC_1_13_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_15_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16230),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37148),
            .ce(N__27533),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_0_c_LC_1_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_0_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_0_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_0_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__17529),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_1_c_inv_LC_1_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_1_c_inv_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_1_c_inv_LC_1_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_1_c_inv_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__17816),
            .in2(N__17804),
            .in3(N__17667),
            .lcout(\b2v_inst11.N_5853_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_0 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_2_c_inv_LC_1_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_2_c_inv_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_2_c_inv_LC_1_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_2_c_inv_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__17786),
            .in2(N__17775),
            .in3(N__18269),
            .lcout(\b2v_inst11.N_5854_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_1 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_3_c_inv_LC_1_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_3_c_inv_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_3_c_inv_LC_1_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_3_c_inv_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__18485),
            .in2(N__18473),
            .in3(N__18246),
            .lcout(\b2v_inst11.N_5855_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_2 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_4_c_inv_LC_1_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_4_c_inv_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_4_c_inv_LC_1_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_4_c_inv_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__18437),
            .in2(N__18456),
            .in3(N__18222),
            .lcout(\b2v_inst11.N_5856_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_3 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_5_c_inv_LC_1_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_5_c_inv_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_5_c_inv_LC_1_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_5_c_inv_LC_1_14_5  (
            .in0(N__18130),
            .in1(N__18425),
            .in2(N__18414),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5857_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_4 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_6_c_inv_LC_1_14_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_6_c_inv_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_6_c_inv_LC_1_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_6_c_inv_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__18392),
            .in2(N__18380),
            .in3(N__18160),
            .lcout(\b2v_inst11.N_5858_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_5 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_7_c_inv_LC_1_14_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_7_c_inv_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_7_c_inv_LC_1_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_7_c_inv_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__18359),
            .in2(N__18348),
            .in3(N__18197),
            .lcout(\b2v_inst11.N_5859_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_6 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_8_c_inv_LC_1_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_8_c_inv_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_8_c_inv_LC_1_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_8_c_inv_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__18332),
            .in2(N__18320),
            .in3(N__17946),
            .lcout(\b2v_inst11.N_5860_i ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_9_c_inv_LC_1_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_9_c_inv_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_9_c_inv_LC_1_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_9_c_inv_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__18302),
            .in2(N__18291),
            .in3(N__17916),
            .lcout(\b2v_inst11.N_5861_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_8 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_10_c_inv_LC_1_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_10_c_inv_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_10_c_inv_LC_1_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_10_c_inv_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__18680),
            .in2(N__18669),
            .in3(N__18111),
            .lcout(\b2v_inst11.N_5862_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_9 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_11_c_inv_LC_1_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_11_c_inv_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_11_c_inv_LC_1_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_11_c_inv_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__18644),
            .in2(N__18633),
            .in3(N__18053),
            .lcout(\b2v_inst11.N_5863_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_10 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_12_c_inv_LC_1_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_12_c_inv_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_12_c_inv_LC_1_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_12_c_inv_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__18611),
            .in2(N__18600),
            .in3(N__18081),
            .lcout(\b2v_inst11.N_5864_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_11 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_13_c_inv_LC_1_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_13_c_inv_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_13_c_inv_LC_1_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_13_c_inv_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__18567),
            .in2(N__18584),
            .in3(N__18023),
            .lcout(\b2v_inst11.N_5865_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_12 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_14_c_inv_LC_1_15_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_14_c_inv_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_14_c_inv_LC_1_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_14_c_inv_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__18533),
            .in2(N__18552),
            .in3(N__18000),
            .lcout(\b2v_inst11.N_5866_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_13 ),
            .carryout(\b2v_inst11.un85_clk_100khz_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_15_c_inv_LC_1_15_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_15_c_inv_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_15_c_inv_LC_1_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_15_c_inv_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__18503),
            .in2(N__18521),
            .in3(N__17973),
            .lcout(\b2v_inst11.N_5867_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_0_cry_14 ),
            .carryout(\b2v_inst11.un85_clk_100khz0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz0_THRU_LUT4_0_LC_1_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz0_THRU_LUT4_0_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz0_THRU_LUT4_0_LC_1_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz0_THRU_LUT4_0_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16296),
            .lcout(\b2v_inst11.un85_clk_100khz0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_2_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_2_1_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_2_1_0  (
            .in0(N__19468),
            .in1(N__16457),
            .in2(N__16479),
            .in3(N__19061),
            .lcout(\b2v_inst36.count_rst_12 ),
            .ltout(\b2v_inst36.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIDBRH1_2_LC_2_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIDBRH1_2_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIDBRH1_2_LC_2_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIDBRH1_2_LC_2_1_1  (
            .in0(_gnd_net_),
            .in1(N__16262),
            .in2(N__16293),
            .in3(N__16945),
            .lcout(\b2v_inst36.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIFESH1_3_LC_2_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIFESH1_3_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIFESH1_3_LC_2_1_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNIFESH1_3_LC_2_1_2  (
            .in0(N__16946),
            .in1(N__16254),
            .in2(_gnd_net_),
            .in3(N__16269),
            .lcout(\b2v_inst36.countZ0Z_3 ),
            .ltout(\b2v_inst36.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIDBRH1_0_2_LC_2_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIDBRH1_0_2_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIDBRH1_0_2_LC_2_1_3 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \b2v_inst36.count_RNIDBRH1_0_2_LC_2_1_3  (
            .in0(N__16290),
            .in1(N__16263),
            .in2(N__16284),
            .in3(N__16947),
            .lcout(\b2v_inst36.un12_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_2_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_2_1_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_2_1_4  (
            .in0(N__19469),
            .in1(N__19062),
            .in2(N__16430),
            .in3(N__16446),
            .lcout(\b2v_inst36.count_rst_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_2_LC_2_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_2_LC_2_1_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_2_LC_2_1_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst36.count_2_LC_2_1_5  (
            .in0(N__19063),
            .in1(N__16478),
            .in2(N__16461),
            .in3(N__19549),
            .lcout(\b2v_inst36.count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36801),
            .ce(N__17011),
            .sr(N__19547));
    defparam \b2v_inst36.count_3_LC_2_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_3_LC_2_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_3_LC_2_1_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst36.count_3_LC_2_1_6  (
            .in0(N__19470),
            .in1(N__19064),
            .in2(N__16431),
            .in3(N__16445),
            .lcout(\b2v_inst36.count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36801),
            .ce(N__17011),
            .sr(N__19547));
    defparam \b2v_inst36.count_7_LC_2_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_7_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_7_LC_2_1_7 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst36.count_7_LC_2_1_7  (
            .in0(N__16311),
            .in1(N__16336),
            .in2(N__19081),
            .in3(N__19548),
            .lcout(\b2v_inst36.count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36801),
            .ce(N__17011),
            .sr(N__19547));
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_2_2_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_2_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__16707),
            .in2(N__16500),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_2_2_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_2_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__16474),
            .in2(_gnd_net_),
            .in3(N__16449),
            .lcout(\b2v_inst36.un2_count_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_1 ),
            .carryout(\b2v_inst36.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_2_2_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_2_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_2_2_2  (
            .in0(_gnd_net_),
            .in1(N__16444),
            .in2(_gnd_net_),
            .in3(N__16416),
            .lcout(\b2v_inst36.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_2 ),
            .carryout(\b2v_inst36.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_2_2_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_2_2_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_2_2_3  (
            .in0(N__19471),
            .in1(_gnd_net_),
            .in2(N__16413),
            .in3(N__16389),
            .lcout(\b2v_inst36.count_rst_10 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_3 ),
            .carryout(\b2v_inst36.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_2_2_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_2_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_2_2_4  (
            .in0(_gnd_net_),
            .in1(N__16385),
            .in2(_gnd_net_),
            .in3(N__16365),
            .lcout(\b2v_inst36.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_4 ),
            .carryout(\b2v_inst36.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_2_2_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_2_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_2_2_5  (
            .in0(_gnd_net_),
            .in1(N__16362),
            .in2(_gnd_net_),
            .in3(N__16344),
            .lcout(\b2v_inst36.un2_count_1_cry_5_c_RNIE2FZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_5 ),
            .carryout(\b2v_inst36.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_2_2_6 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_2_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_2_2_6  (
            .in0(_gnd_net_),
            .in1(N__16332),
            .in2(_gnd_net_),
            .in3(N__16299),
            .lcout(\b2v_inst36.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_6 ),
            .carryout(\b2v_inst36.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_2_2_7 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_2_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_2_2_7  (
            .in0(_gnd_net_),
            .in1(N__16640),
            .in2(_gnd_net_),
            .in3(N__16617),
            .lcout(\b2v_inst36.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_7 ),
            .carryout(\b2v_inst36.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_2_3_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_2_3_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_2_3_0  (
            .in0(N__19459),
            .in1(N__16512),
            .in2(_gnd_net_),
            .in3(N__16614),
            .lcout(\b2v_inst36.count_rst_5 ),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_2_3_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_2_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_2_3_1  (
            .in0(_gnd_net_),
            .in1(N__16606),
            .in2(_gnd_net_),
            .in3(N__16563),
            .lcout(\b2v_inst36.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_9 ),
            .carryout(\b2v_inst36.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_2_3_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_2_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_2_3_2  (
            .in0(_gnd_net_),
            .in1(N__16555),
            .in2(_gnd_net_),
            .in3(N__16527),
            .lcout(\b2v_inst36.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_10 ),
            .carryout(\b2v_inst36.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIM01C_LC_2_3_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIM01C_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIM01C_LC_2_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_11_c_RNIM01C_LC_2_3_3  (
            .in0(N__19462),
            .in1(N__16761),
            .in2(_gnd_net_),
            .in3(N__16524),
            .lcout(\b2v_inst36.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_11 ),
            .carryout(\b2v_inst36.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_2_3_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_2_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_2_3_4  (
            .in0(N__19460),
            .in1(N__16655),
            .in2(_gnd_net_),
            .in3(N__16521),
            .lcout(\b2v_inst36.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_12 ),
            .carryout(\b2v_inst36.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_2_3_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_2_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_2_3_5  (
            .in0(N__19463),
            .in1(N__16716),
            .in2(_gnd_net_),
            .in3(N__16518),
            .lcout(\b2v_inst36.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_13 ),
            .carryout(\b2v_inst36.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_2_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_2_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_2_3_6  (
            .in0(N__19461),
            .in1(N__16845),
            .in2(_gnd_net_),
            .in3(N__16515),
            .lcout(\b2v_inst36.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIR03I1_9_LC_2_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIR03I1_9_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIR03I1_9_LC_2_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIR03I1_9_LC_2_3_7  (
            .in0(N__16733),
            .in1(N__16993),
            .in2(_gnd_net_),
            .in3(N__16753),
            .lcout(\b2v_inst36.un2_count_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_12_LC_2_4_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_12_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_12_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_12_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16770),
            .lcout(\b2v_inst36.count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37027),
            .ce(N__16943),
            .sr(N__19530));
    defparam \b2v_inst36.count_9_LC_2_4_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_9_LC_2_4_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_9_LC_2_4_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst36.count_9_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(N__16755),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37027),
            .ce(N__16943),
            .sr(N__19530));
    defparam \b2v_inst36.count_RNIFSRG1_12_LC_2_4_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIFSRG1_12_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIFSRG1_12_LC_2_4_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIFSRG1_12_LC_2_4_2  (
            .in0(N__16776),
            .in1(N__16935),
            .in2(_gnd_net_),
            .in3(N__16769),
            .lcout(\b2v_inst36.countZ0Z_12 ),
            .ltout(\b2v_inst36.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIR03I1_0_9_LC_2_4_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIR03I1_0_9_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIR03I1_0_9_LC_2_4_3 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst36.count_RNIR03I1_0_9_LC_2_4_3  (
            .in0(N__16938),
            .in1(N__16754),
            .in2(N__16740),
            .in3(N__16737),
            .lcout(\b2v_inst36.un12_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_13_LC_2_4_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_13_LC_2_4_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_13_LC_2_4_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_13_LC_2_4_4  (
            .in0(N__16665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37027),
            .ce(N__16943),
            .sr(N__19530));
    defparam \b2v_inst36.count_RNIJ2UG1_14_LC_2_4_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJ2UG1_14_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJ2UG1_14_LC_2_4_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNIJ2UG1_14_LC_2_4_5  (
            .in0(N__16937),
            .in1(N__17019),
            .in2(_gnd_net_),
            .in3(N__17030),
            .lcout(\b2v_inst36.countZ0Z_14 ),
            .ltout(\b2v_inst36.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_15_LC_2_4_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_15_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_15_LC_2_4_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst36.count_RNI_15_LC_2_4_6  (
            .in0(N__16656),
            .in1(N__16844),
            .in2(N__16710),
            .in3(N__16706),
            .lcout(\b2v_inst36.un12_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIHVSG1_13_LC_2_4_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIHVSG1_13_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIHVSG1_13_LC_2_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNIHVSG1_13_LC_2_4_7  (
            .in0(N__16936),
            .in1(N__16671),
            .in2(_gnd_net_),
            .in3(N__16664),
            .lcout(\b2v_inst36.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_15_LC_2_5_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_15_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_15_LC_2_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_15_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16865),
            .lcout(\b2v_inst36.count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36966),
            .ce(N__16942),
            .sr(N__19542));
    defparam \b2v_inst36.count_14_LC_2_5_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_14_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_14_LC_2_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_14_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17034),
            .lcout(\b2v_inst36.count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36966),
            .ce(N__16942),
            .sr(N__19542));
    defparam \b2v_inst36.curr_state_RNINSDS_0_LC_2_5_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNINSDS_0_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNINSDS_0_LC_2_5_2 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \b2v_inst36.curr_state_RNINSDS_0_LC_2_5_2  (
            .in0(N__23090),
            .in1(N__23036),
            .in2(N__23148),
            .in3(N__27562),
            .lcout(\b2v_inst36.curr_state_RNINSDSZ0Z_0 ),
            .ltout(\b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIL5VG1_15_LC_2_5_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIL5VG1_15_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIL5VG1_15_LC_2_5_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst36.count_RNIL5VG1_15_LC_2_5_3  (
            .in0(N__16866),
            .in1(_gnd_net_),
            .in2(N__16854),
            .in3(N__16851),
            .lcout(\b2v_inst36.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIPLHU_2_LC_2_5_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIPLHU_2_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIPLHU_2_LC_2_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIPLHU_2_LC_2_5_4  (
            .in0(N__19314),
            .in1(N__19325),
            .in2(_gnd_net_),
            .in3(N__19224),
            .lcout(\b2v_inst16.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_2_5_5 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_2_5_5 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \b2v_inst16.curr_state_RNIKEBL_1_LC_2_5_5  (
            .in0(N__27563),
            .in1(N__19798),
            .in2(_gnd_net_),
            .in3(N__20486),
            .lcout(\b2v_inst16.count_en ),
            .ltout(\b2v_inst16.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI12MU_6_LC_2_5_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI12MU_6_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI12MU_6_LC_2_5_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst16.count_RNI12MU_6_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(N__19287),
            .in2(N__16830),
            .in3(N__19305),
            .lcout(\b2v_inst16.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_2_6_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_2_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__16826),
            .in2(N__16815),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_6_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_6_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_6_1  (
            .in0(N__19781),
            .in1(N__16790),
            .in2(_gnd_net_),
            .in3(N__16779),
            .lcout(\b2v_inst16.count_rst_7 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_1 ),
            .carryout(\b2v_inst16.un4_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_6_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17269),
            .in3(N__17238),
            .lcout(\b2v_inst16.un4_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_2 ),
            .carryout(\b2v_inst16.un4_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_6_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__17235),
            .in2(_gnd_net_),
            .in3(N__17202),
            .lcout(\b2v_inst16.un4_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_3 ),
            .carryout(\b2v_inst16.un4_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_6_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__17199),
            .in2(_gnd_net_),
            .in3(N__17151),
            .lcout(\b2v_inst16.un4_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_4 ),
            .carryout(\b2v_inst16.un4_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_6_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_6_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_6_5  (
            .in0(N__19782),
            .in1(N__17147),
            .in2(_gnd_net_),
            .in3(N__17136),
            .lcout(\b2v_inst16.count_rst_11 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_5 ),
            .carryout(\b2v_inst16.un4_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_6_6 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__17132),
            .in2(_gnd_net_),
            .in3(N__17082),
            .lcout(\b2v_inst16.un4_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_6 ),
            .carryout(\b2v_inst16.un4_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_6_7 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17331),
            .in3(N__17079),
            .lcout(\b2v_inst16.un4_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_7 ),
            .carryout(\b2v_inst16.un4_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_7_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__17287),
            .in2(_gnd_net_),
            .in3(N__17076),
            .lcout(\b2v_inst16.un4_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_7_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_7_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_7_1  (
            .in0(N__19773),
            .in1(N__17408),
            .in2(_gnd_net_),
            .in3(N__17073),
            .lcout(\b2v_inst16.count_rst ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_9 ),
            .carryout(\b2v_inst16.un4_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_7_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__17070),
            .in2(_gnd_net_),
            .in3(N__17373),
            .lcout(\b2v_inst16.un4_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_10 ),
            .carryout(\b2v_inst16.un4_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_7_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_7_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_7_3  (
            .in0(N__19774),
            .in1(N__17357),
            .in2(_gnd_net_),
            .in3(N__17370),
            .lcout(\b2v_inst16.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_11 ),
            .carryout(\b2v_inst16.un4_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_2_7_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_2_7_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_2_7_4  (
            .in0(N__19797),
            .in1(N__18911),
            .in2(_gnd_net_),
            .in3(N__17367),
            .lcout(\b2v_inst16.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_12 ),
            .carryout(\b2v_inst16.un4_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_7_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_7_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_7_5  (
            .in0(N__19772),
            .in1(N__18866),
            .in2(_gnd_net_),
            .in3(N__17364),
            .lcout(\b2v_inst16.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_13 ),
            .carryout(\b2v_inst16.un4_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_7_6 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_7_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_7_6  (
            .in0(N__18956),
            .in1(N__19771),
            .in2(_gnd_net_),
            .in3(N__17361),
            .lcout(\b2v_inst16.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIR4KE_12_LC_2_7_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIR4KE_12_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIR4KE_12_LC_2_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIR4KE_12_LC_2_7_7  (
            .in0(N__17385),
            .in1(N__17397),
            .in2(_gnd_net_),
            .in3(N__19245),
            .lcout(\b2v_inst16.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_8_0 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_8_0 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_8_0  (
            .in0(N__19763),
            .in1(N__17345),
            .in2(N__17499),
            .in3(N__17326),
            .lcout(\b2v_inst16.count_rst_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_2_8_1 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_2_8_1 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_2_8_1  (
            .in0(N__17511),
            .in1(N__19762),
            .in2(N__17294),
            .in3(N__17498),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI7BPU_9_LC_2_8_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI7BPU_9_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI7BPU_9_LC_2_8_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNI7BPU_9_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__17433),
            .in2(N__17298),
            .in3(N__19247),
            .lcout(\b2v_inst16.countZ0Z_9 ),
            .ltout(\b2v_inst16.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_9_LC_2_8_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_9_LC_2_8_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_9_LC_2_8_3 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.count_9_LC_2_8_3  (
            .in0(N__17510),
            .in1(N__19765),
            .in2(N__17502),
            .in3(N__17494),
            .lcout(\b2v_inst16.count_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37095),
            .ce(N__19276),
            .sr(N__19123));
    defparam \b2v_inst16.curr_state_RNI_0_LC_2_8_4 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI_0_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI_0_LC_2_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst16.curr_state_RNI_0_LC_2_8_4  (
            .in0(N__19764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.N_3037_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_10_LC_2_8_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_10_LC_2_8_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_10_LC_2_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_10_LC_2_8_5  (
            .in0(N__17420),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37095),
            .ce(N__19276),
            .sr(N__19123));
    defparam \b2v_inst16.count_RNIG7TP_10_LC_2_8_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIG7TP_10_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIG7TP_10_LC_2_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIG7TP_10_LC_2_8_6  (
            .in0(N__17427),
            .in1(N__17421),
            .in2(_gnd_net_),
            .in3(N__19246),
            .lcout(\b2v_inst16.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_12_LC_2_8_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_12_LC_2_8_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_12_LC_2_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_12_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17396),
            .lcout(\b2v_inst16.count_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37095),
            .ce(N__19276),
            .sr(N__19123));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_0_LC_2_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_0_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_0_LC_2_9_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_0_LC_2_9_0  (
            .in0(N__17859),
            .in1(N__17885),
            .in2(_gnd_net_),
            .in3(N__17556),
            .lcout(),
            .ltout(\b2v_inst11.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNI82MVJ62_0_LC_2_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNI82MVJ62_0_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNI82MVJ62_0_LC_2_9_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.curr_state_RNI82MVJ62_0_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__17550),
            .in2(N__17379),
            .in3(N__28390),
            .lcout(\b2v_inst11.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst11.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_2_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_2_9_2 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_LC_2_9_2  (
            .in0(N__28391),
            .in1(_gnd_net_),
            .in2(N__17376),
            .in3(N__17884),
            .lcout(\b2v_inst11.count_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNO_0_LC_2_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_2_9_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \b2v_inst11.pwm_out_RNO_0_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__17855),
            .in2(N__17886),
            .in3(N__28392),
            .lcout(\b2v_inst11.g0_0_0_rep1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_LC_2_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_LC_2_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_LC_2_9_4  (
            .in0(N__19595),
            .in1(N__19624),
            .in2(_gnd_net_),
            .in3(N__19949),
            .lcout(\b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJZ0Z62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_0_LC_2_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_0_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.curr_state_0_LC_2_9_5 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \b2v_inst11.curr_state_0_LC_2_9_5  (
            .in0(N__17860),
            .in1(N__17826),
            .in2(N__19626),
            .in3(N__19594),
            .lcout(\b2v_inst11.curr_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37062),
            .ce(N__27541),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_2_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_2_9_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_0_LC_2_9_6  (
            .in0(N__28393),
            .in1(_gnd_net_),
            .in2(N__17864),
            .in3(N__17880),
            .lcout(\b2v_inst11.g0_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIKEBL_0_LC_2_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIKEBL_0_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIKEBL_0_LC_2_9_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst11.curr_state_RNIKEBL_0_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__27567),
            .in2(_gnd_net_),
            .in3(N__17854),
            .lcout(\b2v_inst11.g0_i_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_0_LC_2_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_0_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_0_LC_2_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_0_LC_2_10_0  (
            .in0(N__20086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20013),
            .lcout(\b2v_inst11.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37140),
            .ce(N__27538),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI03G9_0_LC_2_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI03G9_0_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI03G9_0_LC_2_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI03G9_0_LC_2_10_1  (
            .in0(N__17544),
            .in1(N__28351),
            .in2(_gnd_net_),
            .in3(N__19980),
            .lcout(\b2v_inst11.countZ0Z_0 ),
            .ltout(\b2v_inst11.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_1_LC_2_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_1_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_1_LC_2_10_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \b2v_inst11.count_RNI_1_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__17662),
            .in2(N__17538),
            .in3(N__20012),
            .lcout(),
            .ltout(\b2v_inst11.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI14G9_1_LC_2_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI14G9_1_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI14G9_1_LC_2_10_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \b2v_inst11.count_RNI14G9_1_LC_2_10_3  (
            .in0(N__28394),
            .in1(N__17637),
            .in2(N__17535),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_10_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_10_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(CONSTANT_ONE_NET_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_0_cry_0_c_inv_LC_2_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_0_c_inv_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_0_cry_0_c_inv_LC_2_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_0_cry_0_c_inv_LC_2_10_5  (
            .in0(N__17525),
            .in1(_gnd_net_),
            .in2(N__17532),
            .in3(N__20085),
            .lcout(\b2v_inst11.N_5852_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_1_LC_2_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_1_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_1_LC_2_10_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst11.count_1_LC_2_10_6  (
            .in0(N__20087),
            .in1(N__17661),
            .in2(_gnd_net_),
            .in3(N__20014),
            .lcout(\b2v_inst11.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37140),
            .ce(N__27538),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI0AHN_8_LC_2_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_2_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI0AHN_8_LC_2_10_7  (
            .in0(N__17631),
            .in1(N__28352),
            .in2(_gnd_net_),
            .in3(N__17621),
            .lcout(\b2v_inst11.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI2DIN_9_LC_2_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_2_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI2DIN_9_LC_2_11_0  (
            .in0(N__17598),
            .in1(N__28399),
            .in2(_gnd_net_),
            .in3(N__17606),
            .lcout(\b2v_inst11.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_9_LC_2_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_9_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_9_LC_2_11_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_9_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17610),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37135),
            .ce(N__27535),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIB49T_10_LC_2_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIB49T_10_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIB49T_10_LC_2_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIB49T_10_LC_2_11_2  (
            .in0(N__17580),
            .in1(N__28400),
            .in2(_gnd_net_),
            .in3(N__17588),
            .lcout(\b2v_inst11.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_10_LC_2_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_10_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_10_LC_2_11_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_10_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17592),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37135),
            .ce(N__27535),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIK61M_11_LC_2_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIK61M_11_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIK61M_11_LC_2_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIK61M_11_LC_2_11_4  (
            .in0(N__17562),
            .in1(N__28401),
            .in2(_gnd_net_),
            .in3(N__17570),
            .lcout(\b2v_inst11.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_11_LC_2_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_11_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_11_LC_2_11_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_11_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17574),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37135),
            .ce(N__27535),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIKNAN_2_LC_2_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_2_11_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNIKNAN_2_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__17742),
            .in2(N__17754),
            .in3(N__28398),
            .lcout(\b2v_inst11.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_2_LC_2_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_2_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_2_LC_2_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_2_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17753),
            .lcout(\b2v_inst11.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37135),
            .ce(N__27535),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIM92M_12_LC_2_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIM92M_12_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIM92M_12_LC_2_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIM92M_12_LC_2_12_0  (
            .in0(N__28404),
            .in1(N__17724),
            .in2(_gnd_net_),
            .in3(N__17732),
            .lcout(\b2v_inst11.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_12_LC_2_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_12_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_12_LC_2_12_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_12_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17736),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37134),
            .ce(N__27534),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIMQBN_3_LC_2_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_2_12_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \b2v_inst11.count_RNIMQBN_3_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__28402),
            .in2(N__17709),
            .in3(N__17717),
            .lcout(\b2v_inst11.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_3_LC_2_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_3_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_3_LC_2_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_3_LC_2_12_3  (
            .in0(N__17718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37134),
            .ce(N__27534),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOC3M_13_LC_2_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_2_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOC3M_13_LC_2_12_4  (
            .in0(N__28405),
            .in1(N__17688),
            .in2(_gnd_net_),
            .in3(N__17696),
            .lcout(\b2v_inst11.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_13_LC_2_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_13_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_13_LC_2_12_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_13_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17700),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37134),
            .ce(N__27534),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOTCN_4_LC_2_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_2_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOTCN_4_LC_2_12_6  (
            .in0(N__28403),
            .in1(N__17673),
            .in2(_gnd_net_),
            .in3(N__17681),
            .lcout(\b2v_inst11.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_4_LC_2_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_4_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_4_LC_2_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_4_LC_2_12_7  (
            .in0(N__17682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37134),
            .ce(N__27534),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_2_LC_2_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_2_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_2_LC_2_13_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.count_RNI_2_LC_2_13_0  (
            .in0(N__18270),
            .in1(N__18244),
            .in2(_gnd_net_),
            .in3(N__18220),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_5_LC_2_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_5_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_5_LC_2_13_1 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \b2v_inst11.count_RNI_5_LC_2_13_1  (
            .in0(N__18198),
            .in1(N__18161),
            .in2(N__18141),
            .in3(N__18137),
            .lcout(\b2v_inst11.un79_clk_100khzlto15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_10_LC_2_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_10_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_10_LC_2_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_RNI_10_LC_2_13_2  (
            .in0(N__18110),
            .in1(N__18076),
            .in2(N__18054),
            .in3(N__18024),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_15_LC_2_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_15_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_15_LC_2_13_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst11.count_RNI_15_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__17998),
            .in2(N__17976),
            .in3(N__17971),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_8_LC_2_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_8_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_8_LC_2_13_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.count_RNI_8_LC_2_13_4  (
            .in0(N__17952),
            .in1(N__17945),
            .in2(N__17919),
            .in3(N__17915),
            .lcout(\b2v_inst11.count_RNIZ0Z_8 ),
            .ltout(\b2v_inst11.count_RNIZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNO_0_0_LC_2_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNO_0_0_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNO_0_0_LC_2_13_5 .LUT_INIT=16'b0000001111001111;
    LogicCell40 \b2v_inst11.curr_state_RNO_0_0_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__17865),
            .in2(N__17829),
            .in3(N__19950),
            .lcout(\b2v_inst11.curr_state_3_i_m2_0_rep1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_1_c_inv_LC_2_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_1_c_inv_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_1_c_inv_LC_2_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_1_c_inv_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__17817),
            .in2(N__17805),
            .in3(N__23886),
            .lcout(\b2v_inst11.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_2_c_inv_LC_2_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_2_c_inv_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_2_c_inv_LC_2_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_2_c_inv_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__17787),
            .in2(N__17774),
            .in3(N__24027),
            .lcout(\b2v_inst11.un85_clk_100khz_0_0 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_1 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_3_c_inv_LC_2_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_3_c_inv_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_3_c_inv_LC_2_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_3_c_inv_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__18486),
            .in2(N__18474),
            .in3(N__23766),
            .lcout(\b2v_inst11.un85_clk_100khz_0_1 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_2 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_4_c_inv_LC_2_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_4_c_inv_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_4_c_inv_LC_2_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_4_c_inv_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__18455),
            .in2(N__18441),
            .in3(N__20196),
            .lcout(\b2v_inst11.un85_clk_100khz_0_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_3 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_5_c_inv_LC_2_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_5_c_inv_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_5_c_inv_LC_2_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_5_c_inv_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__18426),
            .in2(N__18413),
            .in3(N__20616),
            .lcout(\b2v_inst11.un85_clk_100khz_0_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_4 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_6_c_inv_LC_2_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_6_c_inv_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_6_c_inv_LC_2_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_6_c_inv_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__18393),
            .in2(N__18381),
            .in3(N__20580),
            .lcout(\b2v_inst11.un85_clk_100khz_0_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_5 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_7_c_inv_LC_2_14_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_7_c_inv_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_7_c_inv_LC_2_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_7_c_inv_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__18347),
            .in2(N__18363),
            .in3(N__20424),
            .lcout(\b2v_inst11.un85_clk_100khz_0_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_6 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_8_c_inv_LC_2_14_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_8_c_inv_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_8_c_inv_LC_2_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_8_c_inv_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__18333),
            .in2(N__18321),
            .in3(N__21762),
            .lcout(\b2v_inst11.un85_clk_100khz_0_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_7 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_9_c_inv_LC_2_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_9_c_inv_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_9_c_inv_LC_2_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_9_c_inv_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__18303),
            .in2(N__18290),
            .in3(N__21868),
            .lcout(\b2v_inst11.un85_clk_100khz_0_7 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_10_c_inv_LC_2_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_10_c_inv_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_10_c_inv_LC_2_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_10_c_inv_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__18681),
            .in2(N__18668),
            .in3(N__22101),
            .lcout(\b2v_inst11.un85_clk_100khz_1_8 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_9 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_11_c_inv_LC_2_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_11_c_inv_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_11_c_inv_LC_2_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_11_c_inv_LC_2_15_2  (
            .in0(N__22068),
            .in1(N__18629),
            .in2(N__18648),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_1_9 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_10 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_12_c_inv_LC_2_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_12_c_inv_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_12_c_inv_LC_2_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_12_c_inv_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__18599),
            .in2(N__18615),
            .in3(N__24102),
            .lcout(\b2v_inst11.un85_clk_100khz_1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_11 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_13_c_inv_LC_2_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_13_c_inv_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_13_c_inv_LC_2_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_13_c_inv_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__18566),
            .in2(N__18585),
            .in3(N__24198),
            .lcout(\b2v_inst11.un85_clk_100khz_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_12 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_14_c_inv_LC_2_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_14_c_inv_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_14_c_inv_LC_2_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_14_c_inv_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__18551),
            .in2(N__18537),
            .in3(N__25362),
            .lcout(\b2v_inst11.un85_clk_100khz_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_13 ),
            .carryout(\b2v_inst11.un85_clk_100khz_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_inv_LC_2_15_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_inv_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_inv_LC_2_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_15_c_inv_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(N__18522),
            .in3(N__25326),
            .lcout(\b2v_inst11.un85_clk_100khz_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_1_cry_14 ),
            .carryout(\b2v_inst11.un85_clk_100khz1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz1_THRU_LUT4_0_LC_2_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz1_THRU_LUT4_0_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz1_THRU_LUT4_0_LC_2_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz1_THRU_LUT4_0_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18492),
            .lcout(\b2v_inst11.un85_clk_100khz1_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__27069),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__23964),
            .in2(N__18698),
            .in3(N__18489),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__18694),
            .in2(N__21972),
            .in3(N__18714),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__22093),
            .in2(N__21945),
            .in3(N__18711),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__21921),
            .in2(N__22100),
            .in3(N__18708),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_16_5  (
            .in0(N__21867),
            .in1(N__22146),
            .in2(N__18699),
            .in3(N__18705),
            .lcout(\b2v_inst11.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22128),
            .in3(N__18702),
            .lcout(\b2v_inst11.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22092),
            .lcout(\b2v_inst11.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9S71_16_LC_4_1_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_4_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIB9S71_16_LC_4_1_0  (
            .in0(N__18743),
            .in1(N__20974),
            .in2(_gnd_net_),
            .in3(N__22612),
            .lcout(\b2v_inst200.un2_count_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_16_LC_4_1_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_16_LC_4_1_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_16_LC_4_1_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_16_LC_4_1_1  (
            .in0(N__20976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36800),
            .ce(N__22541),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNID13N_0_1_LC_4_1_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNID13N_0_1_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNID13N_0_1_LC_4_1_2 .LUT_INIT=16'b0000000001000111;
    LogicCell40 \b2v_inst200.count_RNID13N_0_1_LC_4_1_2  (
            .in0(N__18756),
            .in1(N__22614),
            .in2(N__18729),
            .in3(N__20754),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIOAVU1_1_LC_4_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIOAVU1_1_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIOAVU1_1_LC_4_1_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst200.count_RNIOAVU1_1_LC_4_1_3  (
            .in0(N__20847),
            .in1(N__18735),
            .in2(N__18762),
            .in3(N__22283),
            .lcout(\b2v_inst200.un25_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNID13N_1_LC_4_1_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNID13N_1_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNID13N_1_LC_4_1_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNID13N_1_LC_4_1_4  (
            .in0(N__18725),
            .in1(N__18755),
            .in2(_gnd_net_),
            .in3(N__22611),
            .lcout(\b2v_inst200.un2_count_1_axb_1 ),
            .ltout(\b2v_inst200.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_1_LC_4_1_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_1_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_1_LC_4_1_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst200.count_RNI_1_LC_4_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18759),
            .in3(N__22282),
            .lcout(\b2v_inst200.count_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9S71_0_16_LC_4_1_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9S71_0_16_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9S71_0_16_LC_4_1_6 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \b2v_inst200.count_RNIB9S71_0_16_LC_4_1_6  (
            .in0(N__18744),
            .in1(N__20975),
            .in2(N__20954),
            .in3(N__22613),
            .lcout(\b2v_inst200.un25_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_1_LC_4_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_1_LC_4_1_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_1_LC_4_1_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst200.count_1_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(N__20768),
            .in2(_gnd_net_),
            .in3(N__22284),
            .lcout(\b2v_inst200.count_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36800),
            .ce(N__22541),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3T051_3_LC_4_2_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3T051_3_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3T051_3_LC_4_2_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI3T051_3_LC_4_2_0  (
            .in0(N__18818),
            .in1(N__20725),
            .in2(_gnd_net_),
            .in3(N__22617),
            .lcout(\b2v_inst200.un2_count_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_3_LC_4_2_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_3_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_3_LC_4_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_3_LC_4_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20727),
            .lcout(\b2v_inst200.count_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36755),
            .ce(N__22539),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73351_0_5_LC_4_2_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73351_0_5_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73351_0_5_LC_4_2_2 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \b2v_inst200.count_RNI73351_0_5_LC_4_2_2  (
            .in0(N__20889),
            .in1(N__22621),
            .in2(N__18972),
            .in3(N__20685),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIUF4N4_3_LC_4_2_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIUF4N4_3_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIUF4N4_3_LC_4_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNIUF4N4_3_LC_4_2_3  (
            .in0(N__18810),
            .in1(N__18768),
            .in2(N__18717),
            .in3(N__18792),
            .lcout(\b2v_inst200.un25_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3T051_0_3_LC_4_2_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3T051_0_3_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3T051_0_3_LC_4_2_4 .LUT_INIT=16'b0000000001000111;
    LogicCell40 \b2v_inst200.count_RNI3T051_0_3_LC_4_2_4  (
            .in0(N__20726),
            .in1(N__22619),
            .in2(N__18822),
            .in3(N__20709),
            .lcout(\b2v_inst200.un25_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_13_LC_4_2_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_13_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_13_LC_4_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_13_LC_4_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20805),
            .lcout(\b2v_inst200.count_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36755),
            .ce(N__22539),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50P71_13_LC_4_2_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50P71_13_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50P71_13_LC_4_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI50P71_13_LC_4_2_6  (
            .in0(N__20803),
            .in1(N__18800),
            .in2(_gnd_net_),
            .in3(N__22618),
            .lcout(\b2v_inst200.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50P71_0_13_LC_4_2_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50P71_0_13_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50P71_0_13_LC_4_2_7 .LUT_INIT=16'b0000000000100111;
    LogicCell40 \b2v_inst200.count_RNI50P71_0_13_LC_4_2_7  (
            .in0(N__22620),
            .in1(N__20804),
            .in2(N__18804),
            .in3(N__20789),
            .lcout(\b2v_inst200.un25_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_12_LC_4_3_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_12_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_12_LC_4_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_12_LC_4_3_0  (
            .in0(N__20823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36719),
            .ce(N__22538),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_9_LC_4_3_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_9_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_9_LC_4_3_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_9_LC_4_3_1  (
            .in0(N__20865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36719),
            .ce(N__22538),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIFF751_9_LC_4_3_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIFF751_9_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIFF751_9_LC_4_3_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNIFF751_9_LC_4_3_2  (
            .in0(N__22623),
            .in1(N__18779),
            .in2(_gnd_net_),
            .in3(N__20863),
            .lcout(\b2v_inst200.un2_count_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3TN71_12_LC_4_3_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_4_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI3TN71_12_LC_4_3_3  (
            .in0(N__18786),
            .in1(N__20822),
            .in2(_gnd_net_),
            .in3(N__22625),
            .lcout(\b2v_inst200.countZ0Z_12 ),
            .ltout(\b2v_inst200.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIFF751_0_9_LC_4_3_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIFF751_0_9_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIFF751_0_9_LC_4_3_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst200.count_RNIFF751_0_9_LC_4_3_4  (
            .in0(N__22626),
            .in1(N__18780),
            .in2(N__18771),
            .in3(N__20864),
            .lcout(\b2v_inst200.un25_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73351_5_LC_4_3_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73351_5_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73351_5_LC_4_3_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI73351_5_LC_4_3_5  (
            .in0(N__18968),
            .in1(N__22622),
            .in2(_gnd_net_),
            .in3(N__20683),
            .lcout(\b2v_inst200.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_5_LC_4_3_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_5_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_5_LC_4_3_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_5_LC_4_3_6  (
            .in0(N__20684),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36719),
            .ce(N__22538),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QM71_11_LC_4_3_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_4_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI1QM71_11_LC_4_3_7  (
            .in0(N__22239),
            .in1(N__22250),
            .in2(_gnd_net_),
            .in3(N__22624),
            .lcout(\b2v_inst200.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI1ENE_15_LC_4_4_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI1ENE_15_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI1ENE_15_LC_4_4_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNI1ENE_15_LC_4_4_0  (
            .in0(N__19278),
            .in1(N__18921),
            .in2(_gnd_net_),
            .in3(N__18935),
            .lcout(\b2v_inst16.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_15_LC_4_4_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_15_LC_4_4_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_15_LC_4_4_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_15_LC_4_4_1  (
            .in0(N__18936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36872),
            .ce(N__19277),
            .sr(N__19146));
    defparam \b2v_inst16.count_RNIT7LE_13_LC_4_4_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIT7LE_13_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIT7LE_13_LC_4_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNIT7LE_13_LC_4_4_2  (
            .in0(N__18894),
            .in1(N__18876),
            .in2(_gnd_net_),
            .in3(N__19271),
            .lcout(\b2v_inst16.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_13_LC_4_4_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_13_LC_4_4_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_13_LC_4_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_13_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18893),
            .lcout(\b2v_inst16.count_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36872),
            .ce(N__19277),
            .sr(N__19146));
    defparam \b2v_inst16.count_RNIVAME_14_LC_4_4_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIVAME_14_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIVAME_14_LC_4_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNIVAME_14_LC_4_4_4  (
            .in0(N__18843),
            .in1(N__18828),
            .in2(_gnd_net_),
            .in3(N__19272),
            .lcout(\b2v_inst16.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_14_LC_4_4_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_14_LC_4_4_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_14_LC_4_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_14_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18842),
            .lcout(\b2v_inst16.count_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36872),
            .ce(N__19277),
            .sr(N__19146));
    defparam \b2v_inst200.count_RNI1QV41_2_LC_4_4_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_4_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI1QV41_2_LC_4_4_6  (
            .in0(N__22206),
            .in1(N__22191),
            .in2(_gnd_net_),
            .in3(N__22615),
            .lcout(\b2v_inst200.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50251_4_LC_4_4_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50251_4_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50251_4_LC_4_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI50251_4_LC_4_4_7  (
            .in0(N__22616),
            .in1(N__22164),
            .in2(_gnd_net_),
            .in3(N__22179),
            .lcout(\b2v_inst200.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_2_LC_4_5_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_2_LC_4_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_2_LC_4_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_2_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19332),
            .lcout(\b2v_inst16.count_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36965),
            .ce(N__19257),
            .sr(N__19145));
    defparam \b2v_inst16.count_6_LC_4_5_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_6_LC_4_5_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_6_LC_4_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_6_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19304),
            .lcout(\b2v_inst16.count_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36965),
            .ce(N__19257),
            .sr(N__19145));
    defparam \b2v_inst36.curr_state_0_LC_4_6_0 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_0_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_0_LC_4_6_0 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \b2v_inst36.curr_state_0_LC_4_6_0  (
            .in0(N__23150),
            .in1(N__23021),
            .in2(N__19082),
            .in3(N__23072),
            .lcout(\b2v_inst36.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36873),
            .ce(N__27543),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_1_LC_4_6_1 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_1_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_1_LC_4_6_1 .LUT_INIT=16'b0001010100010000;
    LogicCell40 \b2v_inst36.curr_state_1_LC_4_6_1  (
            .in0(N__23020),
            .in1(N__19073),
            .in2(N__23082),
            .in3(N__23151),
            .lcout(\b2v_inst36.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36873),
            .ce(N__27543),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_4_6_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_4_6_2 .LUT_INIT=16'b0000001000110010;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m6_LC_4_6_2  (
            .in0(N__23153),
            .in1(N__23016),
            .in2(N__23086),
            .in3(N__19072),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIU72Q_1_LC_4_6_3 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIU72Q_1_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIU72Q_1_LC_4_6_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.curr_state_RNIU72Q_1_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__19095),
            .in2(N__19089),
            .in3(N__28330),
            .lcout(\b2v_inst36.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_4_6_4 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_4_6_4 .LUT_INIT=16'b0011100000001000;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m4_LC_4_6_4  (
            .in0(N__23152),
            .in1(N__23022),
            .in2(N__19086),
            .in3(N__19071),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIT62Q_0_LC_4_6_5 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIT62Q_0_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIT62Q_0_LC_4_6_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.curr_state_RNIT62Q_0_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__18981),
            .in2(N__18975),
            .in3(N__28329),
            .lcout(\b2v_inst36.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIRQCA_0_LC_4_6_6 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIRQCA_0_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIRQCA_0_LC_4_6_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \b2v_inst36.curr_state_RNIRQCA_0_LC_4_6_6  (
            .in0(N__23154),
            .in1(N__28343),
            .in2(N__19563),
            .in3(N__23067),
            .lcout(\b2v_inst36.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_LC_4_6_7 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.DSW_PWROK_LC_4_6_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \b2v_inst36.DSW_PWROK_LC_4_6_7  (
            .in0(N__23068),
            .in1(_gnd_net_),
            .in2(N__23029),
            .in3(N__23149),
            .lcout(\b2v_inst36.DSW_PWROK_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36873),
            .ce(N__27543),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI5MK6V3_11_LC_4_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI5MK6V3_11_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI5MK6V3_11_LC_4_7_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNI5MK6V3_11_LC_4_7_0  (
            .in0(N__19350),
            .in1(N__28545),
            .in2(N__26556),
            .in3(N__21125),
            .lcout(\b2v_inst11.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_11_LC_4_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_11_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_11_LC_4_7_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_11_LC_4_7_1  (
            .in0(N__21126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26552),
            .lcout(\b2v_inst11.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37071),
            .ce(N__28532),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_10_LC_4_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_10_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_10_LC_4_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_10_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__26547),
            .in2(_gnd_net_),
            .in3(N__21141),
            .lcout(\b2v_inst11.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37071),
            .ce(N__28532),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIS7D3V3_10_LC_4_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIS7D3V3_10_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIS7D3V3_10_LC_4_7_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_off_RNIS7D3V3_10_LC_4_7_3  (
            .in0(N__28544),
            .in1(N__19344),
            .in2(N__26554),
            .in3(N__21140),
            .lcout(\b2v_inst11.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI7PL6V3_12_LC_4_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI7PL6V3_12_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI7PL6V3_12_LC_4_7_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_off_RNI7PL6V3_12_LC_4_7_5  (
            .in0(N__28546),
            .in1(N__19338),
            .in2(N__26555),
            .in3(N__21110),
            .lcout(\b2v_inst11.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_12_LC_4_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_12_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_12_LC_4_7_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.count_off_12_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21114),
            .in3(N__26548),
            .lcout(\b2v_inst11.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37071),
            .ce(N__28532),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIJMQ2V3_9_LC_4_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIJMQ2V3_9_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIJMQ2V3_9_LC_4_7_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_off_RNIJMQ2V3_9_LC_4_7_7  (
            .in0(N__28543),
            .in1(N__24795),
            .in2(N__26553),
            .in3(N__24806),
            .lcout(\b2v_inst11.count_offZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI74K2V3_3_LC_4_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI74K2V3_3_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI74K2V3_3_LC_4_8_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNI74K2V3_3_LC_4_8_0  (
            .in0(N__19659),
            .in1(N__28533),
            .in2(N__21012),
            .in3(N__26523),
            .lcout(\b2v_inst11.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_3_LC_4_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_3_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_3_LC_4_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_3_LC_4_8_1  (
            .in0(N__26527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21011),
            .lcout(\b2v_inst11.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37007),
            .ce(N__28547),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_13_LC_4_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_13_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_13_LC_4_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_13_LC_4_8_2  (
            .in0(N__21084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26528),
            .lcout(\b2v_inst11.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37007),
            .ce(N__28547),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNID2P6V3_15_LC_4_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNID2P6V3_15_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNID2P6V3_15_LC_4_8_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.count_off_RNID2P6V3_15_LC_4_8_3  (
            .in0(N__26526),
            .in1(N__22938),
            .in2(N__28551),
            .in3(N__22949),
            .lcout(\b2v_inst11.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_14_LC_4_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_14_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_14_LC_4_8_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_14_LC_4_8_4  (
            .in0(N__21264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26529),
            .lcout(\b2v_inst11.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37007),
            .ce(N__28547),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIBVN6V3_14_LC_4_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIBVN6V3_14_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIBVN6V3_14_LC_4_8_5 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.count_off_RNIBVN6V3_14_LC_4_8_5  (
            .in0(N__26525),
            .in1(N__19653),
            .in2(N__28550),
            .in3(N__21263),
            .lcout(\b2v_inst11.count_offZ0Z_14 ),
            .ltout(\b2v_inst11.count_offZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_15_LC_4_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_15_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_15_LC_4_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_15_LC_4_8_6  (
            .in0(N__21098),
            .in1(N__22905),
            .in2(N__19644),
            .in3(N__21251),
            .lcout(\b2v_inst11.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI9SM6V3_13_LC_4_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI9SM6V3_13_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI9SM6V3_13_LC_4_8_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.count_off_RNI9SM6V3_13_LC_4_8_7  (
            .in0(N__26524),
            .in1(N__19641),
            .in2(N__28549),
            .in3(N__21083),
            .lcout(\b2v_inst11.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNI9STGK62_LC_4_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNI9STGK62_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNI9STGK62_LC_4_9_0 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNI9STGK62_LC_4_9_0  (
            .in0(N__19635),
            .in1(N__19948),
            .in2(N__19625),
            .in3(N__19596),
            .lcout(\b2v_inst11.N_6 ),
            .ltout(\b2v_inst11.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_LC_4_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_LC_4_9_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.pwm_out_LC_4_9_1 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \b2v_inst11.pwm_out_LC_4_9_1  (
            .in0(N__19907),
            .in1(N__35808),
            .in2(N__19566),
            .in3(N__19895),
            .lcout(\b2v_inst11.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37001),
            .ce(),
            .sr(N__19920));
    defparam \b2v_inst11.pwm_out_RNINR3DL62_LC_4_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNINR3DL62_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNINR3DL62_LC_4_9_2 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \b2v_inst11.pwm_out_RNINR3DL62_LC_4_9_2  (
            .in0(N__27566),
            .in1(N__19908),
            .in2(N__19899),
            .in3(N__19884),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_en_LC_4_9_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_en_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_en_LC_4_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_en_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__27564),
            .in2(_gnd_net_),
            .in3(N__21054),
            .lcout(\b2v_inst200.count_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIV6I72_0_LC_4_9_4 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIV6I72_0_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIV6I72_0_LC_4_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst16.curr_state_RNIV6I72_0_LC_4_9_4  (
            .in0(N__27565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19815),
            .lcout(\b2v_inst16.delayed_vddq_pwrgd_en ),
            .ltout(\b2v_inst16.delayed_vddq_pwrgd_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNIPAU73_LC_4_9_5 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNIPAU73_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNIPAU73_LC_4_9_5 .LUT_INIT=16'b1010110011111111;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_RNIPAU73_LC_4_9_5  (
            .in0(N__20485),
            .in1(N__20442),
            .in2(N__19851),
            .in3(N__26784),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIBO6I1_0_0_LC_4_9_6 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIBO6I1_0_0_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIBO6I1_0_0_LC_4_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst16.curr_state_RNIBO6I1_0_0_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__19830),
            .in2(_gnd_net_),
            .in3(N__20484),
            .lcout(\b2v_inst16.N_268 ),
            .ltout(\b2v_inst16.N_268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI35HL1_0_LC_4_9_7 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI35HL1_0_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI35HL1_0_LC_4_9_7 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \b2v_inst16.curr_state_RNI35HL1_0_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19809),
            .in3(N__28389),
            .lcout(\b2v_inst16.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_4_10_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_4_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_2_c_RNO_LC_4_10_0  (
            .in0(N__21452),
            .in1(N__21467),
            .in2(N__21438),
            .in3(N__21482),
            .lcout(\b2v_inst20.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_4_10_3 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_4_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_5_c_RNO_LC_4_10_3  (
            .in0(N__21548),
            .in1(N__21533),
            .in2(N__21519),
            .in3(N__21500),
            .lcout(\b2v_inst20.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_0_LC_4_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_0_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_0_LC_4_10_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_RNI_0_LC_4_10_5  (
            .in0(N__20091),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\b2v_inst11.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__31582),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__23850),
            .in2(N__19970),
            .in3(N__23877),
            .lcout(G_2848),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__19966),
            .in2(N__23586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__23878),
            .in2(N__23571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__23556),
            .in2(N__23885),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__23544),
            .in2(N__19971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_s_6_LC_4_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_s_6_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_s_6_LC_4_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_s_6_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(N__23532),
            .in2(_gnd_net_),
            .in3(N__19953),
            .lcout(\b2v_inst11.mult1_un166_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27255),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__21708),
            .in2(N__20120),
            .in3(N__20139),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__20116),
            .in2(N__20103),
            .in3(N__20136),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__20184),
            .in2(N__20241),
            .in3(N__20133),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__20229),
            .in2(N__20192),
            .in3(N__20130),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_12_5  (
            .in0(N__23749),
            .in1(N__20220),
            .in2(N__20121),
            .in3(N__20127),
            .lcout(\b2v_inst11.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20211),
            .in3(N__20124),
            .lcout(\b2v_inst11.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20183),
            .lcout(\b2v_inst11.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__27222),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__25092),
            .in2(N__20162),
            .in3(N__20094),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__20158),
            .in2(N__20340),
            .in3(N__20232),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__20608),
            .in2(N__20316),
            .in3(N__20223),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__20292),
            .in2(N__20615),
            .in3(N__20214),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_13_5  (
            .in0(N__20188),
            .in1(N__20658),
            .in2(N__20163),
            .in3(N__20202),
            .lcout(\b2v_inst11.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__20640),
            .in2(_gnd_net_),
            .in3(N__20199),
            .lcout(\b2v_inst11.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20607),
            .lcout(\b2v_inst11.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__27110),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__21690),
            .in2(N__21731),
            .in3(N__20145),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__21727),
            .in2(N__21678),
            .in3(N__20142),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__21651),
            .in2(N__21761),
            .in3(N__20280),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__21757),
            .in2(N__21897),
            .in3(N__20277),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_14_5  (
            .in0(N__20415),
            .in1(N__21831),
            .in2(N__21732),
            .in3(N__20274),
            .lcout(\b2v_inst11.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21792),
            .in3(N__20271),
            .lcout(\b2v_inst11.mult1_un117_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20268),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__27146),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__20346),
            .in2(N__20378),
            .in3(N__20265),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__20374),
            .in2(N__20262),
            .in3(N__20253),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__20250),
            .in2(N__20423),
            .in3(N__20244),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__20419),
            .in2(N__20397),
            .in3(N__20388),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_15_5  (
            .in0(N__20572),
            .in1(N__20385),
            .in2(N__20379),
            .in3(N__20361),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20358),
            .in3(N__20349),
            .lcout(\b2v_inst11.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_15_7  (
            .in0(N__27114),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__27186),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__21702),
            .in2(N__20546),
            .in3(N__20328),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__20542),
            .in2(N__20325),
            .in3(N__20304),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__20568),
            .in2(N__20301),
            .in3(N__20283),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__20664),
            .in2(N__20576),
            .in3(N__20649),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_16_5  (
            .in0(N__20603),
            .in1(N__20646),
            .in2(N__20547),
            .in3(N__20631),
            .lcout(\b2v_inst11.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20628),
            .in3(N__20619),
            .lcout(\b2v_inst11.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20567),
            .lcout(\b2v_inst11.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_5_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_5_1_0 .LUT_INIT=16'b1111011111000100;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_LC_5_1_0  (
            .in0(N__20529),
            .in1(N__20508),
            .in2(N__20496),
            .in3(N__20435),
            .lcout(\b2v_inst16.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36640),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73Q71_14_LC_5_1_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_5_1_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst200.count_RNI73Q71_14_LC_5_1_1  (
            .in0(N__22609),
            .in1(N__22227),
            .in2(_gnd_net_),
            .in3(N__22212),
            .lcout(\b2v_inst200.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI96451_6_LC_5_1_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI96451_6_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI96451_6_LC_5_1_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI96451_6_LC_5_1_2  (
            .in0(N__22685),
            .in1(N__22674),
            .in2(_gnd_net_),
            .in3(N__22606),
            .lcout(\b2v_inst200.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9551_7_LC_5_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9551_7_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9551_7_LC_5_1_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNIB9551_7_LC_5_1_3  (
            .in0(N__22607),
            .in1(N__22656),
            .in2(_gnd_net_),
            .in3(N__22667),
            .lcout(\b2v_inst200.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDCT71_17_LC_5_1_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_5_1_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIDCT71_17_LC_5_1_4  (
            .in0(N__20919),
            .in1(N__20934),
            .in2(_gnd_net_),
            .in3(N__22610),
            .lcout(\b2v_inst200.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_0_LC_5_1_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_0_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_0_LC_5_1_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst200.count_RNI_0_LC_5_1_5  (
            .in0(N__22287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22314),
            .lcout(),
            .ltout(\b2v_inst200.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_0_LC_5_1_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_0_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_0_LC_5_1_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.count_RNIC03N_0_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(N__22257),
            .in2(N__20772),
            .in3(N__22605),
            .lcout(\b2v_inst200.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_5_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_5_1_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst200.count_RNIOMPC1_10_LC_5_1_7  (
            .in0(N__22608),
            .in1(_gnd_net_),
            .in2(N__22635),
            .in3(N__22650),
            .lcout(\b2v_inst200.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_1_c_LC_5_2_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_1_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_1_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_1_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__22285),
            .in2(N__20769),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_2_1 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__20753),
            .in2(_gnd_net_),
            .in3(N__20736),
            .lcout(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_1 ),
            .carryout(\b2v_inst200.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_2_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__20733),
            .in2(_gnd_net_),
            .in3(N__20712),
            .lcout(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_2 ),
            .carryout(\b2v_inst200.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_2_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__20708),
            .in2(_gnd_net_),
            .in3(N__20694),
            .lcout(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_3 ),
            .carryout(\b2v_inst200.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_2_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__20691),
            .in2(_gnd_net_),
            .in3(N__20670),
            .lcout(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_4 ),
            .carryout(\b2v_inst200.un2_count_1_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_2_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_2_5  (
            .in0(N__22339),
            .in1(N__22457),
            .in2(_gnd_net_),
            .in3(N__20667),
            .lcout(\b2v_inst200.count_1_6 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_5_cZ0 ),
            .carryout(\b2v_inst200.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_2_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__20888),
            .in2(_gnd_net_),
            .in3(N__20877),
            .lcout(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_6 ),
            .carryout(\b2v_inst200.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_7  (
            .in0(N__22340),
            .in1(N__22008),
            .in2(_gnd_net_),
            .in3(N__20874),
            .lcout(\b2v_inst200.count_1_8 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_7 ),
            .carryout(\b2v_inst200.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_3_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__20871),
            .in2(_gnd_net_),
            .in3(N__20853),
            .lcout(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_3_1 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_3_1  (
            .in0(N__22341),
            .in1(N__22403),
            .in2(_gnd_net_),
            .in3(N__20850),
            .lcout(\b2v_inst200.count_1_10 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_9 ),
            .carryout(\b2v_inst200.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_3_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_3_2  (
            .in0(N__22355),
            .in1(N__20843),
            .in2(_gnd_net_),
            .in3(N__20832),
            .lcout(\b2v_inst200.count_1_11 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_10 ),
            .carryout(\b2v_inst200.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_3_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__20829),
            .in2(_gnd_net_),
            .in3(N__20814),
            .lcout(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_11 ),
            .carryout(\b2v_inst200.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_3_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(N__20811),
            .in2(_gnd_net_),
            .in3(N__20793),
            .lcout(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_12 ),
            .carryout(\b2v_inst200.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_3_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__20790),
            .in2(_gnd_net_),
            .in3(N__20775),
            .lcout(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_13 ),
            .carryout(\b2v_inst200.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_5_3_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_5_3_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22020),
            .in3(N__20988),
            .lcout(\b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_14 ),
            .carryout(\b2v_inst200.un2_count_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_7  (
            .in0(N__22342),
            .in1(N__20985),
            .in2(_gnd_net_),
            .in3(N__20958),
            .lcout(\b2v_inst200.count_1_16 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_15 ),
            .carryout(\b2v_inst200.un2_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_4_0 .C_ON=1'b0;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_4_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_4_0  (
            .in0(N__20955),
            .in1(N__22344),
            .in2(_gnd_net_),
            .in3(N__20937),
            .lcout(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_17_LC_5_4_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_17_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_17_LC_5_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_17_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20933),
            .lcout(\b2v_inst200.count_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36810),
            .ce(N__22542),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_5_4_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_5_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__21049),
            .in2(_gnd_net_),
            .in3(N__22343),
            .lcout(\b2v_inst200.N_282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI_1_LC_5_5_0 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI_1_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI_1_LC_5_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst200.curr_state_RNI_1_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21328),
            .lcout(\b2v_inst200.N_2989_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_5_1 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_5_1 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_5_1  (
            .in0(N__21307),
            .in1(N__21350),
            .in2(N__21335),
            .in3(N__27762),
            .lcout(),
            .ltout(\b2v_inst200.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI26MQ4_1_LC_5_5_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI26MQ4_1_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI26MQ4_1_LC_5_5_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst200.curr_state_RNI26MQ4_1_LC_5_5_2  (
            .in0(N__28320),
            .in1(_gnd_net_),
            .in2(N__20910),
            .in3(N__21294),
            .lcout(\b2v_inst200.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_5_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_5_3 .LUT_INIT=16'b0001000010110101;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_5_3  (
            .in0(N__21308),
            .in1(N__20907),
            .in2(N__20892),
            .in3(N__27761),
            .lcout(\b2v_inst200.m6_i_0 ),
            .ltout(\b2v_inst200.m6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_5_4 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_5_4 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_5_4  (
            .in0(N__21050),
            .in1(_gnd_net_),
            .in2(N__21063),
            .in3(N__22354),
            .lcout(),
            .ltout(\b2v_inst200.N_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI19645_0_LC_5_5_5 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI19645_0_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI19645_0_LC_5_5_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.curr_state_RNI19645_0_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__21021),
            .in2(N__21060),
            .in3(N__28319),
            .lcout(\b2v_inst200.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_5_6 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_5_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21057),
            .in3(N__21176),
            .lcout(N_411),
            .ltout(N_411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_0_LC_5_5_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_0_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_0_LC_5_5_7 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \b2v_inst200.curr_state_0_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__22356),
            .in2(N__21030),
            .in3(N__21027),
            .lcout(\b2v_inst200.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36823),
            .ce(N__27544),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_5_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_5_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__22856),
            .in2(N__22901),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_5_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_5_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22842),
            .in3(N__21015),
            .lcout(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_1 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_5_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_5_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23201),
            .in3(N__20997),
            .lcout(\b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_2 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_5_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_5_6_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22992),
            .in3(N__20994),
            .lcout(\b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_3 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_5_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_5_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23361),
            .in3(N__20991),
            .lcout(\b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_4 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_5_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_5_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_5_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23310),
            .in3(N__21153),
            .lcout(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_5 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_5_6_6 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_5_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24609),
            .in3(N__21150),
            .lcout(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_6 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_5_6_7 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_5_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__24525),
            .in2(_gnd_net_),
            .in3(N__21147),
            .lcout(\b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_7 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_5_7_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_5_7_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21198),
            .in3(N__21144),
            .lcout(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_5_7_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_5_7_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21212),
            .in3(N__21129),
            .lcout(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_9 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_5_7_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_5_7_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21225),
            .in3(N__21117),
            .lcout(\b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_10 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_5_7_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_5_7_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21237),
            .in3(N__21102),
            .lcout(\b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_11 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_5_7_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_5_7_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21099),
            .in3(N__21075),
            .lcout(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_12 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_5_7_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_5_7_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21072),
            .in3(N__21255),
            .lcout(\b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_13 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_5_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_5_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_5_7_6  (
            .in0(N__21252),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21240),
            .lcout(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_9_LC_5_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_9_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_9_LC_5_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_9_LC_5_7_7  (
            .in0(N__21236),
            .in1(N__21224),
            .in2(N__21213),
            .in3(N__21197),
            .lcout(\b2v_inst11.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI37MQ4_2_LC_5_8_0 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI37MQ4_2_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI37MQ4_2_LC_5_8_0 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \b2v_inst200.curr_state_RNI37MQ4_2_LC_5_8_0  (
            .in0(N__21159),
            .in1(N__21183),
            .in2(_gnd_net_),
            .in3(N__28257),
            .lcout(\b2v_inst200.curr_state_i_2 ),
            .ltout(\b2v_inst200.curr_state_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_8_1 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_8_1 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \b2v_inst200.HDA_SDO_ATP_LC_5_8_1  (
            .in0(N__21395),
            .in1(_gnd_net_),
            .in2(N__21186),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.HDA_SDO_ATP_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36996),
            .ce(N__27536),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_8_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_8_2 .LUT_INIT=16'b1110111110101010;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_8_2  (
            .in0(N__21358),
            .in1(N__21394),
            .in2(N__27782),
            .in3(N__21381),
            .lcout(\b2v_inst200.i4_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_8_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_8_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst200.curr_state_RNI_0_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__21314),
            .in2(_gnd_net_),
            .in3(N__21177),
            .lcout(\b2v_inst200.N_205 ),
            .ltout(\b2v_inst200.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_2_LC_5_8_4 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_2_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_2_LC_5_8_4 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \b2v_inst200.curr_state_2_LC_5_8_4  (
            .in0(N__21359),
            .in1(N__21379),
            .in2(N__21162),
            .in3(N__27778),
            .lcout(\b2v_inst200.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36996),
            .ce(N__27536),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_5_8_5 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_5_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_7_c_RNO_LC_5_8_5  (
            .in0(N__21573),
            .in1(N__21615),
            .in2(N__21597),
            .in3(N__21633),
            .lcout(\b2v_inst20.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_8_6 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_8_6 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_8_6  (
            .in0(N__28259),
            .in1(N__21405),
            .in2(N__21399),
            .in3(N__21380),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_1_LC_5_8_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_1_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_1_LC_5_8_7 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \b2v_inst200.curr_state_1_LC_5_8_7  (
            .in0(N__27777),
            .in1(N__21360),
            .in2(N__21339),
            .in3(N__21315),
            .lcout(\b2v_inst200.curr_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36996),
            .ce(N__27536),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_c_LC_5_9_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_5_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_c_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__25013),
            .in2(N__23178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\b2v_inst20.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_5_9_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_5_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__24969),
            .in2(_gnd_net_),
            .in3(N__21282),
            .lcout(\b2v_inst20.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_1 ),
            .carryout(\b2v_inst20.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_5_9_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_5_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__24939),
            .in2(_gnd_net_),
            .in3(N__21279),
            .lcout(\b2v_inst20.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_2 ),
            .carryout(\b2v_inst20.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_5_9_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_5_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__24909),
            .in2(_gnd_net_),
            .in3(N__21276),
            .lcout(\b2v_inst20.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_3 ),
            .carryout(\b2v_inst20.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_5_9_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_5_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23256),
            .in3(N__21273),
            .lcout(\b2v_inst20.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_4 ),
            .carryout(\b2v_inst20.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_5_9_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_5_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__23226),
            .in2(_gnd_net_),
            .in3(N__21270),
            .lcout(\b2v_inst20.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_5 ),
            .carryout(\b2v_inst20.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_7_LC_5_9_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_7_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_7_LC_5_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_7_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__22826),
            .in2(_gnd_net_),
            .in3(N__21267),
            .lcout(\b2v_inst20.counterZ0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_6 ),
            .carryout(\b2v_inst20.counter_1_cry_7 ),
            .clk(N__37072),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_8_LC_5_9_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_8_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_8_LC_5_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_8_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__21483),
            .in2(_gnd_net_),
            .in3(N__21471),
            .lcout(\b2v_inst20.counterZ0Z_8 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_7 ),
            .carryout(\b2v_inst20.counter_1_cry_8 ),
            .clk(N__37072),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_9_LC_5_10_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_9_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_9_LC_5_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_9_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__21468),
            .in2(_gnd_net_),
            .in3(N__21456),
            .lcout(\b2v_inst20.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\b2v_inst20.counter_1_cry_9 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_10_LC_5_10_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_10_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_10_LC_5_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_10_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__21453),
            .in2(_gnd_net_),
            .in3(N__21441),
            .lcout(\b2v_inst20.counterZ0Z_10 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_9 ),
            .carryout(\b2v_inst20.counter_1_cry_10 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_11_LC_5_10_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_11_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_11_LC_5_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_11_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__21437),
            .in2(_gnd_net_),
            .in3(N__21423),
            .lcout(\b2v_inst20.counterZ0Z_11 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_10 ),
            .carryout(\b2v_inst20.counter_1_cry_11 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_12_LC_5_10_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_12_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_12_LC_5_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_12_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__23400),
            .in2(_gnd_net_),
            .in3(N__21420),
            .lcout(\b2v_inst20.counterZ0Z_12 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_11 ),
            .carryout(\b2v_inst20.counter_1_cry_12 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_13_LC_5_10_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_13_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_13_LC_5_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_13_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__23427),
            .in2(_gnd_net_),
            .in3(N__21417),
            .lcout(\b2v_inst20.counterZ0Z_13 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_12 ),
            .carryout(\b2v_inst20.counter_1_cry_13 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_14_LC_5_10_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_14_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_14_LC_5_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_14_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__23414),
            .in2(_gnd_net_),
            .in3(N__21414),
            .lcout(\b2v_inst20.counterZ0Z_14 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_13 ),
            .carryout(\b2v_inst20.counter_1_cry_14 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_15_LC_5_10_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_15_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_15_LC_5_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_15_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__23439),
            .in2(_gnd_net_),
            .in3(N__21411),
            .lcout(\b2v_inst20.counterZ0Z_15 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_14 ),
            .carryout(\b2v_inst20.counter_1_cry_15 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_16_LC_5_10_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_16_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_16_LC_5_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_16_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__23496),
            .in2(_gnd_net_),
            .in3(N__21408),
            .lcout(\b2v_inst20.counterZ0Z_16 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_15 ),
            .carryout(\b2v_inst20.counter_1_cry_16 ),
            .clk(N__36997),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_17_LC_5_11_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_17_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_17_LC_5_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_17_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__23484),
            .in2(_gnd_net_),
            .in3(N__21558),
            .lcout(\b2v_inst20.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\b2v_inst20.counter_1_cry_17 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_18_LC_5_11_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_18_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_18_LC_5_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_18_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__23471),
            .in2(_gnd_net_),
            .in3(N__21555),
            .lcout(\b2v_inst20.counterZ0Z_18 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_17 ),
            .carryout(\b2v_inst20.counter_1_cry_18 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_19_LC_5_11_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_19_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_19_LC_5_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_19_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__23457),
            .in2(_gnd_net_),
            .in3(N__21552),
            .lcout(\b2v_inst20.counterZ0Z_19 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_18 ),
            .carryout(\b2v_inst20.counter_1_cry_19 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_20_LC_5_11_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_20_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_20_LC_5_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_20_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__21549),
            .in2(_gnd_net_),
            .in3(N__21537),
            .lcout(\b2v_inst20.counterZ0Z_20 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_19 ),
            .carryout(\b2v_inst20.counter_1_cry_20 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_21_LC_5_11_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_21_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_21_LC_5_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_21_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__21534),
            .in2(_gnd_net_),
            .in3(N__21522),
            .lcout(\b2v_inst20.counterZ0Z_21 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_20 ),
            .carryout(\b2v_inst20.counter_1_cry_21 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_22_LC_5_11_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_22_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_22_LC_5_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_22_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__21518),
            .in2(_gnd_net_),
            .in3(N__21504),
            .lcout(\b2v_inst20.counterZ0Z_22 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_21 ),
            .carryout(\b2v_inst20.counter_1_cry_22 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_23_LC_5_11_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_23_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_23_LC_5_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_23_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__21501),
            .in2(_gnd_net_),
            .in3(N__21489),
            .lcout(\b2v_inst20.counterZ0Z_23 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_22 ),
            .carryout(\b2v_inst20.counter_1_cry_23 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_24_LC_5_11_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_24_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_24_LC_5_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_24_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__23652),
            .in2(_gnd_net_),
            .in3(N__21486),
            .lcout(\b2v_inst20.counterZ0Z_24 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_23 ),
            .carryout(\b2v_inst20.counter_1_cry_24 ),
            .clk(N__37002),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_25_LC_5_12_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_25_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_25_LC_5_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_25_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__23621),
            .in2(_gnd_net_),
            .in3(N__21642),
            .lcout(\b2v_inst20.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\b2v_inst20.counter_1_cry_25 ),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_26_LC_5_12_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_26_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_26_LC_5_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_26_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__23639),
            .in2(_gnd_net_),
            .in3(N__21639),
            .lcout(\b2v_inst20.counterZ0Z_26 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_25 ),
            .carryout(\b2v_inst20.counter_1_cry_26 ),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_27_LC_5_12_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_27_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_27_LC_5_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_27_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__23606),
            .in2(_gnd_net_),
            .in3(N__21636),
            .lcout(\b2v_inst20.counterZ0Z_27 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_26 ),
            .carryout(\b2v_inst20.counter_1_cry_27 ),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_28_LC_5_12_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_28_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_28_LC_5_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_28_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__21632),
            .in2(_gnd_net_),
            .in3(N__21618),
            .lcout(\b2v_inst20.counterZ0Z_28 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_27 ),
            .carryout(\b2v_inst20.counter_1_cry_28 ),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_29_LC_5_12_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_29_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_29_LC_5_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_29_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__21614),
            .in2(_gnd_net_),
            .in3(N__21600),
            .lcout(\b2v_inst20.counterZ0Z_29 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_28 ),
            .carryout(\b2v_inst20.counter_1_cry_29 ),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_30_LC_5_12_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_30_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_30_LC_5_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_30_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__21593),
            .in2(_gnd_net_),
            .in3(N__21579),
            .lcout(\b2v_inst20.counterZ0Z_30 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_29 ),
            .carryout(\b2v_inst20.counter_1_cry_30 ),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_31_LC_5_12_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_31_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_31_LC_5_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.counter_31_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__21572),
            .in2(_gnd_net_),
            .in3(N__21576),
            .lcout(\b2v_inst20.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37143),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_4_l_fx_LC_5_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_4_l_fx_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_4_l_fx_LC_5_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_4_l_fx_LC_5_12_7  (
            .in0(N__23819),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23748),
            .lcout(\b2v_inst11.mult1_un152_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23746),
            .lcout(\b2v_inst11.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27221),
            .lcout(\b2v_inst11.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_7_l_fx_LC_5_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_7_l_fx_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_7_l_fx_LC_5_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_7_l_fx_LC_5_13_2  (
            .in0(N__23699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23747),
            .lcout(\b2v_inst11.mult1_un152_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31987),
            .lcout(\b2v_inst11.N_2943_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27147),
            .lcout(\b2v_inst11.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21875),
            .lcout(\b2v_inst11.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27090),
            .lcout(\b2v_inst11.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27068),
            .lcout(\b2v_inst11.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__27086),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__21684),
            .in2(N__21809),
            .in3(N__21669),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__21805),
            .in2(N__21666),
            .in3(N__21645),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__21909),
            .in2(N__21885),
            .in3(N__21888),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__21884),
            .in2(N__21846),
            .in3(N__21825),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_14_5  (
            .in0(N__21753),
            .in1(N__21822),
            .in2(N__21810),
            .in3(N__21783),
            .lcout(\b2v_inst11.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21780),
            .in3(N__21765),
            .lcout(\b2v_inst11.mult1_un110_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un110_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_5_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_5_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21735),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__23973),
            .in2(N__21989),
            .in3(N__21714),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__21985),
            .in2(N__23898),
            .in3(N__21711),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__24090),
            .in2(N__24147),
            .in3(N__22002),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__24135),
            .in2(N__24098),
            .in3(N__21999),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5  (
            .in0(N__22063),
            .in1(N__24126),
            .in2(N__21990),
            .in3(N__21996),
            .lcout(\b2v_inst11.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24117),
            .in3(N__21993),
            .lcout(\b2v_inst11.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24089),
            .lcout(\b2v_inst11.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__27038),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_16_0_),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(N__27375),
            .in2(N__22037),
            .in3(N__21957),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__22033),
            .in2(N__21954),
            .in3(N__21933),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__22059),
            .in2(N__21930),
            .in3(N__21912),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(N__22152),
            .in2(N__22067),
            .in3(N__22137),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_16_5  (
            .in0(N__22091),
            .in1(N__22134),
            .in2(N__22038),
            .in3(N__22116),
            .lcout(\b2v_inst11.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22113),
            .in3(N__22104),
            .lcout(\b2v_inst11.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22058),
            .lcout(\b2v_inst11.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI2KKU_15_LC_6_1_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI2KKU_15_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI2KKU_15_LC_6_1_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI2KKU_15_LC_6_1_0  (
            .in0(N__22603),
            .in1(N__22472),
            .in2(_gnd_net_),
            .in3(N__22444),
            .lcout(\b2v_inst200.un2_count_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_15_LC_6_1_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_15_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_15_LC_6_1_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_15_LC_6_1_1  (
            .in0(N__22446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(N__22537),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_8_LC_6_1_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_8_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_8_LC_6_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_8_LC_6_1_2  (
            .in0(N__22430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(N__22537),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDC651_8_LC_6_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDC651_8_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDC651_8_LC_6_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIDC651_8_LC_6_1_3  (
            .in0(N__22416),
            .in1(N__22429),
            .in2(_gnd_net_),
            .in3(N__22602),
            .lcout(\b2v_inst200.un2_count_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI2KKU_0_15_LC_6_1_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI2KKU_0_15_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI2KKU_0_15_LC_6_1_4 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \b2v_inst200.count_RNI2KKU_0_15_LC_6_1_4  (
            .in0(N__22604),
            .in1(N__22473),
            .in2(N__22464),
            .in3(N__22445),
            .lcout(\b2v_inst200.un25_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDC651_0_8_LC_6_1_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDC651_0_8_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDC651_0_8_LC_6_1_5 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \b2v_inst200.count_RNIDC651_0_8_LC_6_1_5  (
            .in0(N__22431),
            .in1(N__22415),
            .in2(N__22404),
            .in3(N__22601),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI5RUP8_8_LC_6_1_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI5RUP8_8_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI5RUP8_8_LC_6_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNI5RUP8_8_LC_6_1_6  (
            .in0(N__22386),
            .in1(N__22374),
            .in2(N__22368),
            .in3(N__22365),
            .lcout(\b2v_inst200.count_RNI5RUP8Z0Z_8 ),
            .ltout(\b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_0_LC_6_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_0_LC_6_1_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_0_LC_6_1_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst200.count_0_LC_6_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22290),
            .in3(N__22286),
            .lcout(\b2v_inst200.count_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36436),
            .ce(N__22537),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_11_LC_6_2_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_11_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_11_LC_6_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_11_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22251),
            .lcout(\b2v_inst200.count_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_14_LC_6_2_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_14_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_14_LC_6_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_14_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22226),
            .lcout(\b2v_inst200.count_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_2_LC_6_2_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_2_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_2_LC_6_2_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst200.count_2_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(N__22205),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_4_LC_6_2_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_4_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_4_LC_6_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_4_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22178),
            .lcout(\b2v_inst200.count_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_6_LC_6_2_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_6_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_6_LC_6_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_6_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22686),
            .lcout(\b2v_inst200.count_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_7_LC_6_2_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_7_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_7_LC_6_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_7_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22668),
            .lcout(\b2v_inst200.count_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_10_LC_6_2_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_10_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_10_LC_6_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_10_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22649),
            .lcout(\b2v_inst200.count_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36775),
            .ce(N__22540),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_0_c_LC_6_3_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_0_c_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_0_c_LC_6_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_0_c_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__24348),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNILCP9_LC_6_3_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNILCP9_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNILCP9_LC_6_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_0_c_RNILCP9_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__24275),
            .in2(_gnd_net_),
            .in3(N__22488),
            .lcout(\b2v_inst5.un2_count_1_cry_0_c_RNILCPZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_0 ),
            .carryout(\b2v_inst5.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNIMEQ9_LC_6_3_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNIMEQ9_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNIMEQ9_LC_6_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_1_c_RNIMEQ9_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__25656),
            .in2(_gnd_net_),
            .in3(N__22485),
            .lcout(\b2v_inst5.un2_count_1_cry_1_c_RNIMEQZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_1 ),
            .carryout(\b2v_inst5.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_6_3_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_6_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__24288),
            .in2(_gnd_net_),
            .in3(N__22482),
            .lcout(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_2 ),
            .carryout(\b2v_inst5.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_6_3_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_6_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_6_3_4  (
            .in0(_gnd_net_),
            .in1(N__22739),
            .in2(_gnd_net_),
            .in3(N__22479),
            .lcout(\b2v_inst5.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_3 ),
            .carryout(\b2v_inst5.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIPKT9_LC_6_3_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIPKT9_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIPKT9_LC_6_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_4_c_RNIPKT9_LC_6_3_5  (
            .in0(_gnd_net_),
            .in1(N__25595),
            .in2(_gnd_net_),
            .in3(N__22476),
            .lcout(\b2v_inst5.un2_count_1_cry_4_c_RNIPKTZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_4 ),
            .carryout(\b2v_inst5.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIQMU9_LC_6_3_6 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIQMU9_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIQMU9_LC_6_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_5_c_RNIQMU9_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__25571),
            .in2(_gnd_net_),
            .in3(N__22713),
            .lcout(\b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_5 ),
            .carryout(\b2v_inst5.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIROV9_LC_6_3_7 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIROV9_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIROV9_LC_6_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_6_c_RNIROV9_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(N__25449),
            .in2(_gnd_net_),
            .in3(N__22710),
            .lcout(\b2v_inst5.un2_count_1_cry_6_c_RNIROVZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_6 ),
            .carryout(\b2v_inst5.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_6_4_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_6_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22796),
            .in3(N__22707),
            .lcout(\b2v_inst5.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_6_4_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_6_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(N__26028),
            .in2(_gnd_net_),
            .in3(N__22704),
            .lcout(\b2v_inst5.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_8 ),
            .carryout(\b2v_inst5.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_6_4_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_6_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__25560),
            .in2(_gnd_net_),
            .in3(N__22701),
            .lcout(\b2v_inst5.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_9 ),
            .carryout(\b2v_inst5.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_6_4_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_6_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_6_4_3  (
            .in0(N__25882),
            .in1(N__25482),
            .in2(_gnd_net_),
            .in3(N__22698),
            .lcout(\b2v_inst5.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_10 ),
            .carryout(\b2v_inst5.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_6_4_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_6_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__24362),
            .in2(_gnd_net_),
            .in3(N__22695),
            .lcout(\b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_11 ),
            .carryout(\b2v_inst5.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_6_4_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_6_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26163),
            .in3(N__22692),
            .lcout(\b2v_inst5.un2_count_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_12 ),
            .carryout(\b2v_inst5.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_6_4_6 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_6_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_6_4_6  (
            .in0(_gnd_net_),
            .in1(N__24372),
            .in2(_gnd_net_),
            .in3(N__22689),
            .lcout(\b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_13 ),
            .carryout(\b2v_inst5.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_6_4_7 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_6_4_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_6_4_7  (
            .in0(N__24438),
            .in1(N__25883),
            .in2(_gnd_net_),
            .in3(N__22812),
            .lcout(\b2v_inst5.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIH08H3_4_LC_6_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIH08H3_4_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIH08H3_4_LC_6_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIH08H3_4_LC_6_5_0  (
            .in0(N__22719),
            .in1(N__26250),
            .in2(_gnd_net_),
            .in3(N__22758),
            .lcout(\b2v_inst5.countZ0Z_4 ),
            .ltout(\b2v_inst5.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIU15T1_0_8_LC_6_5_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIU15T1_0_8_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIU15T1_0_8_LC_6_5_1 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \b2v_inst5.count_RNIU15T1_0_8_LC_6_5_1  (
            .in0(N__26252),
            .in1(N__22767),
            .in2(N__22809),
            .in3(N__22806),
            .lcout(\b2v_inst5.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_6_5_2 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_6_5_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_6_5_2  (
            .in0(N__26104),
            .in1(N__22778),
            .in2(N__22797),
            .in3(N__25855),
            .lcout(\b2v_inst5.count_rst_6 ),
            .ltout(\b2v_inst5.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIU15T1_8_LC_6_5_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIU15T1_8_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIU15T1_8_LC_6_5_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.count_RNIU15T1_8_LC_6_5_3  (
            .in0(N__26251),
            .in1(_gnd_net_),
            .in2(N__22800),
            .in3(N__22766),
            .lcout(\b2v_inst5.un2_count_1_axb_8 ),
            .ltout(\b2v_inst5.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_8_LC_6_5_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_8_LC_6_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_8_LC_6_5_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.count_8_LC_6_5_4  (
            .in0(N__26108),
            .in1(N__22779),
            .in2(N__22770),
            .in3(N__25857),
            .lcout(\b2v_inst5.count_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36822),
            .ce(N__26294),
            .sr(N__25991));
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_6_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_6_5_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_6_5_5  (
            .in0(N__25854),
            .in1(N__22751),
            .in2(N__22740),
            .in3(N__26103),
            .lcout(\b2v_inst5.count_rst_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_4_LC_6_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_4_LC_6_5_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_4_LC_6_5_6 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst5.count_4_LC_6_5_6  (
            .in0(N__22752),
            .in1(N__22735),
            .in2(N__26109),
            .in3(N__25856),
            .lcout(\b2v_inst5.count_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36822),
            .ce(N__26294),
            .sr(N__25991));
    defparam \b2v_inst5.count_RNIL9B73_0_LC_6_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL9B73_0_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL9B73_0_LC_6_5_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst5.count_RNIL9B73_0_LC_6_5_7  (
            .in0(N__25853),
            .in1(N__24484),
            .in2(_gnd_net_),
            .in3(N__26102),
            .lcout(\b2v_inst5.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_1_LC_6_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_1_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_1_LC_6_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_1_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__22872),
            .in2(_gnd_net_),
            .in3(N__26473),
            .lcout(\b2v_inst11.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36639),
            .ce(N__28531),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_2_LC_6_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_2_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_2_LC_6_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_2_LC_6_6_1  (
            .in0(N__26471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22923),
            .lcout(\b2v_inst11.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36639),
            .ce(N__28531),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_0_LC_6_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_0_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_0_LC_6_6_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_off_0_LC_6_6_2  (
            .in0(N__22900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26472),
            .lcout(\b2v_inst11.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36639),
            .ce(N__28531),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI51J2V3_2_LC_6_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI51J2V3_2_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI51J2V3_2_LC_6_6_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNI51J2V3_2_LC_6_6_3  (
            .in0(N__22929),
            .in1(N__28502),
            .in2(N__26522),
            .in3(N__22922),
            .lcout(\b2v_inst11.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI5TD0V3_0_LC_6_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI5TD0V3_0_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI5TD0V3_0_LC_6_6_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst11.count_off_RNI5TD0V3_0_LC_6_6_4  (
            .in0(N__22899),
            .in1(N__28500),
            .in2(N__22914),
            .in3(N__26466),
            .lcout(\b2v_inst11.count_offZ0Z_0 ),
            .ltout(\b2v_inst11.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_1_LC_6_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_1_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_1_LC_6_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.count_off_RNI_1_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22875),
            .in3(N__22857),
            .lcout(\b2v_inst11.count_off_RNIZ0Z_1 ),
            .ltout(\b2v_inst11.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI6UD0V3_1_LC_6_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI6UD0V3_1_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI6UD0V3_1_LC_6_6_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNI6UD0V3_1_LC_6_6_6  (
            .in0(N__22866),
            .in1(N__28501),
            .in2(N__22860),
            .in3(N__26467),
            .lcout(\b2v_inst11.count_offZ0Z_1 ),
            .ltout(\b2v_inst11.count_offZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_0_1_LC_6_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_0_1_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_0_1_LC_6_6_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.count_off_RNI_0_1_LC_6_6_7  (
            .in0(N__23306),
            .in1(N__23360),
            .in2(N__22845),
            .in3(N__22841),
            .lcout(\b2v_inst11.un34_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_6_7_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_6_7_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_RNO_LC_6_7_0  (
            .in0(N__23167),
            .in1(N__23248),
            .in2(N__23225),
            .in3(N__22827),
            .lcout(\b2v_inst20.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_5_LC_6_7_1 .C_ON=1'b0;
    defparam \b2v_inst20.counter_5_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_5_LC_6_7_1 .LUT_INIT=16'b0000011000000110;
    LogicCell40 \b2v_inst20.counter_5_LC_6_7_1  (
            .in0(N__23249),
            .in1(N__23265),
            .in2(N__26697),
            .in3(_gnd_net_),
            .lcout(\b2v_inst20.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36955),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_6_LC_6_7_2 .C_ON=1'b0;
    defparam \b2v_inst20.counter_6_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_6_LC_6_7_2 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst20.counter_6_LC_6_7_2  (
            .in0(N__23221),
            .in1(N__26691),
            .in2(_gnd_net_),
            .in3(N__23235),
            .lcout(\b2v_inst20.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36955),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_3_LC_6_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_3_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_3_LC_6_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_3_LC_6_7_4  (
            .in0(N__24605),
            .in1(N__22988),
            .in2(N__23205),
            .in3(N__24521),
            .lcout(\b2v_inst11.un34_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_LC_6_7_5 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_LC_6_7_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst20.tmp_1_LC_6_7_5  (
            .in0(N__26693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28258),
            .lcout(SYNTHESIZED_WIRE_1keep_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36955),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_LC_6_7_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_1_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_1_LC_6_7_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_1_LC_6_7_6  (
            .in0(N__23168),
            .in1(N__25017),
            .in2(_gnd_net_),
            .in3(N__26692),
            .lcout(\b2v_inst20.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36955),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI3E27_0_LC_6_7_7 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI3E27_0_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI3E27_0_LC_6_7_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst36.curr_state_RNI3E27_0_LC_6_7_7  (
            .in0(N__23147),
            .in1(N__23091),
            .in2(_gnd_net_),
            .in3(N__23040),
            .lcout(\b2v_inst36.curr_state_RNI3E27Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI97L2V3_4_LC_6_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI97L2V3_4_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI97L2V3_4_LC_6_8_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNI97L2V3_4_LC_6_8_0  (
            .in0(N__22956),
            .in1(N__28526),
            .in2(N__22974),
            .in3(N__26531),
            .lcout(\b2v_inst11.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_4_LC_6_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_4_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_4_LC_6_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_4_LC_6_8_1  (
            .in0(N__26533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22970),
            .lcout(\b2v_inst11.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36891),
            .ce(N__28548),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_15_LC_6_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_15_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_15_LC_6_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_15_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__22950),
            .in2(_gnd_net_),
            .in3(N__26537),
            .lcout(\b2v_inst11.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36891),
            .ce(N__28548),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_5_LC_6_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_5_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_5_LC_6_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_5_LC_6_8_3  (
            .in0(N__26534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23372),
            .lcout(\b2v_inst11.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36891),
            .ce(N__28548),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIBAM2V3_5_LC_6_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIBAM2V3_5_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIBAM2V3_5_LC_6_8_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNIBAM2V3_5_LC_6_8_4  (
            .in0(N__23382),
            .in1(N__28527),
            .in2(N__23376),
            .in3(N__26532),
            .lcout(\b2v_inst11.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_6_LC_6_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_6_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_6_LC_6_8_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_6_LC_6_8_5  (
            .in0(N__26535),
            .in1(_gnd_net_),
            .in2(N__23333),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36891),
            .ce(N__28548),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIDDN2V3_6_LC_6_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIDDN2V3_6_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIDDN2V3_6_LC_6_8_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNIDDN2V3_6_LC_6_8_6  (
            .in0(N__23343),
            .in1(N__28525),
            .in2(N__23337),
            .in3(N__26530),
            .lcout(\b2v_inst11.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_7_LC_6_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_7_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_7_LC_6_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_7_LC_6_8_7  (
            .in0(N__26536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24632),
            .lcout(\b2v_inst11.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36891),
            .ce(N__28548),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_LC_6_9_0 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_0_c_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_LC_6_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__24984),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\b2v_inst20.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_LC_6_9_1 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_1_c_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_LC_6_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__23286),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_0 ),
            .carryout(\b2v_inst20.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_LC_6_9_2 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_2_c_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_LC_6_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_2_c_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__23277),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_1 ),
            .carryout(\b2v_inst20.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_LC_6_9_3 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_3_c_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_LC_6_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_3_c_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__23388),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_2 ),
            .carryout(\b2v_inst20.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_LC_6_9_4 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_4_c_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_LC_6_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_4_c_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__23445),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_3 ),
            .carryout(\b2v_inst20.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_LC_6_9_5 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_5_c_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_LC_6_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_5_c_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__23517),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_4 ),
            .carryout(\b2v_inst20.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_LC_6_9_6 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_6_c_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_LC_6_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_6_c_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__23592),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_5 ),
            .carryout(\b2v_inst20.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_LC_6_9_7 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_7_c_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_LC_6_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_7_c_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__23505),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_6 ),
            .carryout(b2v_inst20_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_6_10_0.C_ON=1'b0;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_6_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23499),
            .lcout(b2v_inst20_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_6_10_2 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_6_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_4_c_RNO_LC_6_10_2  (
            .in0(N__23495),
            .in1(N__23483),
            .in2(N__23472),
            .in3(N__23456),
            .lcout(\b2v_inst20.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.G_149_LC_6_10_3 .C_ON=1'b0;
    defparam \b2v_inst5.G_149_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.G_149_LC_6_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst5.G_149_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__34240),
            .in2(_gnd_net_),
            .in3(N__26654),
            .lcout(G_149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_6_10_5 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_6_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_3_c_RNO_LC_6_10_5  (
            .in0(N__23438),
            .in1(N__23426),
            .in2(N__23415),
            .in3(N__23399),
            .lcout(\b2v_inst20.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_rep1_LC_6_10_6 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_rep1_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_rep1_LC_6_10_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst20.tmp_1_rep1_LC_6_10_6  (
            .in0(N__34241),
            .in1(_gnd_net_),
            .in2(N__26672),
            .in3(_gnd_net_),
            .lcout(SYNTHESIZED_WIRE_1keep_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36909),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_6_10_7 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_6_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_6_c_RNO_LC_6_10_7  (
            .in0(N__23651),
            .in1(N__23640),
            .in2(N__23625),
            .in3(N__23607),
            .lcout(\b2v_inst20.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__31460),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__25026),
            .in2(N__23990),
            .in3(N__23574),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__23986),
            .in2(N__23832),
            .in3(N__23559),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__23796),
            .in2(N__24020),
            .in3(N__23547),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__24016),
            .in2(N__23778),
            .in3(N__23535),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_11_5  (
            .in0(N__23873),
            .in1(N__23709),
            .in2(N__23991),
            .in3(N__23523),
            .lcout(\b2v_inst11.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23676),
            .in3(N__23520),
            .lcout(\b2v_inst11.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_11_7  (
            .in0(N__31461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_6_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_6_12_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_2_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31302),
            .in3(N__26813),
            .lcout(\b2v_inst11.N_366 ),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(N__25101),
            .in2(N__23841),
            .in3(N__23823),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__23820),
            .in2(N__23805),
            .in3(N__23790),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(N__23787),
            .in2(N__23765),
            .in3(N__23769),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__23761),
            .in2(N__23721),
            .in3(N__23703),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_12_5  (
            .in0(N__24012),
            .in1(N__23700),
            .in2(N__23685),
            .in3(N__23667),
            .lcout(\b2v_inst11.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23664),
            .in3(N__24030),
            .lcout(\b2v_inst11.mult1_un152_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23994),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27315),
            .lcout(\b2v_inst11.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27339),
            .lcout(\b2v_inst11.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_6_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_6_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27360),
            .lcout(\b2v_inst11.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27039),
            .lcout(\b2v_inst11.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_0_LC_6_13_5 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_0_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_0_LC_6_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_0_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27786),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_6_LC_6_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_6_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_6_LC_6_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_6_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33879),
            .lcout(\b2v_inst11.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37063),
            .ce(N__33837),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__27359),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__23907),
            .in2(N__24068),
            .in3(N__23889),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__24064),
            .in2(N__24042),
            .in3(N__24138),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__24186),
            .in2(N__24243),
            .in3(N__24129),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__24231),
            .in2(N__24194),
            .in3(N__24120),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_14_5  (
            .in0(N__24094),
            .in1(N__24222),
            .in2(N__24069),
            .in3(N__24108),
            .lcout(\b2v_inst11.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24213),
            .in3(N__24105),
            .lcout(\b2v_inst11.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24185),
            .lcout(\b2v_inst11.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__27335),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__24051),
            .in2(N__24164),
            .in3(N__24033),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__24160),
            .in2(N__25176),
            .in3(N__24234),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__25347),
            .in2(N__25437),
            .in3(N__24225),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__25416),
            .in2(N__25355),
            .in3(N__24216),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5  (
            .in0(N__24190),
            .in1(N__25401),
            .in2(N__24165),
            .in3(N__24204),
            .lcout(\b2v_inst11.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25386),
            .in3(N__24201),
            .lcout(\b2v_inst11.mult1_un75_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25346),
            .lcout(\b2v_inst11.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_15_LC_7_1_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_15_LC_7_1_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_15_LC_7_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_15_LC_7_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24456),
            .lcout(\b2v_inst5.count_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36427),
            .ce(N__26310),
            .sr(N__25990));
    defparam \b2v_inst5.count_RNIL6AH3_6_LC_7_2_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL6AH3_6_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL6AH3_6_LC_7_2_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst5.count_RNIL6AH3_6_LC_7_2_0  (
            .in0(N__26266),
            .in1(N__24317),
            .in2(N__24306),
            .in3(N__25966),
            .lcout(\b2v_inst5.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_5_LC_7_2_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_5_LC_7_2_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_5_LC_7_2_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst5.count_5_LC_7_2_1  (
            .in0(N__24336),
            .in1(_gnd_net_),
            .in2(N__25989),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36774),
            .ce(N__26270),
            .sr(N__25988));
    defparam \b2v_inst5.count_RNIJ39H3_5_LC_7_2_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIJ39H3_5_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIJ39H3_5_LC_7_2_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst5.count_RNIJ39H3_5_LC_7_2_2  (
            .in0(N__26265),
            .in1(N__24335),
            .in2(N__24327),
            .in3(N__25965),
            .lcout(\b2v_inst5.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_6_LC_7_2_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_6_LC_7_2_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_6_LC_7_2_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst5.count_6_LC_7_2_3  (
            .in0(N__25970),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24318),
            .lcout(\b2v_inst5.count_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36774),
            .ce(N__26270),
            .sr(N__25988));
    defparam \b2v_inst5.count_RNIH6CN3_13_LC_7_2_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIH6CN3_13_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIH6CN3_13_LC_7_2_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst5.count_RNIH6CN3_13_LC_7_2_4  (
            .in0(N__26118),
            .in1(_gnd_net_),
            .in2(N__26278),
            .in3(N__24294),
            .lcout(\b2v_inst5.countZ0Z_13 ),
            .ltout(\b2v_inst5.countZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_13_LC_7_2_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_13_LC_7_2_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_13_LC_7_2_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_13_LC_7_2_5  (
            .in0(N__26136),
            .in1(N__25976),
            .in2(N__24297),
            .in3(N__26090),
            .lcout(\b2v_inst5.count_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36774),
            .ce(N__26270),
            .sr(N__25988));
    defparam \b2v_inst5.count_RNIFT6H3_3_LC_7_2_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIFT6H3_3_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIFT6H3_3_LC_7_2_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst5.count_RNIFT6H3_3_LC_7_2_6  (
            .in0(N__26264),
            .in1(N__25631),
            .in2(N__25614),
            .in3(N__25964),
            .lcout(\b2v_inst5.countZ0Z_3 ),
            .ltout(\b2v_inst5.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI_1_LC_7_2_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI_1_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI_1_LC_7_2_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst5.count_RNI_1_LC_7_2_7  (
            .in0(N__25655),
            .in1(N__24279),
            .in2(N__24282),
            .in3(N__26155),
            .lcout(\b2v_inst5.un12_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIBN4H3_1_LC_7_3_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIBN4H3_1_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIBN4H3_1_LC_7_3_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst5.count_RNIBN4H3_1_LC_7_3_0  (
            .in0(N__24263),
            .in1(N__26223),
            .in2(N__24252),
            .in3(N__25897),
            .lcout(\b2v_inst5.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_1_LC_7_3_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_1_LC_7_3_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_1_LC_7_3_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst5.count_1_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__25978),
            .in2(_gnd_net_),
            .in3(N__24264),
            .lcout(\b2v_inst5.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36512),
            .ce(N__26287),
            .sr(N__25977));
    defparam \b2v_inst5.count_12_LC_7_3_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_12_LC_7_3_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_12_LC_7_3_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst5.count_12_LC_7_3_2  (
            .in0(N__24405),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25902),
            .lcout(\b2v_inst5.count_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36512),
            .ce(N__26287),
            .sr(N__25977));
    defparam \b2v_inst5.count_RNIF3BN3_12_LC_7_3_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIF3BN3_12_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIF3BN3_12_LC_7_3_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \b2v_inst5.count_RNIF3BN3_12_LC_7_3_3  (
            .in0(N__25898),
            .in1(N__24404),
            .in2(N__24396),
            .in3(N__26256),
            .lcout(\b2v_inst5.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_14_LC_7_3_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_14_LC_7_3_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_14_LC_7_3_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst5.count_14_LC_7_3_4  (
            .in0(N__24381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25903),
            .lcout(\b2v_inst5.count_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36512),
            .ce(N__26287),
            .sr(N__25977));
    defparam \b2v_inst5.count_RNIJ9DN3_14_LC_7_3_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIJ9DN3_14_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIJ9DN3_14_LC_7_3_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \b2v_inst5.count_RNIJ9DN3_14_LC_7_3_5  (
            .in0(N__24387),
            .in1(N__24380),
            .in2(N__25958),
            .in3(N__26257),
            .lcout(\b2v_inst5.countZ0Z_14 ),
            .ltout(\b2v_inst5.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIMP4T1_0_0_LC_7_3_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIMP4T1_0_0_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIMP4T1_0_0_LC_7_3_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst5.count_RNIMP4T1_0_0_LC_7_3_6  (
            .in0(N__24434),
            .in1(N__24485),
            .in2(N__24366),
            .in3(N__24363),
            .lcout(\b2v_inst5.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_0_LC_7_3_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_0_LC_7_3_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_0_LC_7_3_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst5.count_0_LC_7_3_7  (
            .in0(N__24486),
            .in1(N__25979),
            .in2(_gnd_net_),
            .in3(N__26089),
            .lcout(\b2v_inst5.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36512),
            .ce(N__26287),
            .sr(N__25977));
    defparam \b2v_inst5.curr_state_1_LC_7_4_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_1_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_1_LC_7_4_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst5.curr_state_1_LC_7_4_0  (
            .in0(N__24420),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36744),
            .ce(N__27539),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIRH7S1_0_LC_7_4_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIRH7S1_0_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIRH7S1_0_LC_7_4_1 .LUT_INIT=16'b1000000010001000;
    LogicCell40 \b2v_inst5.curr_state_RNIRH7S1_0_LC_7_4_1  (
            .in0(N__24679),
            .in1(N__35827),
            .in2(N__27735),
            .in3(N__24666),
            .lcout(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0 ),
            .ltout(\b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_7_4_2 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_7_4_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_7_4_2  (
            .in0(_gnd_net_),
            .in1(N__24507),
            .in2(N__24351),
            .in3(N__24494),
            .lcout(\b2v_inst5.un2_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIKEUB2_1_LC_7_4_3 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIKEUB2_1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIKEUB2_1_LC_7_4_3 .LUT_INIT=16'b0000110011111100;
    LogicCell40 \b2v_inst5.curr_state_RNIKEUB2_1_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(N__24342),
            .in2(N__28325),
            .in3(N__24419),
            .lcout(\b2v_inst5.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst5.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI_1_LC_7_4_4 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI_1_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI_1_LC_7_4_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst5.curr_state_RNI_1_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24510),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.curr_state_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIMP4T1_0_LC_7_4_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIMP4T1_0_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIMP4T1_0_LC_7_4_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \b2v_inst5.count_RNIMP4T1_0_LC_7_4_5  (
            .in0(N__24506),
            .in1(_gnd_net_),
            .in2(N__24498),
            .in3(N__26221),
            .lcout(\b2v_inst5.count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_7_4_6 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_7_4_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(N__24471),
            .in2(_gnd_net_),
            .in3(N__26081),
            .lcout(N_413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNILCEN3_15_LC_7_4_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNILCEN3_15_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNILCEN3_15_LC_7_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNILCEN3_15_LC_7_4_7  (
            .in0(N__24465),
            .in1(N__26222),
            .in2(_gnd_net_),
            .in3(N__24449),
            .lcout(\b2v_inst5.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_7_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_7_5_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst5.curr_state_RNI65HI_0_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__24705),
            .in2(N__28324),
            .in3(N__24411),
            .lcout(\b2v_inst5.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst5.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_7_5_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_7_5_1 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m6_i_LC_7_5_1  (
            .in0(N__24664),
            .in1(N__27732),
            .in2(N__24423),
            .in3(N__24716),
            .lcout(\b2v_inst5.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_LC_7_5_2 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.RSMRSTn_LC_7_5_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst5.RSMRSTn_LC_7_5_2  (
            .in0(N__27731),
            .in1(_gnd_net_),
            .in2(N__24699),
            .in3(N__24663),
            .lcout(RSMRSTn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36611),
            .ce(N__27537),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_7_5_3 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_7_5_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_LC_7_5_3  (
            .in0(N__28790),
            .in1(N__24681),
            .in2(_gnd_net_),
            .in3(N__24715),
            .lcout(\b2v_inst5.m4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNID8DP1_0_LC_7_5_4 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNID8DP1_0_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNID8DP1_0_LC_7_5_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst5.curr_state_RNID8DP1_0_LC_7_5_4  (
            .in0(N__27733),
            .in1(_gnd_net_),
            .in2(N__24698),
            .in3(N__24662),
            .lcout(curr_state_RNID8DP1_0_0),
            .ltout(curr_state_RNID8DP1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_0_LC_7_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_0_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_0_LC_7_5_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \b2v_inst5.curr_state_0_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__24680),
            .in2(N__24720),
            .in3(N__24717),
            .lcout(\b2v_inst5.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36611),
            .ce(N__27537),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI65HI_0_0_LC_7_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI65HI_0_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI65HI_0_0_LC_7_5_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst5.curr_state_RNI65HI_0_0_LC_7_5_6  (
            .in0(N__24694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.N_2856_i ),
            .ltout(\b2v_inst5.N_2856_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIVF6A1_0_LC_7_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIVF6A1_0_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIVF6A1_0_LC_7_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.curr_state_RNIVF6A1_0_LC_7_5_7  (
            .in0(N__24665),
            .in1(N__27734),
            .in2(N__24645),
            .in3(N__28260),
            .lcout(\b2v_inst5.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIFGO2V3_7_LC_7_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIFGO2V3_7_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIFGO2V3_7_LC_7_6_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNIFGO2V3_7_LC_7_6_0  (
            .in0(N__24642),
            .in1(N__28499),
            .in2(N__24633),
            .in3(N__26457),
            .lcout(\b2v_inst11.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_8_LC_7_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_8_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_8_LC_7_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_8_LC_7_6_1  (
            .in0(N__26458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24545),
            .lcout(\b2v_inst11.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36745),
            .ce(N__28524),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_1_1_LC_7_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_1_1_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_1_1_LC_7_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_off_RNI_1_1_LC_7_6_2  (
            .in0(N__24591),
            .in1(N__24579),
            .in2(N__24573),
            .in3(N__24558),
            .lcout(\b2v_inst11.count_off_RNI_1Z0Z_1 ),
            .ltout(\b2v_inst11.count_off_RNI_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI794G3_1_LC_7_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI794G3_1_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI794G3_1_LC_7_6_3 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \b2v_inst11.func_state_RNI794G3_1_LC_7_6_3  (
            .in0(N__24822),
            .in1(N__32305),
            .in2(N__24552),
            .in3(N__28003),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNICMPB4_0_LC_7_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNICMPB4_0_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNICMPB4_0_LC_7_6_4 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \b2v_inst11.func_state_RNICMPB4_0_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__28718),
            .in2(N__24549),
            .in3(N__30761),
            .lcout(\b2v_inst11.func_state_RNICMPB4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIHJP2V3_8_LC_7_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIHJP2V3_8_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIHJP2V3_8_LC_7_6_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst11.count_off_RNIHJP2V3_8_LC_7_6_6  (
            .in0(N__24546),
            .in1(N__26460),
            .in2(N__24534),
            .in3(N__28498),
            .lcout(\b2v_inst11.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_9_LC_7_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_9_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_9_LC_7_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_9_LC_7_6_7  (
            .in0(N__26459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24813),
            .lcout(\b2v_inst11.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36745),
            .ce(N__28524),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI6IFF4_0_1_LC_7_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI6IFF4_0_1_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI6IFF4_0_1_LC_7_7_0 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \b2v_inst11.func_state_RNI6IFF4_0_1_LC_7_7_0  (
            .in0(N__26628),
            .in1(N__37346),
            .in2(N__28719),
            .in3(N__24768),
            .lcout(\b2v_inst11.func_state_RNI6IFF4_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI05F44_1_LC_7_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI05F44_1_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI05F44_1_LC_7_7_1 .LUT_INIT=16'b1100111111011111;
    LogicCell40 \b2v_inst11.func_state_RNI05F44_1_LC_7_7_1  (
            .in0(N__38982),
            .in1(N__26583),
            .in2(N__37357),
            .in3(N__33940),
            .lcout(\b2v_inst11.N_76 ),
            .ltout(\b2v_inst11.N_76_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNII89R8_0_LC_7_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNII89R8_0_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNII89R8_0_LC_7_7_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst11.func_state_RNII89R8_0_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__24759),
            .in2(N__24783),
            .in3(N__24780),
            .lcout(\b2v_inst11.func_state_1_m2_1 ),
            .ltout(\b2v_inst11.func_state_1_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNICD8EB_1_LC_7_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNICD8EB_1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNICD8EB_1_LC_7_7_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst11.func_state_RNICD8EB_1_LC_7_7_3  (
            .in0(N__24878),
            .in1(N__26773),
            .in2(N__24774),
            .in3(N__26732),
            .lcout(\b2v_inst11.func_state ),
            .ltout(\b2v_inst11.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNITPVU_1_LC_7_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNITPVU_1_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNITPVU_1_LC_7_7_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \b2v_inst11.func_state_RNITPVU_1_LC_7_7_4  (
            .in0(N__38562),
            .in1(N__38725),
            .in2(N__24771),
            .in3(N__28240),
            .lcout(\b2v_inst11.N_339 ),
            .ltout(\b2v_inst11.N_339_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI6IFF4_1_LC_7_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI6IFF4_1_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI6IFF4_1_LC_7_7_5 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \b2v_inst11.func_state_RNI6IFF4_1_LC_7_7_5  (
            .in0(N__37350),
            .in1(N__26627),
            .in2(N__24762),
            .in3(N__28714),
            .lcout(\b2v_inst11.func_state_RNI6IFF4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_RNIPUMD_LC_7_7_6 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_RNIPUMD_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.DSW_PWROK_RNIPUMD_LC_7_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst36.DSW_PWROK_RNIPUMD_LC_7_7_6  (
            .in0(N__24753),
            .in1(N__24741),
            .in2(_gnd_net_),
            .in3(N__28241),
            .lcout(dsw_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_LC_7_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_1_LC_7_7_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst11.func_state_1_LC_7_7_7  (
            .in0(N__24879),
            .in1(N__26774),
            .in2(N__24888),
            .in3(N__26733),
            .lcout(\b2v_inst11.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37018),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI3NQD_1_LC_7_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI3NQD_1_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI3NQD_1_LC_7_8_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI3NQD_1_LC_7_8_0  (
            .in0(N__28893),
            .in1(N__38983),
            .in2(N__38565),
            .in3(N__32266),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_51_and_i_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNILBJP_1_LC_7_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNILBJP_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNILBJP_1_LC_7_8_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \b2v_inst11.func_state_RNILBJP_1_LC_7_8_1  (
            .in0(N__34261),
            .in1(N__28800),
            .in2(N__24870),
            .in3(N__28107),
            .lcout(\b2v_inst11.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_7_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_7_8_2 .LUT_INIT=16'b0101011111011111;
    LogicCell40 \b2v_inst11.VCCST_EN_i_0_o3_0_LC_7_8_2  (
            .in0(N__38554),
            .in1(N__34259),
            .in2(N__28115),
            .in3(N__28795),
            .lcout(VCCST_EN_i_0_o3_0),
            .ltout(VCCST_EN_i_0_o3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un1_vddq_en_LC_7_8_3 .C_ON=1'b0;
    defparam \b2v_inst16.un1_vddq_en_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un1_vddq_en_LC_7_8_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst16.un1_vddq_en_LC_7_8_3  (
            .in0(N__24867),
            .in1(_gnd_net_),
            .in2(N__24849),
            .in3(_gnd_net_),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_en_0_x1_LC_7_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_en_0_x1_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_en_0_x1_LC_7_8_4 .LUT_INIT=16'b1000110011001100;
    LogicCell40 \b2v_inst11.count_clk_en_0_x1_LC_7_8_4  (
            .in0(N__38555),
            .in1(N__34258),
            .in2(N__38675),
            .in3(N__28794),
            .lcout(),
            .ltout(\b2v_inst11.count_clk_en_0_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_en_0_ns_LC_7_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_en_0_ns_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_en_0_ns_LC_7_8_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_en_0_ns_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24825),
            .in3(N__26673),
            .lcout(\b2v_inst11.count_clk_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_7_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_7_8_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_7_8_6  (
            .in0(N__38556),
            .in1(N__34260),
            .in2(N__38676),
            .in3(N__28796),
            .lcout(\b2v_inst11.N_185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVT4P1_1_LC_7_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVT4P1_1_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVT4P1_1_LC_7_8_7 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \b2v_inst11.func_state_RNIVT4P1_1_LC_7_8_7  (
            .in0(N__30767),
            .in1(N__37356),
            .in2(N__39060),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_7_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_7_9_0 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_7_9_0  (
            .in0(N__34265),
            .in1(N__28116),
            .in2(N__38674),
            .in3(N__28809),
            .lcout(v5s_enn),
            .ltout(v5s_enn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIKAJP_2_LC_7_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIKAJP_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIKAJP_2_LC_7_9_1 .LUT_INIT=16'b0000010100001110;
    LogicCell40 \b2v_inst11.dutycycle_RNIKAJP_2_LC_7_9_1  (
            .in0(N__39001),
            .in1(N__32304),
            .in2(N__25020),
            .in3(N__31295),
            .lcout(\b2v_inst11.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_0_LC_7_9_2 .C_ON=1'b0;
    defparam \b2v_inst20.counter_0_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_0_LC_7_9_2 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \b2v_inst20.counter_0_LC_7_9_2  (
            .in0(N__26669),
            .in1(_gnd_net_),
            .in2(N__25012),
            .in3(_gnd_net_),
            .lcout(\b2v_inst20.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37088),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_LC_7_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_LC_7_9_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_1_LC_7_9_3  (
            .in0(N__38528),
            .in1(N__38645),
            .in2(N__39085),
            .in3(N__34800),
            .lcout(\b2v_inst11.func_state_RNIDQ4A1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_7_9_4 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_7_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_RNO_LC_7_9_4  (
            .in0(N__25002),
            .in1(N__24961),
            .in2(N__24938),
            .in3(N__24904),
            .lcout(\b2v_inst20.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_2_LC_7_9_5 .C_ON=1'b0;
    defparam \b2v_inst20.counter_2_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_2_LC_7_9_5 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \b2v_inst20.counter_2_LC_7_9_5  (
            .in0(N__24978),
            .in1(_gnd_net_),
            .in2(N__24968),
            .in3(N__26670),
            .lcout(\b2v_inst20.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37088),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_3_LC_7_9_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_3_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_3_LC_7_9_6 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \b2v_inst20.counter_3_LC_7_9_6  (
            .in0(N__24934),
            .in1(_gnd_net_),
            .in2(N__26680),
            .in3(N__24948),
            .lcout(\b2v_inst20.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37088),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_4_LC_7_9_7 .C_ON=1'b0;
    defparam \b2v_inst20.counter_4_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_4_LC_7_9_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_4_LC_7_9_7  (
            .in0(N__24905),
            .in1(N__24918),
            .in2(_gnd_net_),
            .in3(N__26671),
            .lcout(\b2v_inst20.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37088),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI498D2_5_LC_7_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI498D2_5_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI498D2_5_LC_7_10_0 .LUT_INIT=16'b1111111100001101;
    LogicCell40 \b2v_inst11.dutycycle_RNI498D2_5_LC_7_10_0  (
            .in0(N__25041),
            .in1(N__39296),
            .in2(N__29087),
            .in3(N__29151),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIB79JE_3_LC_7_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIB79JE_3_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIB79JE_3_LC_7_10_1 .LUT_INIT=16'b0101111101011101;
    LogicCell40 \b2v_inst11.dutycycle_RNIB79JE_3_LC_7_10_1  (
            .in0(N__37345),
            .in1(N__30824),
            .in2(N__24891),
            .in3(N__25071),
            .lcout(\b2v_inst11.dutycycle_eena_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVK_LC_7_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVK_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVK_LC_7_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVK_LC_7_10_2  (
            .in0(N__31179),
            .in1(N__35946),
            .in2(_gnd_net_),
            .in3(N__30534),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVKZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIKJFD2_LC_7_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIKJFD2_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIKJFD2_LC_7_10_3 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIKJFD2_LC_7_10_3  (
            .in0(N__39057),
            .in1(N__38641),
            .in2(N__25044),
            .in3(N__25032),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_7_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_7_10_4 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_5_LC_7_10_4  (
            .in0(N__32303),
            .in1(N__39059),
            .in2(_gnd_net_),
            .in3(N__35947),
            .lcout(\b2v_inst11.N_236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI34G9_0_LC_7_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI34G9_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI34G9_0_LC_7_10_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.func_state_RNI34G9_0_LC_7_10_5  (
            .in0(N__39297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32301),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINGLA1_1_LC_7_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINGLA1_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINGLA1_1_LC_7_10_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNINGLA1_1_LC_7_10_6  (
            .in0(N__38404),
            .in1(N__34251),
            .in2(N__25035),
            .in3(N__39056),
            .lcout(\b2v_inst11.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_7_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_7_10_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_9_LC_7_10_7  (
            .in0(N__39058),
            .in1(N__38159),
            .in2(_gnd_net_),
            .in3(N__32302),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31296),
            .lcout(\b2v_inst11.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_14_0_LC_7_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_14_0_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_14_0_LC_7_11_1 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_14_0_LC_7_11_1  (
            .in0(N__26832),
            .in1(N__28860),
            .in2(N__34194),
            .in3(N__34036),
            .lcout(\b2v_inst11.dutycycle_RNI_14Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_13_0_LC_7_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_13_0_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_13_0_LC_7_11_2 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_13_0_LC_7_11_2  (
            .in0(N__28859),
            .in1(N__25050),
            .in2(N__34049),
            .in3(N__34189),
            .lcout(),
            .ltout(\b2v_inst11.N_3055_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIK9J85_5_LC_7_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIK9J85_5_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIK9J85_5_LC_7_11_3 .LUT_INIT=16'b1010111110101100;
    LogicCell40 \b2v_inst11.dutycycle_RNIK9J85_5_LC_7_11_3  (
            .in0(N__25059),
            .in1(N__26883),
            .in2(N__25083),
            .in3(N__36019),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_172_m3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIRO179_3_LC_7_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIRO179_3_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIRO179_3_LC_7_11_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \b2v_inst11.dutycycle_RNIRO179_3_LC_7_11_4  (
            .in0(N__26898),
            .in1(N__25080),
            .in2(N__25074),
            .in3(N__26952),
            .lcout(\b2v_inst11.un1_dutycycle_172_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_6_1_LC_7_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_6_1_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_6_1_LC_7_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.func_state_RNI_6_1_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__38850),
            .in2(_gnd_net_),
            .in3(N__34032),
            .lcout(\b2v_inst11.N_19_i ),
            .ltout(\b2v_inst11.N_19_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNII7Q52_5_LC_7_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNII7Q52_5_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNII7Q52_5_LC_7_11_6 .LUT_INIT=16'b0000001011110010;
    LogicCell40 \b2v_inst11.dutycycle_RNII7Q52_5_LC_7_11_6  (
            .in0(N__38484),
            .in1(N__38615),
            .in2(N__25065),
            .in3(N__26877),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_172_m0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_5_LC_7_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_5_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_5_LC_7_11_7 .LUT_INIT=16'b0011111100101100;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_5_LC_7_11_7  (
            .in0(N__34823),
            .in1(N__28858),
            .in2(N__25062),
            .in3(N__36020),
            .lcout(\b2v_inst11.un1_dutycycle_172_m0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_0  (
            .in0(N__38346),
            .in1(N__29276),
            .in2(_gnd_net_),
            .in3(N__28956),
            .lcout(),
            .ltout(\b2v_inst11.g0_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_0_LC_7_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_0_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_0_LC_7_12_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_0_LC_7_12_1  (
            .in0(N__31454),
            .in1(N__31577),
            .in2(N__25053),
            .in3(N__37749),
            .lcout(\b2v_inst11.N_293_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_0_LC_7_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_0_LC_7_12_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_0_LC_7_12_2  (
            .in0(N__34024),
            .in1(N__25113),
            .in2(N__31583),
            .in3(N__31453),
            .lcout(\b2v_inst11.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_12_LC_7_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_12_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_12_LC_7_12_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_12_LC_7_12_3  (
            .in0(N__29278),
            .in1(N__37747),
            .in2(N__28964),
            .in3(N__38347),
            .lcout(\b2v_inst11.g0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_12_LC_7_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_12_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_12_LC_7_12_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_12_LC_7_12_4  (
            .in0(N__37748),
            .in1(N__29279),
            .in2(N__38352),
            .in3(N__28960),
            .lcout(\b2v_inst11.g0_3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_13_LC_7_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_13_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_13_LC_7_12_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_13_LC_7_12_5  (
            .in0(N__34591),
            .in1(N__35084),
            .in2(N__37935),
            .in3(N__35193),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_15_LC_7_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_15_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_15_LC_7_12_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_15_LC_7_12_6  (
            .in0(N__29331),
            .in1(N__38168),
            .in2(N__25107),
            .in3(N__37594),
            .lcout(\b2v_inst11.N_363 ),
            .ltout(\b2v_inst11.N_363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_7_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_7_12_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_12_LC_7_12_7  (
            .in0(N__29277),
            .in1(_gnd_net_),
            .in2(N__25104),
            .in3(N__37746),
            .lcout(\b2v_inst11.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27248),
            .lcout(\b2v_inst11.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27185),
            .lcout(\b2v_inst11.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_7_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_7_13_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_8_LC_7_13_3  (
            .in0(N__39055),
            .in1(N__37930),
            .in2(_gnd_net_),
            .in3(N__32310),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_1_LC_7_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_1_LC_7_13_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_1_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27288),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_3_sf_LC_7_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_3_sf_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_3_sf_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_3_sf_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29446),
            .lcout(\b2v_inst11.mult1_un54_sum_s_3_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25155),
            .in3(N__25146),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29394),
            .in3(N__25143),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__30946),
            .in2(N__29460),
            .in3(N__25140),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__30947),
            .in2(N__29493),
            .in3(N__25137),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_7_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_7_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__27408),
            .in2(_gnd_net_),
            .in3(N__25134),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25131),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25261),
            .lcout(\b2v_inst11.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27438),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__25262),
            .in2(N__25128),
            .in3(N__25116),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__25272),
            .in2(N__25266),
            .in3(N__25248),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__25198),
            .in2(N__25245),
            .in3(N__25236),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__25233),
            .in2(N__25205),
            .in3(N__25227),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_15_5  (
            .in0(N__25321),
            .in1(N__25224),
            .in2(N__25185),
            .in3(N__25218),
            .lcout(\b2v_inst11.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_15_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_15_6  (
            .in0(N__25215),
            .in1(N__27407),
            .in2(N__25206),
            .in3(N__25209),
            .lcout(\b2v_inst11.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25197),
            .lcout(\b2v_inst11.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27311),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_16_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__27423),
            .in2(N__25295),
            .in3(N__25167),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_7_16_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_7_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__25291),
            .in2(N__25164),
            .in3(N__25428),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_7_16_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_7_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__25317),
            .in2(N__25425),
            .in3(N__25410),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_7_16_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_7_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__25407),
            .in2(N__25325),
            .in3(N__25395),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_7_16_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_7_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_7_16_5  (
            .in0(N__25351),
            .in1(N__25392),
            .in2(N__25296),
            .in3(N__25377),
            .lcout(\b2v_inst11.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_7_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_7_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25374),
            .in3(N__25365),
            .lcout(\b2v_inst11.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_7_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_7_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25316),
            .lcout(\b2v_inst11.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNI440L1_LC_8_1_0 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNI440L1_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNI440L1_LC_8_1_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_c_RNI440L1_LC_8_1_0  (
            .in0(N__33137),
            .in1(N__29717),
            .in2(N__29738),
            .in3(N__29780),
            .lcout(\b2v_inst6.count_rst_11 ),
            .ltout(\b2v_inst6.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNINOEF5_3_LC_8_1_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNINOEF5_3_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNINOEF5_3_LC_8_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNINOEF5_3_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__25508),
            .in2(N__25278),
            .in3(N__33450),
            .lcout(\b2v_inst6.un2_count_1_axb_3 ),
            .ltout(\b2v_inst6.un2_count_1_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_3_LC_8_1_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_3_LC_8_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_3_LC_8_1_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.count_3_LC_8_1_2  (
            .in0(N__33140),
            .in1(N__29718),
            .in2(N__25275),
            .in3(N__29783),
            .lcout(\b2v_inst6.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36437),
            .ce(N__33456),
            .sr(N__33236));
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNI561L1_LC_8_1_3 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNI561L1_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNI561L1_LC_8_1_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_c_RNI561L1_LC_8_1_3  (
            .in0(N__29781),
            .in1(N__29672),
            .in2(N__29699),
            .in3(N__33138),
            .lcout(\b2v_inst6.count_rst_10 ),
            .ltout(\b2v_inst6.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIPRFF5_4_LC_8_1_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIPRFF5_4_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIPRFF5_4_LC_8_1_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNIPRFF5_4_LC_8_1_4  (
            .in0(N__33451),
            .in1(_gnd_net_),
            .in2(N__25518),
            .in3(N__25490),
            .lcout(\b2v_inst6.un2_count_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNINOEF5_0_3_LC_8_1_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNINOEF5_0_3_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNINOEF5_0_3_LC_8_1_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst6.count_RNINOEF5_0_3_LC_8_1_5  (
            .in0(N__25515),
            .in1(N__25509),
            .in2(_gnd_net_),
            .in3(N__33453),
            .lcout(),
            .ltout(\b2v_inst6.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIGKUUA_4_LC_8_1_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIGKUUA_4_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIGKUUA_4_LC_8_1_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \b2v_inst6.count_RNIGKUUA_4_LC_8_1_6  (
            .in0(N__33452),
            .in1(N__25500),
            .in2(N__25494),
            .in3(N__25491),
            .lcout(\b2v_inst6.count_1_i_a3_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_4_LC_8_1_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_4_LC_8_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_4_LC_8_1_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.count_4_LC_8_1_7  (
            .in0(N__29782),
            .in1(N__33139),
            .in2(N__29698),
            .in3(N__29673),
            .lcout(\b2v_inst6.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36437),
            .ce(N__33456),
            .sr(N__33236));
    defparam \b2v_inst5.count_7_LC_8_2_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_7_LC_8_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_7_LC_8_2_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst5.count_7_LC_8_2_0  (
            .in0(N__25464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25963),
            .lcout(\b2v_inst5.count_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36834),
            .ce(N__26276),
            .sr(N__25998));
    defparam \b2v_inst5.count_RNID0AN3_11_LC_8_2_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNID0AN3_11_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNID0AN3_11_LC_8_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst5.count_RNID0AN3_11_LC_8_2_1  (
            .in0(N__26262),
            .in1(N__25694),
            .in2(_gnd_net_),
            .in3(N__25711),
            .lcout(\b2v_inst5.un2_count_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_11_LC_8_2_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_11_LC_8_2_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_11_LC_8_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_11_LC_8_2_2  (
            .in0(N__25713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36834),
            .ce(N__26276),
            .sr(N__25998));
    defparam \b2v_inst5.count_RNIN9BH3_7_LC_8_2_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIN9BH3_7_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIN9BH3_7_LC_8_2_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \b2v_inst5.count_RNIN9BH3_7_LC_8_2_3  (
            .in0(N__25960),
            .in1(N__25470),
            .in2(N__26277),
            .in3(N__25463),
            .lcout(\b2v_inst5.countZ0Z_7 ),
            .ltout(\b2v_inst5.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNID0AN3_0_11_LC_8_2_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNID0AN3_0_11_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNID0AN3_0_11_LC_8_2_4 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \b2v_inst5.count_RNID0AN3_0_11_LC_8_2_4  (
            .in0(N__25712),
            .in1(N__25695),
            .in2(N__25683),
            .in3(N__26263),
            .lcout(\b2v_inst5.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_2_LC_8_2_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_2_LC_8_2_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_2_LC_8_2_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst5.count_2_LC_8_2_5  (
            .in0(N__25961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25680),
            .lcout(\b2v_inst5.count_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36834),
            .ce(N__26276),
            .sr(N__25998));
    defparam \b2v_inst5.count_RNIDQ5H3_2_LC_8_2_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIDQ5H3_2_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIDQ5H3_2_LC_8_2_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst5.count_RNIDQ5H3_2_LC_8_2_6  (
            .in0(N__25679),
            .in1(N__26258),
            .in2(N__25665),
            .in3(N__25959),
            .lcout(\b2v_inst5.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_3_LC_8_2_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_3_LC_8_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_3_LC_8_2_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst5.count_3_LC_8_2_7  (
            .in0(N__25962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25635),
            .lcout(\b2v_inst5.count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36834),
            .ce(N__26276),
            .sr(N__25998));
    defparam \b2v_inst5.count_RNI7BCA2_10_LC_8_3_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI7BCA2_10_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI7BCA2_10_LC_8_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst5.count_RNI7BCA2_10_LC_8_3_0  (
            .in0(N__26253),
            .in1(N__25524),
            .in2(_gnd_net_),
            .in3(N__26352),
            .lcout(\b2v_inst5.un2_count_1_axb_10 ),
            .ltout(\b2v_inst5.un2_count_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_10_LC_8_3_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_10_LC_8_3_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_10_LC_8_3_1 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_10_LC_8_3_1  (
            .in0(N__25541),
            .in1(N__25975),
            .in2(N__25605),
            .in3(N__26086),
            .lcout(\b2v_inst5.count_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37014),
            .ce(N__26306),
            .sr(N__25980));
    defparam \b2v_inst5.count_RNI3QEK5_11_LC_8_3_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI3QEK5_11_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI3QEK5_11_LC_8_3_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst5.count_RNI3QEK5_11_LC_8_3_2  (
            .in0(N__25602),
            .in1(N__25596),
            .in2(N__25584),
            .in3(N__25575),
            .lcout(\b2v_inst5.un12_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_8_3_3 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_8_3_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_8_3_3  (
            .in0(N__25556),
            .in1(N__25974),
            .in2(N__25542),
            .in3(N__26085),
            .lcout(\b2v_inst5.count_rst_4 ),
            .ltout(\b2v_inst5.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI7BCA2_0_10_LC_8_3_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI7BCA2_0_10_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI7BCA2_0_10_LC_8_3_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \b2v_inst5.count_RNI7BCA2_0_10_LC_8_3_4  (
            .in0(N__26254),
            .in1(N__26351),
            .in2(N__26343),
            .in3(N__26016),
            .lcout(),
            .ltout(\b2v_inst5.un12_clk_100khz_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI870S9_8_LC_8_3_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI870S9_8_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI870S9_8_LC_8_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.count_RNI870S9_8_LC_8_3_5  (
            .in0(N__26340),
            .in1(N__26328),
            .in2(N__26322),
            .in3(N__26319),
            .lcout(\b2v_inst5.N_1_i ),
            .ltout(\b2v_inst5.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_9_LC_8_3_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_9_LC_8_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_9_LC_8_3_6 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst5.count_9_LC_8_3_6  (
            .in0(N__26046),
            .in1(N__25981),
            .in2(N__26313),
            .in3(N__26017),
            .lcout(\b2v_inst5.count_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37014),
            .ce(N__26306),
            .sr(N__25980));
    defparam \b2v_inst5.count_RNIRFDH3_9_LC_8_3_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRFDH3_9_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRFDH3_9_LC_8_3_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \b2v_inst5.count_RNIRFDH3_9_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__26255),
            .in2(N__26172),
            .in3(N__25794),
            .lcout(\b2v_inst5.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_4_0 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_4_0 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_4_0  (
            .in0(N__26162),
            .in1(N__26135),
            .in2(N__25896),
            .in3(N__26087),
            .lcout(\b2v_inst5.count_rst_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_8_4_1 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_8_4_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_8_4_1  (
            .in0(N__26088),
            .in1(N__26045),
            .in2(N__26027),
            .in3(N__25849),
            .lcout(\b2v_inst5.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_8_4_2 .C_ON=1'b0;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_8_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.un8_rsmrst_pwrgd_4_LC_8_4_2  (
            .in0(N__25788),
            .in1(N__25773),
            .in2(N__25761),
            .in3(N__25740),
            .lcout(SYNTHESIZED_WIRE_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI_1_LC_8_4_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI_1_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI_1_LC_8_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.curr_state_RNI_1_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27466),
            .lcout(\b2v_inst6.N_3011_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_8_4_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_8_4_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_8_4_4  (
            .in0(N__25728),
            .in1(N__38730),
            .in2(N__26394),
            .in3(N__34817),
            .lcout(\b2v_inst6.N_192 ),
            .ltout(\b2v_inst6.N_192_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_8_4_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_8_4_5 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_8_4_5  (
            .in0(N__27645),
            .in1(_gnd_net_),
            .in2(N__26373),
            .in3(N__27861),
            .lcout(\b2v_inst6.N_241 ),
            .ltout(\b2v_inst6.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_1_LC_8_4_6 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_1_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_1_LC_8_4_6 .LUT_INIT=16'b0000010100001111;
    LogicCell40 \b2v_inst6.curr_state_1_LC_8_4_6  (
            .in0(N__27467),
            .in1(_gnd_net_),
            .in2(N__26370),
            .in3(N__29820),
            .lcout(\b2v_inst6.curr_state_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36836),
            .ce(N__27545),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIG8KAH_7_LC_8_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIG8KAH_7_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIG8KAH_7_LC_8_5_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.count_clk_RNIG8KAH_7_LC_8_5_0  (
            .in0(N__30153),
            .in1(N__29977),
            .in2(_gnd_net_),
            .in3(N__26361),
            .lcout(),
            .ltout(\b2v_inst11.count_clk_RNIG8KAHZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNITV5AU_7_LC_8_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNITV5AU_7_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNITV5AU_7_LC_8_5_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.count_clk_RNITV5AU_7_LC_8_5_1  (
            .in0(N__27948),
            .in1(N__30440),
            .in2(N__26367),
            .in3(N__32296),
            .lcout(\b2v_inst11.count_clk_RNITV5AUZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI7SOFB_1_LC_8_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI7SOFB_1_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI7SOFB_1_LC_8_5_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \b2v_inst11.count_clk_RNI7SOFB_1_LC_8_5_2  (
            .in0(N__30479),
            .in1(N__27958),
            .in2(N__32946),
            .in3(N__29978),
            .lcout(\b2v_inst11.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIB2RFB_1_LC_8_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIB2RFB_1_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIB2RFB_1_LC_8_5_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst11.count_clk_RNIB2RFB_1_LC_8_5_3  (
            .in0(N__27960),
            .in1(N__30151),
            .in2(_gnd_net_),
            .in3(N__30480),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIG510T_5_LC_8_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIG510T_5_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIG510T_5_LC_8_5_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.count_clk_RNIG510T_5_LC_8_5_4  (
            .in0(N__32945),
            .in1(N__27947),
            .in2(N__26364),
            .in3(N__29979),
            .lcout(\b2v_inst11.count_clk_RNIG510TZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI7SOFB_0_1_LC_8_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI7SOFB_0_1_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI7SOFB_0_1_LC_8_5_5 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \b2v_inst11.count_clk_RNI7SOFB_0_1_LC_8_5_5  (
            .in0(N__27959),
            .in1(N__32944),
            .in2(_gnd_net_),
            .in3(N__30478),
            .lcout(\b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1 ),
            .ltout(\b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIG510T_0_7_LC_8_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIG510T_0_7_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIG510T_0_7_LC_8_5_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst11.count_clk_RNIG510T_0_7_LC_8_5_6  (
            .in0(N__30152),
            .in1(N__27946),
            .in2(N__26355),
            .in3(N__29976),
            .lcout(\b2v_inst11.N_428 ),
            .ltout(\b2v_inst11.N_428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_3_LC_8_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_3_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_3_LC_8_5_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_3_LC_8_5_7  (
            .in0(N__39094),
            .in1(N__30441),
            .in2(N__26565),
            .in3(N__32297),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_332_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.N_224_i_LC_8_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.N_224_i_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.N_224_i_LC_8_6_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.N_224_i_LC_8_6_0  (
            .in0(N__39284),
            .in1(N__34771),
            .in2(N__38417),
            .in3(N__28328),
            .lcout(\b2v_inst11.N_224_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNILG61T1_5_LC_8_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNILG61T1_5_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNILG61T1_5_LC_8_6_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst11.count_clk_RNILG61T1_5_LC_8_6_1  (
            .in0(N__28579),
            .in1(N__27990),
            .in2(N__26601),
            .in3(N__26562),
            .lcout(\b2v_inst11.count_clk_RNILG61T1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_8_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_8_6_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_8_6_2  (
            .in0(N__39285),
            .in1(N__34769),
            .in2(N__38418),
            .in3(N__28326),
            .lcout(\b2v_inst11.N_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_4_i_a2_sx_LC_8_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_4_i_a2_sx_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_4_i_a2_sx_LC_8_6_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \b2v_inst11.un1_func_state25_4_i_a2_sx_LC_8_6_3  (
            .in0(N__38722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39286),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_4_i_a2_sxZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_4_i_a2_LC_8_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_4_i_a2_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_4_i_a2_LC_8_6_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \b2v_inst11.un1_func_state25_4_i_a2_LC_8_6_4  (
            .in0(N__28770),
            .in1(N__28142),
            .in2(N__26412),
            .in3(N__28085),
            .lcout(\b2v_inst11.N_417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_6_5 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_6_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__28078),
            .in2(N__28146),
            .in3(N__28769),
            .lcout(rsmrstn),
            .ltout(rsmrstn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_8_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_8_6_6 .LUT_INIT=16'b0001111110011111;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_8_6_6  (
            .in0(N__38563),
            .in1(N__38718),
            .in2(N__26409),
            .in3(N__28327),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNI1EKN3_LC_8_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNI1EKN3_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNI1EKN3_LC_8_6_7 .LUT_INIT=16'b1111111101010111;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNI1EKN3_LC_8_6_7  (
            .in0(N__34770),
            .in1(N__38564),
            .in2(N__38729),
            .in3(N__26406),
            .lcout(\b2v_inst11.N_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_8_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_8_7_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_8_7_0  (
            .in0(N__30749),
            .in1(N__28158),
            .in2(_gnd_net_),
            .in3(N__34059),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_331_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_fast_LC_8_7_1 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_fast_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_fast_LC_8_7_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst20.tmp_1_fast_LC_8_7_1  (
            .in0(N__28145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26681),
            .lcout(SYNTHESIZED_WIRE_1keep_3_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36969),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_2_1_LC_8_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_8_7_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.func_state_RNI_2_1_LC_8_7_2  (
            .in0(N__30747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39053),
            .lcout(\b2v_inst11.func_state_RNI_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI5DLR_1_LC_8_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI5DLR_1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI5DLR_1_LC_8_7_3 .LUT_INIT=16'b1010000000010001;
    LogicCell40 \b2v_inst11.func_state_RNI5DLR_1_LC_8_7_3  (
            .in0(N__32276),
            .in1(N__38981),
            .in2(N__28734),
            .in3(N__30748),
            .lcout(\b2v_inst11.func_state_1_ss0_i_0_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_1_LC_8_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_1_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_1_LC_8_7_4 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_1_LC_8_7_4  (
            .in0(N__38724),
            .in1(N__39288),
            .in2(N__30377),
            .in3(N__32277),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_8_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_8_7_5 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_8_7_5  (
            .in0(N__26777),
            .in1(N__26619),
            .in2(N__26613),
            .in3(N__26610),
            .lcout(\b2v_inst11.un1_func_state25_6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_8_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_8_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_8_7_6  (
            .in0(N__26597),
            .in1(N__28733),
            .in2(N__34818),
            .in3(N__32274),
            .lcout(),
            .ltout(\b2v_inst11.N_337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_8_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_8_7_7 .LUT_INIT=16'b1111001111110001;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_8_7_7  (
            .in0(N__32275),
            .in1(N__38980),
            .in2(N__26586),
            .in3(N__28892),
            .lcout(\b2v_inst11.func_state_1_m2s2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNITU8B9_0_LC_8_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNITU8B9_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNITU8B9_0_LC_8_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.func_state_RNITU8B9_0_LC_8_8_0  (
            .in0(N__28017),
            .in1(N__26577),
            .in2(_gnd_net_),
            .in3(N__26571),
            .lcout(\b2v_inst11.func_state_1_m2_0 ),
            .ltout(\b2v_inst11.func_state_1_m2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIM28UB_0_LC_8_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIM28UB_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIM28UB_0_LC_8_8_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst11.func_state_RNIM28UB_0_LC_8_8_1  (
            .in0(N__26775),
            .in1(N__26747),
            .in2(N__26796),
            .in3(N__26734),
            .lcout(\b2v_inst11.func_stateZ0Z_0 ),
            .ltout(\b2v_inst11.func_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_0_LC_8_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_0_LC_8_8_2 .LUT_INIT=16'b1011111111001100;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_0_LC_8_8_2  (
            .in0(N__39294),
            .in1(N__38560),
            .in2(N__26793),
            .in3(N__38693),
            .lcout(\b2v_inst11.g3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_LC_8_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_8_8_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_LC_8_8_3  (
            .in0(N__38967),
            .in1(N__31395),
            .in2(_gnd_net_),
            .in3(N__32249),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_LC_8_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_0_LC_8_8_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst11.func_state_0_LC_8_8_4  (
            .in0(N__26748),
            .in1(N__26790),
            .in2(N__26739),
            .in3(N__26776),
            .lcout(\b2v_inst11.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36980),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_8_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_8_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29224),
            .lcout(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI6M5R2_1_LC_8_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI6M5R2_1_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI6M5R2_1_LC_8_8_6 .LUT_INIT=16'b1111010101010101;
    LogicCell40 \b2v_inst11.func_state_RNI6M5R2_1_LC_8_8_6  (
            .in0(N__26735),
            .in1(_gnd_net_),
            .in2(N__26715),
            .in3(N__37402),
            .lcout(\b2v_inst11.func_state_RNI6M5R2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a3_1_LC_8_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a3_1_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a3_1_LC_8_8_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \b2v_inst11.un1_clk_100khz_52_and_i_a3_1_LC_8_8_7  (
            .in0(N__38561),
            .in1(_gnd_net_),
            .in2(N__38717),
            .in3(N__34801),
            .lcout(\b2v_inst11.un1_clk_100khz_25_and_i_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_8_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_8_9_0 .LUT_INIT=16'b1100001111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_2_LC_8_9_0  (
            .in0(N__31297),
            .in1(N__26712),
            .in2(N__26706),
            .in3(N__31423),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_8_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_8_9_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_4_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__26854),
            .in2(_gnd_net_),
            .in3(N__35002),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_8_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_8_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_3_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__34362),
            .in2(_gnd_net_),
            .in3(N__38310),
            .lcout(\b2v_inst11.d_N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQH45K_5_LC_8_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQH45K_5_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQH45K_5_LC_8_9_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIQH45K_5_LC_8_9_3  (
            .in0(N__34455),
            .in1(N__35789),
            .in2(N__33924),
            .in3(N__34466),
            .lcout(\b2v_inst11.dutycycleZ1Z_5 ),
            .ltout(\b2v_inst11.dutycycleZ1Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_8_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_8_9_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_5_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26838),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ),
            .ltout(\b2v_inst11.dutycycle_RNI_1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_8_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_8_9_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_0_LC_8_9_5  (
            .in0(N__38311),
            .in1(N__31463),
            .in2(N__26835),
            .in3(N__31532),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_0_LC_8_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_0_LC_8_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_0_LC_8_9_6  (
            .in0(N__31533),
            .in1(N__31424),
            .in2(N__26823),
            .in3(N__38312),
            .lcout(\b2v_inst11.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_0_LC_8_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_0_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_0_LC_8_9_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_0_LC_8_9_7  (
            .in0(N__31425),
            .in1(N__31534),
            .in2(N__38343),
            .in3(N__26819),
            .lcout(\b2v_inst11.dutycycle_RNI_9Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_2_LC_8_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_2_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_2_LC_8_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_2_LC_8_10_0  (
            .in0(N__28902),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28666),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_LC_8_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_LC_8_10_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_LC_8_10_1  (
            .in0(N__28629),
            .in1(N__30637),
            .in2(N__32307),
            .in3(N__28901),
            .lcout(\b2v_inst11.N_159 ),
            .ltout(\b2v_inst11.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_2_LC_8_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_2_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_2_LC_8_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_2_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26799),
            .in3(N__28670),
            .lcout(\b2v_inst11.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_1_2_LC_8_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_1_2_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_1_2_LC_8_10_3 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_1_2_LC_8_10_3  (
            .in0(N__28630),
            .in1(N__30438),
            .in2(N__28678),
            .in3(N__34183),
            .lcout(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_0_LC_8_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_0_LC_8_10_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_0_LC_8_10_4  (
            .in0(N__26855),
            .in1(N__38847),
            .in2(_gnd_net_),
            .in3(N__26892),
            .lcout(\b2v_inst11.dutycycle_RNI_11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_8_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_8_10_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_14_LC_8_10_5  (
            .in0(N__32284),
            .in1(_gnd_net_),
            .in2(N__39093),
            .in3(N__35211),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_10_LC_8_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_10_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_10_LC_8_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_10_LC_8_10_6  (
            .in0(N__35472),
            .in1(N__39012),
            .in2(_gnd_net_),
            .in3(N__32282),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_8_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_8_10_7 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_13_LC_8_10_7  (
            .in0(N__32283),
            .in1(_gnd_net_),
            .in2(N__39092),
            .in3(N__34605),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_0_2_LC_8_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_0_2_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_0_2_LC_8_11_0 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_0_2_LC_8_11_0  (
            .in0(N__32292),
            .in1(N__26946),
            .in2(N__31290),
            .in3(N__36175),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_172_m3_d_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_2_LC_8_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_2_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_2_LC_8_11_1 .LUT_INIT=16'b0000000111100001;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_2_LC_8_11_1  (
            .in0(N__26931),
            .in1(N__26915),
            .in2(N__26886),
            .in3(N__30429),
            .lcout(\b2v_inst11.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_8_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_8_11_2 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_8_11_2  (
            .in0(N__32294),
            .in1(N__26862),
            .in2(_gnd_net_),
            .in3(N__36177),
            .lcout(\b2v_inst11.dutycycle_RNIDQ4A1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_2_LC_8_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_2_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_2_LC_8_11_3 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_2_LC_8_11_3  (
            .in0(N__36176),
            .in1(N__27015),
            .in2(N__31291),
            .in3(N__32293),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_172_m4_rn_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQK9K2_0_2_LC_8_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_0_2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQK9K2_0_2_LC_8_11_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIQK9K2_0_2_LC_8_11_4  (
            .in0(N__32295),
            .in1(N__36178),
            .in2(N__26871),
            .in3(N__26868),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_172_m4_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI7FEU3_0_LC_8_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI7FEU3_0_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI7FEU3_0_LC_8_11_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI7FEU3_0_LC_8_11_5  (
            .in0(N__26861),
            .in1(N__27014),
            .in2(N__26955),
            .in3(N__30428),
            .lcout(\b2v_inst11.un1_dutycycle_172_m4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_16_0_LC_8_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_16_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_16_0_LC_8_11_6 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_16_0_LC_8_11_6  (
            .in0(N__26916),
            .in1(N__26939),
            .in2(N__34193),
            .in3(N__28861),
            .lcout(\b2v_inst11.N_3057_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_17_0_LC_8_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_17_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_17_0_LC_8_11_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_17_0_LC_8_11_7  (
            .in0(N__26940),
            .in1(N__28862),
            .in2(_gnd_net_),
            .in3(N__34187),
            .lcout(\b2v_inst11.N_3055_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_8_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_8_12_0 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_3_LC_8_12_0  (
            .in0(N__34388),
            .in1(_gnd_net_),
            .in2(N__38859),
            .in3(N__34986),
            .lcout(\b2v_inst11.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__29241),
            .in2(_gnd_net_),
            .in3(N__38851),
            .lcout(),
            .ltout(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5AV24_4_LC_8_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5AV24_4_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5AV24_4_LC_8_12_2 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \b2v_inst11.dutycycle_RNI5AV24_4_LC_8_12_2  (
            .in0(N__34976),
            .in1(N__37508),
            .in2(N__26925),
            .in3(N__37408),
            .lcout(\b2v_inst11.dutycycle_RNI5AV24Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_8_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_8_12_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_0_LC_8_12_3  (
            .in0(N__31554),
            .in1(N__26922),
            .in2(N__34047),
            .in3(N__31449),
            .lcout(\b2v_inst11.g1_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_LC_8_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_8_12_4 .LUT_INIT=16'b0000000011111101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_LC_8_12_4  (
            .in0(N__26907),
            .in1(N__31552),
            .in2(N__31462),
            .in3(N__34188),
            .lcout(),
            .ltout(\b2v_inst11.g2_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_LC_8_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_8_12_5 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_LC_8_12_5  (
            .in0(N__29178),
            .in1(N__34978),
            .in2(N__26901),
            .in3(N__34387),
            .lcout(\b2v_inst11.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_0_LC_8_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_0_LC_8_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_0_LC_8_12_6  (
            .in0(N__31448),
            .in1(N__31553),
            .in2(N__38858),
            .in3(N__29327),
            .lcout(\b2v_inst11.dutycycle_RNI_10Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_8_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_8_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_0_LC_8_12_7  (
            .in0(N__31555),
            .in1(N__34977),
            .in2(_gnd_net_),
            .in3(N__31444),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIPKS23_4_LC_8_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIPKS23_4_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIPKS23_4_LC_8_13_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNIPKS23_4_LC_8_13_0  (
            .in0(N__35799),
            .in1(N__36173),
            .in2(N__26997),
            .in3(N__27003),
            .lcout(\b2v_inst11.dutycycle_RNIPKS23Z0Z_4 ),
            .ltout(\b2v_inst11.dutycycle_RNIPKS23Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_4_LC_8_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_4_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_4_LC_8_13_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \b2v_inst11.dutycycle_4_LC_8_13_1  (
            .in0(N__26982),
            .in1(N__37361),
            .in2(N__27006),
            .in3(N__26996),
            .lcout(\b2v_inst11.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37069),
            .ce(),
            .sr(N__36341));
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_8_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_8_13_2 .LUT_INIT=16'b1111010100001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_2_LC_8_13_2  (
            .in0(N__31443),
            .in1(N__31299),
            .in2(N__35009),
            .in3(N__36011),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08U_LC_8_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08U_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08U_LC_8_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08U_LC_8_13_3  (
            .in0(N__31128),
            .in1(N__30969),
            .in2(_gnd_net_),
            .in3(N__36010),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08UZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIM7549_4_LC_8_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIM7549_4_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIM7549_4_LC_8_13_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \b2v_inst11.dutycycle_RNIM7549_4_LC_8_13_4  (
            .in0(N__26995),
            .in1(N__26981),
            .in2(N__37362),
            .in3(N__26973),
            .lcout(\b2v_inst11.dutycycleZ0Z_6 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_8_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_8_13_5 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_3_LC_8_13_5  (
            .in0(N__38345),
            .in1(N__31442),
            .in2(N__26967),
            .in3(N__34381),
            .lcout(),
            .ltout(\b2v_inst11.un1_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_LC_8_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_8_13_6 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_LC_8_13_6  (
            .in0(N__29529),
            .in1(N__26961),
            .in2(N__26964),
            .in3(N__36012),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_13_7 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_3_LC_8_13_7  (
            .in0(N__38344),
            .in1(N__31441),
            .in2(_gnd_net_),
            .in3(N__34380),
            .lcout(\b2v_inst11.d_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_8_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_8_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_0_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__34389),
            .in2(N__31581),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_0 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_8_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_8_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__31570),
            .in2(N__27234),
            .in3(N__27195),
            .lcout(\b2v_inst11.mult1_un138_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_8_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_8_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__27192),
            .in2(N__31301),
            .in3(N__27165),
            .lcout(\b2v_inst11.mult1_un131_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_1 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_8_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_8_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__31289),
            .in2(N__27162),
            .in3(N__27126),
            .lcout(\b2v_inst11.mult1_un124_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_2 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_8_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_8_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__29525),
            .in2(N__27123),
            .in3(N__27093),
            .lcout(\b2v_inst11.mult1_un117_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_3 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_8_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_8_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__29514),
            .in2(N__36060),
            .in3(N__27072),
            .lcout(\b2v_inst11.mult1_un110_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_4 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_8_14_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_8_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__31746),
            .in2(N__36061),
            .in3(N__27042),
            .lcout(\b2v_inst11.mult1_un103_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_5 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_8_14_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_8_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__35468),
            .in2(N__32028),
            .in3(N__27018),
            .lcout(\b2v_inst11.mult1_un96_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_6 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_8_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_8_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__31969),
            .in2(N__31872),
            .in3(N__27363),
            .lcout(\b2v_inst11.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_8_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_8_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__37766),
            .in2(N__37653),
            .in3(N__27342),
            .lcout(\b2v_inst11.mult1_un82_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_8 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_8_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_8_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__34600),
            .in2(N__27417),
            .in3(N__27318),
            .lcout(\b2v_inst11.mult1_un75_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_9 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_8_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_8_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__29592),
            .in2(N__35210),
            .in3(N__27294),
            .lcout(\b2v_inst11.mult1_un68_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_8_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_8_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__29379),
            .in2(N__37595),
            .in3(N__27291),
            .lcout(\b2v_inst11.mult1_un61_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_8_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_8_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__31794),
            .in2(N__34608),
            .in3(N__27267),
            .lcout(\b2v_inst11.mult1_un47_sum_1 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_8_15_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_8_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__35203),
            .in2(N__31758),
            .in3(N__27264),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_8_15_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_8_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__37588),
            .in2(N__29586),
            .in3(N__27261),
            .lcout(\b2v_inst11.mult1_un40_sum_i_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_8_16_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_8_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__37589),
            .in2(N__29577),
            .in3(N__27258),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\b2v_inst11.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_8_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_8_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.CO2_THRU_LUT4_0_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27441),
            .lcout(\b2v_inst11.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27437),
            .lcout(\b2v_inst11.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_13_LC_8_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_8_16_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_13_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29538),
            .in3(N__34604),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_m_0_6_LC_8_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_m_0_6_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_m_0_6_LC_8_16_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_m_0_6_LC_8_16_6  (
            .in0(N__29414),
            .in1(N__29507),
            .in2(N__29448),
            .in3(N__29476),
            .lcout(\b2v_inst11.mult1_un47_sum_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_8_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_8_16_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__27389),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_9_LC_9_1_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_9_LC_9_1_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_9_LC_9_1_0 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst6.count_9_LC_9_1_0  (
            .in0(N__29894),
            .in1(N__29796),
            .in2(N__33209),
            .in3(N__29877),
            .lcout(\b2v_inst6.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36709),
            .ce(N__33463),
            .sr(N__33237));
    defparam \b2v_inst6.count_RNI18KF5_8_LC_9_1_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI18KF5_8_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI18KF5_8_LC_9_1_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNI18KF5_8_LC_9_1_1  (
            .in0(N__27575),
            .in1(N__27605),
            .in2(_gnd_net_),
            .in3(N__33460),
            .lcout(\b2v_inst6.un2_count_1_axb_8 ),
            .ltout(\b2v_inst6.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNI9E5L1_LC_9_1_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNI9E5L1_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNI9E5L1_LC_9_1_2 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_c_RNI9E5L1_LC_9_1_2  (
            .in0(N__33141),
            .in1(N__29793),
            .in2(N__27366),
            .in3(N__29912),
            .lcout(\b2v_inst6.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI3BLF5_9_LC_9_1_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI3BLF5_9_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI3BLF5_9_LC_9_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNI3BLF5_9_LC_9_1_3  (
            .in0(N__27584),
            .in1(N__27596),
            .in2(_gnd_net_),
            .in3(N__33461),
            .lcout(\b2v_inst6.un2_count_1_axb_9 ),
            .ltout(\b2v_inst6.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIAG6L1_LC_9_1_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIAG6L1_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIAG6L1_LC_9_1_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_c_RNIAG6L1_LC_9_1_4  (
            .in0(N__33142),
            .in1(N__29794),
            .in2(N__27609),
            .in3(N__29876),
            .lcout(\b2v_inst6.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI18KF5_0_8_LC_9_1_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI18KF5_0_8_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI18KF5_0_8_LC_9_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNI18KF5_0_8_LC_9_1_5  (
            .in0(N__27576),
            .in1(N__27606),
            .in2(_gnd_net_),
            .in3(N__33464),
            .lcout(),
            .ltout(\b2v_inst6.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI4J9VA_9_LC_9_1_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI4J9VA_9_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI4J9VA_9_LC_9_1_6 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \b2v_inst6.count_RNI4J9VA_9_LC_9_1_6  (
            .in0(N__27597),
            .in1(N__33462),
            .in2(N__27588),
            .in3(N__27585),
            .lcout(\b2v_inst6.count_1_i_a3_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_8_LC_9_1_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_8_LC_9_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_8_LC_9_1_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.count_8_LC_9_1_7  (
            .in0(N__29795),
            .in1(N__33143),
            .in2(N__29916),
            .in3(N__29930),
            .lcout(\b2v_inst6.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36709),
            .ce(N__33463),
            .sr(N__33237));
    defparam \b2v_inst6.curr_state_0_LC_9_2_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_0_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_0_LC_9_2_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \b2v_inst6.curr_state_0_LC_9_2_0  (
            .in0(N__29813),
            .in1(N__27875),
            .in2(N__27468),
            .in3(N__27626),
            .lcout(\b2v_inst6.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36835),
            .ce(N__27546),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_0_0_LC_9_2_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_0_0_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_0_0_LC_9_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst6.count_RNI_0_0_LC_9_2_1  (
            .in0(N__33530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33551),
            .lcout(\b2v_inst6.N_394 ),
            .ltout(\b2v_inst6.N_394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_9_2_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_9_2_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_9_2_2  (
            .in0(N__27465),
            .in1(_gnd_net_),
            .in2(N__27483),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst6.m6_i_a3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIS68V1_1_LC_9_2_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIS68V1_1_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIS68V1_1_LC_9_2_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \b2v_inst6.curr_state_RNIS68V1_1_LC_9_2_3  (
            .in0(N__27480),
            .in1(N__33611),
            .in2(N__27471),
            .in3(N__28382),
            .lcout(\b2v_inst6.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst6.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_2_4 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_2_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_2_4  (
            .in0(N__27627),
            .in1(N__29779),
            .in2(N__27444),
            .in3(N__27876),
            .lcout(),
            .ltout(\b2v_inst6.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIR58V1_0_LC_9_2_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIR58V1_0_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIR58V1_0_LC_9_2_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.curr_state_RNIR58V1_0_LC_9_2_5  (
            .in0(_gnd_net_),
            .in1(N__27801),
            .in2(N__27795),
            .in3(N__28383),
            .lcout(\b2v_inst6.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNICV5H1_0_LC_9_2_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNICV5H1_0_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNICV5H1_0_LC_9_2_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst6.count_RNICV5H1_0_LC_9_2_6  (
            .in0(N__33552),
            .in1(N__33529),
            .in2(_gnd_net_),
            .in3(N__33101),
            .lcout(),
            .ltout(\b2v_inst6.count_RNICV5H1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNISGKB5_0_LC_9_2_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNISGKB5_0_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNISGKB5_0_LC_9_2_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNISGKB5_0_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(N__33510),
            .in2(N__27792),
            .in3(N__33459),
            .lcout(\b2v_inst6.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIAQ3L3_LC_9_3_0 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIAQ3L3_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIAQ3L3_LC_9_3_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIAQ3L3_LC_9_3_0  (
            .in0(N__27625),
            .in1(N__27899),
            .in2(N__27888),
            .in3(N__35832),
            .lcout(),
            .ltout(\b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_LC_9_3_1 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_LC_9_3_1 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27789),
            .in3(N__29112),
            .lcout(N_222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI_0_LC_9_3_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI_0_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI_0_LC_9_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.curr_state_RNI_0_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27640),
            .lcout(\b2v_inst6.N_2992_i ),
            .ltout(\b2v_inst6.N_2992_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIKIRD1_0_0_LC_9_3_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIKIRD1_0_0_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIKIRD1_0_0_LC_9_3_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIKIRD1_0_0_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(N__27841),
            .in2(N__27738),
            .in3(N__27858),
            .lcout(\b2v_inst6.N_276_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst31.un6_output_LC_9_3_4 .C_ON=1'b0;
    defparam \b2v_inst31.un6_output_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst31.un6_output_LC_9_3_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst31.un6_output_LC_9_3_4  (
            .in0(N__27730),
            .in1(N__27705),
            .in2(N__29118),
            .in3(N__27693),
            .lcout(vccinaux_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIKIRD1_0_LC_9_3_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIKIRD1_0_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIKIRD1_0_LC_9_3_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIKIRD1_0_LC_9_3_5  (
            .in0(N__27641),
            .in1(N__27842),
            .in2(_gnd_net_),
            .in3(N__27859),
            .lcout(\b2v_inst6.curr_state_RNIKIRD1Z0Z_0 ),
            .ltout(\b2v_inst6.curr_state_RNIKIRD1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_9_3_6 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_9_3_6 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_LC_9_3_6  (
            .in0(N__27887),
            .in1(N__27900),
            .in2(N__27891),
            .in3(N__35833),
            .lcout(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36673),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNICV5H1_0_LC_9_3_7 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNICV5H1_0_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNICV5H1_0_LC_9_3_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst6.curr_state_RNICV5H1_0_LC_9_3_7  (
            .in0(N__27874),
            .in1(N__27860),
            .in2(N__28410),
            .in3(N__27843),
            .lcout(\b2v_inst6.curr_state_RNICV5H1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_LC_9_4_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_LC_9_4_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__30083),
            .in2(_gnd_net_),
            .in3(N__30283),
            .lcout(),
            .ltout(\b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI1LVK5_0_LC_9_4_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI1LVK5_0_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI1LVK5_0_LC_9_4_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI1LVK5_0_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__27816),
            .in2(N__27828),
            .in3(N__33803),
            .lcout(\b2v_inst11.count_clkZ0Z_0 ),
            .ltout(\b2v_inst11.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_1_LC_9_4_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_1_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_1_LC_9_4_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_1_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__30113),
            .in2(N__27825),
            .in3(N__30284),
            .lcout(\b2v_inst11.count_clk_RNIZ0Z_1 ),
            .ltout(\b2v_inst11.count_clk_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI2MVK5_1_LC_9_4_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI2MVK5_1_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI2MVK5_1_LC_9_4_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI2MVK5_1_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__27809),
            .in2(N__27822),
            .in3(N__33802),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_1 ),
            .ltout(\b2v_inst11.un1_count_clk_2_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_1_LC_9_4_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_1_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_1_LC_9_4_4 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \b2v_inst11.count_clk_1_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__30084),
            .in2(N__27819),
            .in3(N__30286),
            .lcout(\b2v_inst11.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36840),
            .ce(N__33808),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_0_LC_9_4_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_0_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_0_LC_9_4_5 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst11.count_clk_0_LC_9_4_5  (
            .in0(N__30285),
            .in1(_gnd_net_),
            .in2(N__30094),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36840),
            .ce(N__33808),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI2MVK5_0_1_LC_9_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI2MVK5_0_1_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI2MVK5_0_1_LC_9_4_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \b2v_inst11.count_clk_RNI2MVK5_0_1_LC_9_4_6  (
            .in0(N__27810),
            .in1(_gnd_net_),
            .in2(N__33830),
            .in3(N__27966),
            .lcout(\b2v_inst11.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVE6Q5_11_LC_9_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVE6Q5_11_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVE6Q5_11_LC_9_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_clk_RNIVE6Q5_11_LC_9_4_7  (
            .in0(N__30174),
            .in1(N__30201),
            .in2(_gnd_net_),
            .in3(N__33807),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI0TCLB_0_2_LC_9_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI0TCLB_0_2_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI0TCLB_0_2_LC_9_5_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.count_clk_RNI0TCLB_0_2_LC_9_5_0  (
            .in0(N__33639),
            .in1(N__27918),
            .in2(N__32883),
            .in3(N__32811),
            .lcout(\b2v_inst11.N_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI10NQ5_3_LC_9_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI10NQ5_3_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI10NQ5_3_LC_9_5_1 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \b2v_inst11.count_clk_RNI10NQ5_3_LC_9_5_1  (
            .in0(N__27909),
            .in1(N__30044),
            .in2(N__33831),
            .in3(N__30253),
            .lcout(\b2v_inst11.count_clkZ0Z_3 ),
            .ltout(\b2v_inst11.count_clkZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI0TCLB_2_LC_9_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI0TCLB_2_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI0TCLB_2_LC_9_5_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \b2v_inst11.count_clk_RNI0TCLB_2_LC_9_5_2  (
            .in0(N__32879),
            .in1(N__32810),
            .in2(N__27936),
            .in3(N__30521),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIG510T_7_LC_9_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIG510T_7_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIG510T_7_LC_9_5_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \b2v_inst11.count_clk_RNIG510T_7_LC_9_5_3  (
            .in0(N__33638),
            .in1(N__27933),
            .in2(N__27927),
            .in3(N__30150),
            .lcout(\b2v_inst11.count_clk_RNIG510TZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI10NQ5_2_3_LC_9_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI10NQ5_2_3_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI10NQ5_2_3_LC_9_5_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst11.count_clk_RNI10NQ5_2_3_LC_9_5_4  (
            .in0(N__27924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30522),
            .lcout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_0_LC_9_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_0_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_0_LC_9_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_0_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__30252),
            .in2(_gnd_net_),
            .in3(N__30043),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI10NQ5_0_3_LC_9_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI10NQ5_0_3_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI10NQ5_0_3_LC_9_5_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI10NQ5_0_3_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__27908),
            .in2(N__27912),
            .in3(N__33812),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_3_LC_9_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_3_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_3_LC_9_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_clk_3_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__30045),
            .in2(_gnd_net_),
            .in3(N__30254),
            .lcout(\b2v_inst11.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36862),
            .ce(N__33836),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNILIMRT_7_LC_9_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNILIMRT_7_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNILIMRT_7_LC_9_6_0 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \b2v_inst11.count_clk_RNILIMRT_7_LC_9_6_0  (
            .in0(N__39086),
            .in1(N__30644),
            .in2(N__38416),
            .in3(N__28047),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIJ9H9T_5_LC_9_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIJ9H9T_5_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIJ9H9T_5_LC_9_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNIJ9H9T_5_LC_9_6_1  (
            .in0(N__39272),
            .in1(N__28580),
            .in2(N__30768),
            .in3(N__29304),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIOM65U_1_LC_9_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIOM65U_1_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIOM65U_1_LC_9_6_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \b2v_inst11.func_state_RNIOM65U_1_LC_9_6_2  (
            .in0(N__38409),
            .in1(N__39091),
            .in2(N__28041),
            .in3(N__38848),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIIGCET1_1_LC_9_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIIGCET1_1_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIIGCET1_1_LC_9_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.func_state_RNIIGCET1_1_LC_9_6_3  (
            .in0(N__30370),
            .in1(N__28028),
            .in2(N__28038),
            .in3(N__28035),
            .lcout(\b2v_inst11.func_state_RNIIGCET1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_1_LC_9_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_9_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_1_LC_9_6_4  (
            .in0(N__39087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30753),
            .lcout(\b2v_inst11.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIAK492_0_LC_9_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIAK492_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIAK492_0_LC_9_6_5 .LUT_INIT=16'b0000111101111111;
    LogicCell40 \b2v_inst11.func_state_RNIAK492_0_LC_9_6_5  (
            .in0(N__30645),
            .in1(N__38408),
            .in2(N__39159),
            .in3(N__28029),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m2_am_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINCPR4_0_LC_9_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINCPR4_0_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINCPR4_0_LC_9_6_6 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \b2v_inst11.func_state_RNINCPR4_0_LC_9_6_6  (
            .in0(N__28705),
            .in1(N__28004),
            .in2(N__28020),
            .in3(N__30754),
            .lcout(\b2v_inst11.func_state_RNINCPR4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8BVM1_0_LC_9_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8BVM1_0_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8BVM1_0_LC_9_6_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst11.func_state_RNI8BVM1_0_LC_9_6_7  (
            .in0(N__28005),
            .in1(_gnd_net_),
            .in2(N__30769),
            .in3(N__28593),
            .lcout(\b2v_inst11.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_9_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_9_7_0 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \b2v_inst11.VCCST_EN_i_0_i_LC_9_7_0  (
            .in0(N__28113),
            .in1(N__28387),
            .in2(N__28815),
            .in3(N__38515),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_0_LC_9_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_9_7_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.func_state_RNI_0_0_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__39054),
            .in2(_gnd_net_),
            .in3(N__30634),
            .lcout(\b2v_inst11.func_state_RNI_0Z0Z_0 ),
            .ltout(\b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_9_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_9_7_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__28587),
            .in2(N__28563),
            .in3(N__28157),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_en_LC_9_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_en_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_en_LC_9_7_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \b2v_inst11.count_off_en_LC_9_7_3  (
            .in0(N__28560),
            .in1(N__35782),
            .in2(N__28554),
            .in3(N__28608),
            .lcout(\b2v_inst11.count_off_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_9_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_9_7_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_9_7_4  (
            .in0(N__38704),
            .in1(N__38516),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_7_5 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_7_5  (
            .in0(N__28144),
            .in1(N__28112),
            .in2(N__28413),
            .in3(N__28810),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_9_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_9_7_6 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_9_7_6  (
            .in0(N__39273),
            .in1(N__38517),
            .in2(N__38723),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ),
            .ltout(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_9_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_9_7_7 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_9_7_7  (
            .in0(N__28388),
            .in1(N__28114),
            .in2(N__28161),
            .in3(N__28814),
            .lcout(\b2v_inst11.N_382_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIG2BA2_0_LC_9_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIG2BA2_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIG2BA2_0_LC_9_8_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \b2v_inst11.func_state_RNIG2BA2_0_LC_9_8_0  (
            .in0(N__28740),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37641),
            .lcout(),
            .ltout(\b2v_inst11.g0_4_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIOFQO2_0_LC_9_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIOFQO2_0_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIOFQO2_0_LC_9_8_1 .LUT_INIT=16'b1111000111111011;
    LogicCell40 \b2v_inst11.func_state_RNIOFQO2_0_LC_9_8_1  (
            .in0(N__28143),
            .in1(N__28111),
            .in2(N__28050),
            .in3(N__28808),
            .lcout(\b2v_inst11.N_140_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_0_0_LC_9_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_0_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_0_0_LC_9_8_2 .LUT_INIT=16'b0001000110010001;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_0_0_LC_9_8_2  (
            .in0(N__38679),
            .in1(N__38553),
            .in2(N__30643),
            .in3(N__39287),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_7_LC_9_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_7_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_7_LC_9_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_7_LC_9_8_3  (
            .in0(N__38036),
            .in1(N__39127),
            .in2(_gnd_net_),
            .in3(N__32248),
            .lcout(\b2v_inst11.dutycycle_RNI_9Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_ss0_i_0_x2_LC_9_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_ss0_i_0_x2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_1_ss0_i_0_x2_LC_9_8_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.func_state_1_ss0_i_0_x2_LC_9_8_4  (
            .in0(N__38677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38552),
            .lcout(\b2v_inst11.N_160_i ),
            .ltout(\b2v_inst11.N_160_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI5DLR_0_LC_9_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI5DLR_0_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI5DLR_0_LC_9_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI5DLR_0_LC_9_8_5  (
            .in0(N__28631),
            .in1(N__28671),
            .in2(N__28722),
            .in3(N__30629),
            .lcout(\b2v_inst11.func_state_RNI5DLRZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI2MQD_0_LC_9_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI2MQD_0_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI2MQD_0_LC_9_8_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI2MQD_0_LC_9_8_6  (
            .in0(N__38678),
            .in1(N__30633),
            .in2(N__28679),
            .in3(N__28632),
            .lcout(\b2v_inst11.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_9_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_9_8_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_9_8_7  (
            .in0(N__34058),
            .in1(N__30430),
            .in2(N__28680),
            .in3(N__28628),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_313_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIL4TIA_1_LC_9_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIL4TIA_1_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIL4TIA_1_LC_9_9_0 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIL4TIA_1_LC_9_9_0  (
            .in0(N__28934),
            .in1(N__35790),
            .in2(N__29169),
            .in3(N__28599),
            .lcout(\b2v_inst11.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2B_LC_9_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2B_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2B_LC_9_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2B_LC_9_9_1  (
            .in0(N__31320),
            .in1(N__30561),
            .in2(_gnd_net_),
            .in3(N__35919),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2BZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNI6TFA1_LC_9_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNI6TFA1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNI6TFA1_LC_9_9_2 .LUT_INIT=16'b1110111110101011;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNI6TFA1_LC_9_9_2  (
            .in0(N__30436),
            .in1(N__39117),
            .in2(N__28602),
            .in3(N__30627),
            .lcout(\b2v_inst11.dutycycle_1_0_1 ),
            .ltout(\b2v_inst11.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_LC_9_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_1_LC_9_9_3 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \b2v_inst11.dutycycle_1_LC_9_9_3  (
            .in0(N__29162),
            .in1(N__35798),
            .in2(N__28938),
            .in3(N__28935),
            .lcout(\b2v_inst11.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36973),
            .ce(),
            .sr(N__36324));
    defparam \b2v_inst11.dutycycle_0_LC_9_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_0_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_0_LC_9_9_4 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \b2v_inst11.dutycycle_0_LC_9_9_4  (
            .in0(N__28923),
            .in1(N__29028),
            .in2(N__28917),
            .in3(N__35792),
            .lcout(\b2v_inst11.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36973),
            .ce(),
            .sr(N__36324));
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_LC_9_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_0_LC_9_9_5 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_0_LC_9_9_5  (
            .in0(N__30628),
            .in1(N__30437),
            .in2(N__31556),
            .in3(N__39128),
            .lcout(\b2v_inst11.dutycycle_1_0_0 ),
            .ltout(\b2v_inst11.dutycycle_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIR0IIA_0_LC_9_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIR0IIA_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIR0IIA_0_LC_9_9_6 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIR0IIA_0_LC_9_9_6  (
            .in0(N__28913),
            .in1(N__29027),
            .in2(N__28905),
            .in3(N__35791),
            .lcout(\b2v_inst11.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_0_LC_9_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_0_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_0_LC_9_9_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_0_LC_9_9_7  (
            .in0(N__31527),
            .in1(N__35920),
            .in2(N__31455),
            .in3(N__38274),
            .lcout(\b2v_inst11.dutycycle_RNI_8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_0_LC_9_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_0_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_1_0_LC_9_10_0 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_1_0_LC_9_10_0  (
            .in0(N__32285),
            .in1(N__36174),
            .in2(N__28872),
            .in3(N__28885),
            .lcout(),
            .ltout(\b2v_inst11.func_state_RNIDQ4A1_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIQK9K2_1_LC_9_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIQK9K2_1_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIQK9K2_1_LC_9_10_1 .LUT_INIT=16'b1110000011110001;
    LogicCell40 \b2v_inst11.func_state_RNIQK9K2_1_LC_9_10_1  (
            .in0(N__34050),
            .in1(N__28871),
            .in2(N__28830),
            .in3(N__28827),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIH3DN3_1_LC_9_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIH3DN3_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIH3DN3_1_LC_9_10_2 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \b2v_inst11.func_state_RNIH3DN3_1_LC_9_10_2  (
            .in0(N__39295),
            .in1(_gnd_net_),
            .in2(N__28821),
            .in3(N__29088),
            .lcout(\b2v_inst11.N_186_i ),
            .ltout(\b2v_inst11.N_186_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIH6AK7_2_LC_9_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIH6AK7_2_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIH6AK7_2_LC_9_10_3 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \b2v_inst11.dutycycle_RNIH6AK7_2_LC_9_10_3  (
            .in0(N__37340),
            .in1(N__29149),
            .in2(N__28818),
            .in3(N__29190),
            .lcout(\b2v_inst11.dutycycle_eena_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_9_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_9_10_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_0_LC_9_10_4  (
            .in0(N__31394),
            .in1(N__34051),
            .in2(N__31557),
            .in3(N__38846),
            .lcout(\b2v_inst11.un1_dutycycle_96_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5HTD8_1_LC_9_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5HTD8_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5HTD8_1_LC_9_10_5 .LUT_INIT=16'b0101010011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI5HTD8_1_LC_9_10_5  (
            .in0(N__29124),
            .in1(N__31393),
            .in2(N__29107),
            .in3(N__37342),
            .lcout(\b2v_inst11.dutycycle_eena_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNII85R5_1_LC_9_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNII85R5_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNII85R5_1_LC_9_10_6 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \b2v_inst11.func_state_RNII85R5_1_LC_9_10_6  (
            .in0(N__29150),
            .in1(N__29297),
            .in2(N__29108),
            .in3(N__29130),
            .lcout(\b2v_inst11.N_117_f0_1 ),
            .ltout(\b2v_inst11.N_117_f0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5HTD8_0_LC_9_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5HTD8_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5HTD8_0_LC_9_10_7 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI5HTD8_0_LC_9_10_7  (
            .in0(N__29089),
            .in1(N__31528),
            .in2(N__29031),
            .in3(N__37341),
            .lcout(\b2v_inst11.dutycycle_eena ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_9_LC_9_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_9_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_9_LC_9_11_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst11.dutycycle_9_LC_9_11_0  (
            .in0(N__35361),
            .in1(N__35345),
            .in2(N__35852),
            .in3(N__35325),
            .lcout(\b2v_inst11.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37068),
            .ce(),
            .sr(N__36325));
    defparam \b2v_inst11.dutycycle_2_LC_9_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_2_LC_9_11_1 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_2_LC_9_11_1 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \b2v_inst11.dutycycle_2_LC_9_11_1  (
            .in0(N__29019),
            .in1(N__29009),
            .in2(N__35856),
            .in3(N__28989),
            .lcout(\b2v_inst11.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37068),
            .ce(),
            .sr(N__36325));
    defparam \b2v_inst11.dutycycle_RNITBE6C_2_LC_9_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITBE6C_2_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITBE6C_2_LC_9_11_3 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNITBE6C_2_LC_9_11_3  (
            .in0(N__29018),
            .in1(N__35817),
            .in2(N__29010),
            .in3(N__28988),
            .lcout(\b2v_inst11.dutycycleZ0Z_1 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_LC_9_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_9_11_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_LC_9_11_4  (
            .in0(N__34165),
            .in1(N__28980),
            .in2(N__28968),
            .in3(N__28965),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_9_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_9_11_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_2_LC_9_11_5  (
            .in0(N__32268),
            .in1(_gnd_net_),
            .in2(N__39160),
            .in3(N__31257),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_2_LC_9_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_2_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_2_LC_9_11_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_2_LC_9_11_6  (
            .in0(N__31258),
            .in1(N__39095),
            .in2(_gnd_net_),
            .in3(N__32267),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_1_LC_9_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_9_11_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst11.func_state_RNI_1_1_LC_9_11_7  (
            .in0(N__32269),
            .in1(_gnd_net_),
            .in2(N__39161),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.func_state_RNI_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICO933_12_LC_9_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICO933_12_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICO933_12_LC_9_12_0 .LUT_INIT=16'b0101010111011111;
    LogicCell40 \b2v_inst11.dutycycle_RNICO933_12_LC_9_12_0  (
            .in0(N__37344),
            .in1(N__37704),
            .in2(N__29247),
            .in3(N__29199),
            .lcout(\b2v_inst11.dutycycle_eena_9 ),
            .ltout(\b2v_inst11.dutycycle_eena_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNII1EI5_12_LC_9_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNII1EI5_12_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNII1EI5_12_LC_9_12_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \b2v_inst11.dutycycle_RNII1EI5_12_LC_9_12_1  (
            .in0(N__35779),
            .in1(N__31088),
            .in2(N__29286),
            .in3(N__29363),
            .lcout(\b2v_inst11.dutycycleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNICO933_1_LC_9_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNICO933_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNICO933_1_LC_9_12_2 .LUT_INIT=16'b0011001101111111;
    LogicCell40 \b2v_inst11.func_state_RNICO933_1_LC_9_12_2  (
            .in0(N__29243),
            .in1(N__37343),
            .in2(N__29280),
            .in3(N__29198),
            .lcout(\b2v_inst11.dutycycle_eena_7 ),
            .ltout(\b2v_inst11.dutycycle_eena_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_11_LC_9_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_11_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_11_LC_9_12_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst11.dutycycle_11_LC_9_12_3  (
            .in0(N__29355),
            .in1(N__31598),
            .in2(N__29283),
            .in3(N__35781),
            .lcout(\b2v_inst11.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37126),
            .ce(),
            .sr(N__36326));
    defparam \b2v_inst11.dutycycle_RNI_2_12_LC_9_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_12_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_12_LC_9_12_4 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_12_LC_9_12_4  (
            .in0(N__29275),
            .in1(N__37705),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst11.N_360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5AV24_2_LC_9_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5AV24_2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5AV24_2_LC_9_12_5 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI5AV24_2_LC_9_12_5  (
            .in0(N__29242),
            .in1(N__37500),
            .in2(N__29208),
            .in3(N__29205),
            .lcout(\b2v_inst11.N_234_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_12_LC_9_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_12_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_12_LC_9_12_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \b2v_inst11.dutycycle_12_LC_9_12_6  (
            .in0(N__29364),
            .in1(N__35780),
            .in2(N__29373),
            .in3(N__31089),
            .lcout(\b2v_inst11.dutycycleZ1Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37126),
            .ce(),
            .sr(N__36326));
    defparam \b2v_inst11.dutycycle_RNIFMPT5_11_LC_9_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIFMPT5_11_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIFMPT5_11_LC_9_12_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIFMPT5_11_LC_9_12_7  (
            .in0(N__29354),
            .in1(N__31599),
            .in2(N__35831),
            .in3(N__29346),
            .lcout(\b2v_inst11.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_9_LC_9_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_9_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_9_LC_9_13_0 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_9_LC_9_13_0  (
            .in0(N__38160),
            .in1(N__35545),
            .in2(N__38351),
            .in3(N__34953),
            .lcout(\b2v_inst11.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_8_LC_9_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_8_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_8_LC_9_13_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_8_LC_9_13_1  (
            .in0(N__34955),
            .in1(N__38336),
            .in2(N__37934),
            .in3(N__35070),
            .lcout(),
            .ltout(\b2v_inst11.N_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_LC_9_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_9_13_2 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_LC_9_13_2  (
            .in0(N__29340),
            .in1(N__35370),
            .in2(N__29334),
            .in3(N__31948),
            .lcout(\b2v_inst11.un1_dutycycle_53_55_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_9_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_9_13_3 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_3_LC_9_13_3  (
            .in0(N__35544),
            .in1(_gnd_net_),
            .in2(N__34993),
            .in3(N__34355),
            .lcout(\b2v_inst11.N_355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_9_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_9_13_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_9_LC_9_13_4  (
            .in0(N__38161),
            .in1(N__34954),
            .in2(_gnd_net_),
            .in3(N__38329),
            .lcout(),
            .ltout(\b2v_inst11.g0_6_a5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_7_LC_9_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_7_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_7_LC_9_13_5 .LUT_INIT=16'b0101011101010111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_7_LC_9_13_5  (
            .in0(N__38023),
            .in1(N__29310),
            .in2(N__29313),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_9_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_9_13_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_3_LC_9_13_6  (
            .in0(N__34356),
            .in1(N__37923),
            .in2(_gnd_net_),
            .in3(N__38328),
            .lcout(\b2v_inst11.g0_6_a5_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_15_LC_9_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_9_13_7 .LUT_INIT=16'b1100110010011001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_15_LC_9_13_7  (
            .in0(N__39175),
            .in1(N__37593),
            .in2(_gnd_net_),
            .in3(N__32309),
            .lcout(\b2v_inst11.un1_dutycycle_94_axb_15_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_9_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_9_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_7_LC_9_14_0  (
            .in0(N__34982),
            .in1(N__38034),
            .in2(_gnd_net_),
            .in3(N__34382),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_11_LC_9_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_11_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_11_LC_9_14_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_11_LC_9_14_1  (
            .in0(N__39171),
            .in1(N__31970),
            .in2(_gnd_net_),
            .in3(N__32308),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_9_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_9_14_2 .LUT_INIT=16'b1010011010011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_7_LC_9_14_2  (
            .in0(N__37916),
            .in1(N__38035),
            .in2(N__35010),
            .in3(N__34383),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_LC_9_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_9_14_3 .LUT_INIT=16'b1111111110001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_LC_9_14_3  (
            .in0(N__34962),
            .in1(N__37915),
            .in2(N__35554),
            .in3(N__38136),
            .lcout(\b2v_inst11.un1_dutycycle_53_44_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_6_i_l_fx_LC_9_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_6_i_l_fx_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_6_i_l_fx_LC_9_14_5 .LUT_INIT=16'b0000000111111110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_6_i_l_fx_LC_9_14_5  (
            .in0(N__29442),
            .in1(N__29413),
            .in2(N__29481),
            .in3(N__29508),
            .lcout(\b2v_inst11.mult1_un54_sum_axb_6_i_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_5_i_l_ofx_LC_9_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_5_i_l_ofx_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_5_i_l_ofx_LC_9_14_6 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_5_i_l_ofx_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__29441),
            .in2(N__29415),
            .in3(N__29477),
            .lcout(\b2v_inst11.mult1_un54_sum_axb_5_i_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_1_axbxc3_LC_9_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_1_axbxc3_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_1_axbxc3_LC_9_14_7 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_1_axbxc3_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29447),
            .in3(N__29409),
            .lcout(\b2v_inst11.mult1_un47_sum1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_9_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_9_15_0 .LUT_INIT=16'b1110011100011000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_11_LC_9_15_0  (
            .in0(N__35466),
            .in1(N__29601),
            .in2(N__31984),
            .in3(N__31818),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_9_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_9_15_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_15_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29382),
            .in3(N__37583),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_LC_9_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_9_15_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_LC_9_15_2  (
            .in0(N__38337),
            .in1(N__34875),
            .in2(N__35490),
            .in3(N__29568),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_6 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_9_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_11_LC_9_15_3  (
            .in0(N__35199),
            .in1(N__35467),
            .in2(N__29595),
            .in3(N__31965),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_15_LC_9_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_15_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_15_LC_9_15_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_15_LC_9_15_4  (
            .in0(N__37584),
            .in1(_gnd_net_),
            .in2(N__29628),
            .in3(N__35195),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_14_LC_9_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_9_15_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_14_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35209),
            .in3(N__29627),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_9_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_9_15_7 .LUT_INIT=16'b0111000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_11_LC_9_15_7  (
            .in0(N__29567),
            .in1(N__35486),
            .in2(N__35083),
            .in3(N__31961),
            .lcout(\b2v_inst11.un1_dutycycle_53_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_9_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_9_16_0 .LUT_INIT=16'b0011001100111011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_8_LC_9_16_0  (
            .in0(N__35555),
            .in1(N__37927),
            .in2(N__29616),
            .in3(N__38162),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_9_LC_9_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_9_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_9_LC_9_16_1 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_9_LC_9_16_1  (
            .in0(N__38331),
            .in1(N__35556),
            .in2(N__38169),
            .in3(N__35007),
            .lcout(\b2v_inst11.N_35_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_9_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_9_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_10_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__35464),
            .in2(_gnd_net_),
            .in3(N__34598),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_9_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_9_16_3 .LUT_INIT=16'b0110100110100101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_9_LC_9_16_3  (
            .in0(N__38167),
            .in1(N__29559),
            .in2(N__29553),
            .in3(N__29550),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_9_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_9_16_4 .LUT_INIT=16'b0011001101110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_9_LC_9_16_4  (
            .in0(N__35008),
            .in1(N__38166),
            .in2(N__35085),
            .in3(N__38332),
            .lcout(),
            .ltout(\b2v_inst11.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_9_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_9_16_5 .LUT_INIT=16'b1111111101110101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_10_LC_9_16_5  (
            .in0(N__35465),
            .in1(N__37928),
            .in2(N__29640),
            .in3(N__29637),
            .lcout(),
            .ltout(\b2v_inst11.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_9_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_9_16_6 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_11_LC_9_16_6  (
            .in0(N__31985),
            .in1(N__34599),
            .in2(N__29631),
            .in3(N__37756),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_LC_9_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_LC_9_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_LC_9_16_7  (
            .in0(N__38330),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35006),
            .lcout(\b2v_inst11.g0_6_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNI8C4L1_LC_11_1_0 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNI8C4L1_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNI8C4L1_LC_11_1_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_c_RNI8C4L1_LC_11_1_0  (
            .in0(N__29815),
            .in1(N__29958),
            .in2(N__33230),
            .in3(N__29945),
            .lcout(\b2v_inst6.count_rst_7 ),
            .ltout(\b2v_inst6.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIV4JF5_7_LC_11_1_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIV4JF5_7_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIV4JF5_7_LC_11_1_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNIV4JF5_7_LC_11_1_1  (
            .in0(_gnd_net_),
            .in1(N__32447),
            .in2(N__29607),
            .in3(N__33408),
            .lcout(\b2v_inst6.un2_count_1_axb_7 ),
            .ltout(\b2v_inst6.un2_count_1_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_7_LC_11_1_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_7_LC_11_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_7_LC_11_1_2 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.count_7_LC_11_1_2  (
            .in0(N__29818),
            .in1(N__33198),
            .in2(N__29604),
            .in3(N__29946),
            .lcout(\b2v_inst6.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36861),
            .ce(N__33418),
            .sr(N__33196));
    defparam \b2v_inst6.count_5_LC_11_1_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_5_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_5_LC_11_1_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.count_5_LC_11_1_3  (
            .in0(N__29655),
            .in1(N__29819),
            .in2(N__32330),
            .in3(N__33195),
            .lcout(\b2v_inst6.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36861),
            .ce(N__33418),
            .sr(N__33196));
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNIJOFS1_LC_11_1_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNIJOFS1_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNIJOFS1_LC_11_1_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_c_RNIJOFS1_LC_11_1_4  (
            .in0(N__29816),
            .in1(N__32404),
            .in2(N__33231),
            .in3(N__29855),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNILTEO5_11_LC_11_1_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNILTEO5_11_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNILTEO5_11_LC_11_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNILTEO5_11_LC_11_1_5  (
            .in0(_gnd_net_),
            .in1(N__29826),
            .in2(N__29832),
            .in3(N__33409),
            .lcout(\b2v_inst6.countZ0Z_11 ),
            .ltout(\b2v_inst6.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_11_LC_11_1_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_11_LC_11_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_11_LC_11_1_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.count_11_LC_11_1_6  (
            .in0(N__29817),
            .in1(N__33197),
            .in2(N__29829),
            .in3(N__29856),
            .lcout(\b2v_inst6.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36861),
            .ce(N__33418),
            .sr(N__33196));
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNI682L1_LC_11_1_7 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNI682L1_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNI682L1_LC_11_1_7 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_c_RNI682L1_LC_11_1_7  (
            .in0(N__29654),
            .in1(N__33188),
            .in2(N__32331),
            .in3(N__29814),
            .lcout(\b2v_inst6.count_rst_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_2_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__32429),
            .in2(N__33590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNIN2P3_LC_11_2_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNIN2P3_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNIN2P3_LC_11_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_RNIN2P3_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(N__32460),
            .in2(_gnd_net_),
            .in3(N__29742),
            .lcout(\b2v_inst6.un2_count_1_cry_1_c_RNIN2PZ0Z3 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_1 ),
            .carryout(\b2v_inst6.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__29739),
            .in2(_gnd_net_),
            .in3(N__29703),
            .lcout(\b2v_inst6.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_2 ),
            .carryout(\b2v_inst6.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_2_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(N__29700),
            .in2(_gnd_net_),
            .in3(N__29658),
            .lcout(\b2v_inst6.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_3 ),
            .carryout(\b2v_inst6.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__32323),
            .in2(_gnd_net_),
            .in3(N__29646),
            .lcout(\b2v_inst6.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_4 ),
            .carryout(\b2v_inst6.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_2_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_2_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32598),
            .in3(N__29643),
            .lcout(\b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_5 ),
            .carryout(\b2v_inst6.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_6 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_6  (
            .in0(_gnd_net_),
            .in1(N__29957),
            .in2(_gnd_net_),
            .in3(N__29937),
            .lcout(\b2v_inst6.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_6 ),
            .carryout(\b2v_inst6.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_2_7 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(N__29934),
            .in2(_gnd_net_),
            .in3(N__29898),
            .lcout(\b2v_inst6.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_7 ),
            .carryout(\b2v_inst6.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_3_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__29895),
            .in2(_gnd_net_),
            .in3(N__29862),
            .lcout(\b2v_inst6.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIVI14_LC_11_3_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIVI14_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIVI14_LC_11_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst6.un2_count_1_cry_9_c_RNIVI14_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__32553),
            .in2(_gnd_net_),
            .in3(N__29859),
            .lcout(\b2v_inst6.un2_count_1_cry_9_c_RNIVIZ0Z14 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_9 ),
            .carryout(\b2v_inst6.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__32408),
            .in2(_gnd_net_),
            .in3(N__29844),
            .lcout(\b2v_inst6.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_10 ),
            .carryout(\b2v_inst6.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNI8RAB_LC_11_3_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNI8RAB_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNI8RAB_LC_11_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst6.un2_count_1_cry_11_c_RNI8RAB_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__32559),
            .in2(_gnd_net_),
            .in3(N__29841),
            .lcout(\b2v_inst6.un2_count_1_cry_11_c_RNI8RABZ0 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_11 ),
            .carryout(\b2v_inst6.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNI9TBB_LC_11_3_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNI9TBB_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNI9TBB_LC_11_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst6.un2_count_1_cry_12_c_RNI9TBB_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__30009),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(\b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_12 ),
            .carryout(\b2v_inst6.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNIR6IO5_LC_11_3_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNIR6IO5_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNIR6IO5_LC_11_3_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_13_c_RNIR6IO5_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32514),
            .in3(N__29835),
            .lcout(\b2v_inst6.un2_count_1_cry_13_c_RNIR6IOZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_13 ),
            .carryout(\b2v_inst6.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNIN0KS1_LC_11_3_6 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNIN0KS1_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNIN0KS1_LC_11_3_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_14_c_RNIN0KS1_LC_11_3_6  (
            .in0(N__33163),
            .in1(_gnd_net_),
            .in2(N__32775),
            .in3(N__30012),
            .lcout(\b2v_inst6.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIP3HO5_13_LC_11_3_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIP3HO5_13_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIP3HO5_13_LC_11_3_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \b2v_inst6.count_RNIP3HO5_13_LC_11_3_7  (
            .in0(N__32734),
            .in1(N__33162),
            .in2(N__32766),
            .in3(N__33410),
            .lcout(\b2v_inst6.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI1I7Q5_0_12_LC_11_4_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI1I7Q5_0_12_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI1I7Q5_0_12_LC_11_4_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \b2v_inst11.count_clk_RNI1I7Q5_0_12_LC_11_4_0  (
            .in0(N__30682),
            .in1(N__32688),
            .in2(N__32709),
            .in3(N__30792),
            .lcout(\b2v_inst11.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIM2RL5_0_10_LC_11_4_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIM2RL5_0_10_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIM2RL5_0_10_LC_11_4_1 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \b2v_inst11.count_clk_RNIM2RL5_0_10_LC_11_4_1  (
            .in0(N__30126),
            .in1(N__30339),
            .in2(N__30801),
            .in3(N__30683),
            .lcout(\b2v_inst11.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVE6Q5_0_11_LC_11_4_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVE6Q5_0_11_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVE6Q5_0_11_LC_11_4_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \b2v_inst11.count_clk_RNIVE6Q5_0_11_LC_11_4_2  (
            .in0(N__30173),
            .in1(N__30200),
            .in2(N__30687),
            .in3(N__30799),
            .lcout(\b2v_inst11.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI3L8Q5_0_13_LC_11_4_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI3L8Q5_0_13_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI3L8Q5_0_13_LC_11_4_3 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI3L8Q5_0_13_LC_11_4_3  (
            .in0(N__32670),
            .in1(N__32651),
            .in2(N__30800),
            .in3(N__30681),
            .lcout(),
            .ltout(\b2v_inst11.count_clkZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIPOH4N_10_LC_11_4_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIPOH4N_10_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIPOH4N_10_LC_11_4_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNIPOH4N_10_LC_11_4_4  (
            .in0(N__30003),
            .in1(N__29997),
            .in2(N__29991),
            .in3(N__29988),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_o2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIPOH4N_0_10_LC_11_4_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIPOH4N_0_10_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIPOH4N_0_10_LC_11_4_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNIPOH4N_0_10_LC_11_4_5  (
            .in0(N__33909),
            .in1(N__30095),
            .in2(N__29982),
            .in3(N__30846),
            .lcout(\b2v_inst11.N_175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_10_LC_11_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_10_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_10_LC_11_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_10_LC_11_4_6  (
            .in0(N__30338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37087),
            .ce(N__33797),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIM2RL5_10_LC_11_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIM2RL5_10_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIM2RL5_10_LC_11_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst11.count_clk_RNIM2RL5_10_LC_11_4_7  (
            .in0(N__30125),
            .in1(N__30337),
            .in2(_gnd_net_),
            .in3(N__33796),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_11_5_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_11_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__30117),
            .in2(N__30099),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_11_5_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_11_5_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_11_5_1  (
            .in0(N__30289),
            .in1(_gnd_net_),
            .in2(N__32841),
            .in3(N__30060),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_11_5_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_11_5_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30057),
            .in3(N__30030),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_11_5_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_11_5_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_11_5_3  (
            .in0(N__30287),
            .in1(_gnd_net_),
            .in2(N__32873),
            .in3(N__30027),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_11_5_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_11_5_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_11_5_4  (
            .in0(N__30296),
            .in1(N__32973),
            .in2(_gnd_net_),
            .in3(N__30024),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_11_5_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_11_5_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_11_5_5  (
            .in0(N__30290),
            .in1(_gnd_net_),
            .in2(N__33631),
            .in3(N__30021),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_11_5_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_11_5_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_11_5_6  (
            .in0(N__30297),
            .in1(_gnd_net_),
            .in2(N__32892),
            .in3(N__30018),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_11_5_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_11_5_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_11_5_7  (
            .in0(N__30288),
            .in1(N__30520),
            .in2(_gnd_net_),
            .in3(N__30015),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_11_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_11_6_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_11_6_0  (
            .in0(N__30264),
            .in1(N__30470),
            .in2(_gnd_net_),
            .in3(N__30351),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_11_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_11_6_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_11_6_1  (
            .in0(N__30279),
            .in1(N__30348),
            .in2(_gnd_net_),
            .in3(N__30324),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_11_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_11_6_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_11_6_2  (
            .in0(N__30265),
            .in1(N__30321),
            .in2(_gnd_net_),
            .in3(N__30309),
            .lcout(\b2v_inst11.count_clk_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_11_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_11_6_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_11_6_3  (
            .in0(N__30280),
            .in1(N__32715),
            .in2(_gnd_net_),
            .in3(N__30306),
            .lcout(\b2v_inst11.count_clk_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_11_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_11_6_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_11_6_4  (
            .in0(N__30266),
            .in1(N__32676),
            .in2(_gnd_net_),
            .in3(N__30303),
            .lcout(\b2v_inst11.count_clk_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_11_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_11_6_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_11_6_5  (
            .in0(N__30281),
            .in1(N__30845),
            .in2(_gnd_net_),
            .in3(N__30300),
            .lcout(\b2v_inst11.count_clk_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_11_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_11_6_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_11_6_6  (
            .in0(N__33905),
            .in1(N__30282),
            .in2(_gnd_net_),
            .in3(N__30204),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_11_LC_11_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_11_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_11_LC_11_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_11_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30199),
            .lcout(\b2v_inst11.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37034),
            .ce(N__33756),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI9CRQ5_0_7_LC_11_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI9CRQ5_0_7_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI9CRQ5_0_7_LC_11_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI9CRQ5_0_7_LC_11_7_0  (
            .in0(N__32924),
            .in1(N__33731),
            .in2(_gnd_net_),
            .in3(N__32909),
            .lcout(\b2v_inst11.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_7_LC_11_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_7_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_7_LC_11_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_7_LC_11_7_1  (
            .in0(N__32910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36967),
            .ce(N__33835),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIBFSQ5_8_LC_11_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIBFSQ5_8_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIBFSQ5_8_LC_11_7_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNIBFSQ5_8_LC_11_7_2  (
            .in0(N__30486),
            .in1(N__33730),
            .in2(_gnd_net_),
            .in3(N__30497),
            .lcout(\b2v_inst11.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_8_LC_11_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_8_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_8_LC_11_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_8_LC_11_7_3  (
            .in0(N__30498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36967),
            .ce(N__33835),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIDITQ5_9_LC_11_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIDITQ5_9_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIDITQ5_9_LC_11_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNIDITQ5_9_LC_11_7_4  (
            .in0(N__30447),
            .in1(N__33732),
            .in2(_gnd_net_),
            .in3(N__30455),
            .lcout(\b2v_inst11.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_9_LC_11_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_9_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_9_LC_11_7_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_9_LC_11_7_5  (
            .in0(N__30456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36967),
            .ce(N__33835),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_4_LC_11_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_4_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_4_LC_11_7_6 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_4_LC_11_7_6  (
            .in0(N__32147),
            .in1(N__39132),
            .in2(_gnd_net_),
            .in3(N__35027),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_4_LC_11_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_4_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_4_LC_11_7_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_4_LC_11_7_7  (
            .in0(N__35028),
            .in1(_gnd_net_),
            .in2(N__39176),
            .in3(N__32146),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_11_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_11_8_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__30439),
            .in2(_gnd_net_),
            .in3(N__32163),
            .lcout(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0 ),
            .ltout(\b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI0O4B5_1_LC_11_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI0O4B5_1_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI0O4B5_1_LC_11_8_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \b2v_inst11.func_state_RNI0O4B5_1_LC_11_8_1  (
            .in0(N__30699),
            .in1(N__30782),
            .in2(N__30381),
            .in3(N__30378),
            .lcout(\b2v_inst11.count_clk_en ),
            .ltout(\b2v_inst11.count_clk_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI5O9Q5_14_LC_11_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI5O9Q5_14_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI5O9Q5_14_LC_11_8_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst11.count_clk_RNI5O9Q5_14_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__30651),
            .in2(N__30849),
            .in3(N__30662),
            .lcout(\b2v_inst11.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNID7Q51_0_LC_11_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNID7Q51_0_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNID7Q51_0_LC_11_8_3 .LUT_INIT=16'b0111000000010000;
    LogicCell40 \b2v_inst11.func_state_RNID7Q51_0_LC_11_8_3  (
            .in0(N__30636),
            .in1(N__39158),
            .in2(N__30828),
            .in3(N__30770),
            .lcout(\b2v_inst11.func_state_RNID7Q51Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIJGA54_1_LC_11_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIJGA54_1_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIJGA54_1_LC_11_8_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \b2v_inst11.func_state_RNIJGA54_1_LC_11_8_4  (
            .in0(N__30771),
            .in1(N__30705),
            .in2(N__39184),
            .in3(N__30698),
            .lcout(\b2v_inst11.func_state_RNIJGA54Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_14_LC_11_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_14_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_14_LC_11_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_14_LC_11_8_5  (
            .in0(N__30663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37099),
            .ce(N__33801),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_0_LC_11_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_11_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNI_1_0_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30635),
            .lcout(\b2v_inst11.N_2904_i ),
            .ltout(\b2v_inst11.N_2904_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_11_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_11_8_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_1_LC_11_8_7  (
            .in0(N__31456),
            .in1(_gnd_net_),
            .in2(N__30579),
            .in3(N__39154),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_LC_11_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__31558),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_RNID26_LC_11_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_RNID26_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_RNID26_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_RNID26_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__30576),
            .in2(N__31440),
            .in3(N__30552),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_1 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_0_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s1_c_RNIE7GA_LC_11_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s1_c_RNIE7GA_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s1_c_RNIE7GA_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_s1_c_RNIE7GA_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__31298),
            .in2(N__30549),
            .in3(N__30987),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_1_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s1_c_RNIFCQ4_LC_11_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s1_c_RNIFCQ4_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s1_c_RNIFCQ4_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_s1_c_RNIFCQ4_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__31110),
            .in2(N__34323),
            .in3(N__30984),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_2_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s1_c_RNIGH4F_LC_11_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s1_c_RNIGH4F_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s1_c_RNIGH4F_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_3_s1_c_RNIGH4F_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__35025),
            .in2(N__30981),
            .in3(N__30954),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_3_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s1_c_RNIHME9_LC_11_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s1_c_RNIHME9_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s1_c_RNIHME9_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_s1_c_RNIHME9_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__30951),
            .in2(N__32985),
            .in3(N__30903),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_4_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s1_c_RNIIRO3_LC_11_9_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s1_c_RNIIRO3_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s1_c_RNIIRO3_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_s1_c_RNIIRO3_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__38227),
            .in2(N__31029),
            .in3(N__30900),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_5_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s1_c_RNIJ03E_LC_11_9_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s1_c_RNIJ03E_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s1_c_RNIJ03E_LC_11_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_s1_c_RNIJ03E_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__38032),
            .in2(N__30897),
            .in3(N__30882),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_7 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_6_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s1_c_RNIK5D8_LC_11_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s1_c_RNIK5D8_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s1_c_RNIK5D8_LC_11_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_7_s1_c_RNIK5D8_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__37911),
            .in2(N__30996),
            .in3(N__30879),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_8 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s1_c_RNILAN2_LC_11_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s1_c_RNILAN2_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s1_c_RNILAN2_LC_11_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_8_s1_c_RNILAN2_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__38158),
            .in2(N__30876),
            .in3(N__30864),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_9 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_8_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s1_c_RNIMF1D_LC_11_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s1_c_RNIMF1D_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s1_c_RNIMF1D_LC_11_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_9_s1_c_RNIMF1D_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__30861),
            .in2(N__35462),
            .in3(N__30852),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_9_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s1_c_RNIU1R8_LC_11_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s1_c_RNIU1R8_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s1_c_RNIU1R8_LC_11_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_10_s1_c_RNIU1R8_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__31983),
            .in2(N__31017),
            .in3(N__31074),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_10_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s1_c_RNIV653_LC_11_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s1_c_RNIV653_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s1_c_RNIV653_LC_11_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_11_s1_c_RNIV653_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__37767),
            .in2(N__32055),
            .in3(N__31071),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_11_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s1_c_RNI0CFD_LC_11_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s1_c_RNI0CFD_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s1_c_RNI0CFD_LC_11_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_12_s1_c_RNI0CFD_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__34606),
            .in2(N__31068),
            .in3(N__31053),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_12_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s1_c_RNI1HP7_LC_11_10_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s1_c_RNI1HP7_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s1_c_RNI1HP7_LC_11_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_13_s1_c_RNI1HP7_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__35204),
            .in2(N__31050),
            .in3(N__31035),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_13_s1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_s1_c_RNI2M32_LC_11_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_s1_c_RNI2M32_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_s1_c_RNI2M32_LC_11_10_7 .LUT_INIT=16'b0011011011001001;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_14_s1_c_RNI2M32_LC_11_10_7  (
            .in0(N__39084),
            .in1(N__37596),
            .in2(N__32278),
            .in3(N__31032),
            .lcout(\b2v_inst11.un1_dutycycle_94_s1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_11_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_11_11_0 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_6_LC_11_11_0  (
            .in0(N__38257),
            .in1(_gnd_net_),
            .in2(N__32273),
            .in3(N__39168),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_11_LC_11_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_11_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_11_LC_11_11_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_11_LC_11_11_1  (
            .in0(N__39170),
            .in1(N__31986),
            .in2(_gnd_net_),
            .in3(N__32204),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJ9_LC_11_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJ9_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJ9_LC_11_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJ9_LC_11_11_2  (
            .in0(N__31005),
            .in1(N__31152),
            .in2(_gnd_net_),
            .in3(N__36009),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_11_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_11_11_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_8_LC_11_11_3  (
            .in0(N__39169),
            .in1(_gnd_net_),
            .in2(N__37929),
            .in3(N__32203),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_12_LC_11_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_12_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_12_LC_11_11_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_12_LC_11_11_4  (
            .in0(N__32199),
            .in1(N__37768),
            .in2(_gnd_net_),
            .in3(N__39167),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_11_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_11_11_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_6_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__38258),
            .in2(N__39185),
            .in3(N__32196),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_11_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_11_11_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_9_LC_11_11_6  (
            .in0(N__32198),
            .in1(N__38154),
            .in2(_gnd_net_),
            .in3(N__39166),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_11_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_11_11_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_3_LC_11_11_7  (
            .in0(N__39165),
            .in1(_gnd_net_),
            .in2(N__34379),
            .in3(N__32197),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_7_LC_11_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_7_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_7_LC_11_12_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_7_LC_11_12_0  (
            .in0(N__32182),
            .in1(_gnd_net_),
            .in2(N__38033),
            .in3(N__39139),
            .lcout(\b2v_inst11.dutycycle_RNI_10Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_11_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_11_12_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_3_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__34354),
            .in2(N__39178),
            .in3(N__32181),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_14_LC_11_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_14_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_14_LC_11_12_2 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_14_LC_11_12_2  (
            .in0(N__32185),
            .in1(N__39146),
            .in2(_gnd_net_),
            .in3(N__35189),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_10_LC_11_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_10_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_10_LC_11_12_3 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_10_LC_11_12_3  (
            .in0(N__35434),
            .in1(_gnd_net_),
            .in2(N__39179),
            .in3(N__32183),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EG1_LC_11_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EG1_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EG1_LC_11_12_4 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EG1_LC_11_12_4  (
            .in0(N__36211),
            .in1(N__36004),
            .in2(N__31101),
            .in3(N__31638),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EGZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_13_LC_11_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_13_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_13_LC_11_12_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_13_LC_11_12_5  (
            .in0(N__34563),
            .in1(_gnd_net_),
            .in2(N__39180),
            .in3(N__32184),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNI8SPR1_LC_11_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNI8SPR1_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNI8SPR1_LC_11_12_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNI8SPR1_LC_11_12_6  (
            .in0(N__36049),
            .in1(N__31608),
            .in2(N__36230),
            .in3(N__31659),
            .lcout(\b2v_inst11.dutycycle_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_LC_11_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_LC_11_12_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \b2v_inst11.func_state_RNI_1_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39177),
            .in3(N__32180),
            .lcout(\b2v_inst11.N_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_LC_11_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__31584),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIC05_LC_11_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIC05_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIC05_LC_11_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIC05_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__31464),
            .in2(N__31332),
            .in3(N__31305),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_1 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_0_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNID5FA_LC_11_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNID5FA_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNID5FA_LC_11_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNID5FA_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__31300),
            .in2(N__31194),
            .in3(N__31164),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_1_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNIEAP4_LC_11_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNIEAP4_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNIEAP4_LC_11_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNIEAP4_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__34378),
            .in2(N__31161),
            .in3(N__31143),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_2_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIFF3F_LC_11_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIFF3F_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIFF3F_LC_11_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIFF3F_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__35011),
            .in2(N__31140),
            .in3(N__31116),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_3_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIGKD9_LC_11_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIGKD9_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIGKD9_LC_11_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIGKD9_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34209),
            .in3(N__31113),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_4_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIHPN3_LC_11_13_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIHPN3_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIHPN3_LC_11_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIHPN3_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__38295),
            .in2(N__31734),
            .in3(N__31722),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_5_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNIIU1E_LC_11_13_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNIIU1E_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNIIU1E_LC_11_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNIIU1E_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__31719),
            .in2(N__38022),
            .in3(N__31713),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_7 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_6_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIJ3C8_LC_11_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIJ3C8_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIJ3C8_LC_11_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIJ3C8_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__31710),
            .in2(N__37875),
            .in3(N__31698),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_8 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIK8M2_LC_11_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIK8M2_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIK8M2_LC_11_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIK8M2_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__31695),
            .in2(N__38135),
            .in3(N__31686),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_9 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_8_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNILD0D_LC_11_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNILD0D_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNILD0D_LC_11_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNILD0D_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__31683),
            .in2(N__35435),
            .in3(N__31674),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_9_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNITVP8_LC_11_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNITVP8_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNITVP8_LC_11_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNITVP8_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__31671),
            .in2(N__31989),
            .in3(N__31650),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_10_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIU443_LC_11_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIU443_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIU443_LC_11_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIU443_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__31647),
            .in2(N__37769),
            .in3(N__31629),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_11_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIV9ED_LC_11_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIV9ED_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIV9ED_LC_11_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIV9ED_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__34567),
            .in2(N__31626),
            .in3(N__31611),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_12_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI0FO7_LC_11_14_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI0FO7_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI0FO7_LC_11_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI0FO7_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__35188),
            .in2(N__31857),
            .in3(N__31845),
            .lcout(\b2v_inst11.un1_dutycycle_94_s0_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_13_s0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3A64_LC_11_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3A64_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3A64_LC_11_14_7 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3A64_LC_11_14_7  (
            .in0(N__31842),
            .in1(N__31830),
            .in2(N__36068),
            .in3(N__31821),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3AZ0Z64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_11_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_11_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_15_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__37540),
            .in2(_gnd_net_),
            .in3(N__37762),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_11_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_11_15_1 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_6_LC_11_15_1  (
            .in0(N__38342),
            .in1(N__34874),
            .in2(N__31809),
            .in3(N__35069),
            .lcout(\b2v_inst11.un1_dutycycle_53_31 ),
            .ltout(\b2v_inst11.un1_dutycycle_53_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_11_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_11_15_2 .LUT_INIT=16'b0000001111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_13_LC_11_15_2  (
            .in0(N__34569),
            .in1(N__31779),
            .in2(N__31797),
            .in3(N__37764),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_11_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_11_15_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_13_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35194),
            .in3(N__34568),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_14_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_11_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_11_15_4 .LUT_INIT=16'b0001111011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_12_LC_11_15_4  (
            .in0(N__31785),
            .in1(N__31778),
            .in2(N__31764),
            .in3(N__37763),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_11_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_11_15_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_14_LC_11_15_5  (
            .in0(N__35169),
            .in1(_gnd_net_),
            .in2(N__31761),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_11_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_11_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_9_LC_11_15_6  (
            .in0(N__38309),
            .in1(N__38123),
            .in2(N__36069),
            .in3(N__32040),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_12_LC_11_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_12_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_12_LC_11_15_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_12_LC_11_15_7  (
            .in0(N__37765),
            .in1(N__39186),
            .in2(_gnd_net_),
            .in3(N__32306),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_LC_11_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_11_16_0 .LUT_INIT=16'b1111100011100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_LC_11_16_0  (
            .in0(N__34368),
            .in1(N__38027),
            .in2(N__35026),
            .in3(N__37871),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_7 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_LC_11_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_LC_11_16_1 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_LC_11_16_1  (
            .in0(N__38340),
            .in1(_gnd_net_),
            .in2(N__32034),
            .in3(N__38131),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_10_LC_11_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_10_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_10_LC_11_16_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_10_LC_11_16_2  (
            .in0(N__35463),
            .in1(_gnd_net_),
            .in2(N__32031),
            .in3(N__31883),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIF1_LC_11_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIF1_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIF1_LC_11_16_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIF1_LC_11_16_3  (
            .in0(N__36224),
            .in1(N__32013),
            .in2(N__36059),
            .in3(N__32001),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_11_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_11_16_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_7_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__38028),
            .in2(_gnd_net_),
            .in3(N__38338),
            .lcout(\b2v_inst11.un1_i2_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_7_LC_11_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_7_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_7_LC_11_16_5 .LUT_INIT=16'b0001110000111000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_7_LC_11_16_5  (
            .in0(N__37870),
            .in1(N__35016),
            .in2(N__38037),
            .in3(N__34369),
            .lcout(),
            .ltout(\b2v_inst11.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_11_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_11_16_6 .LUT_INIT=16'b0111001011100100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_7_LC_11_16_6  (
            .in0(N__38130),
            .in1(N__38029),
            .in2(N__31992),
            .in3(N__38339),
            .lcout(\b2v_inst11.un1_N_5 ),
            .ltout(\b2v_inst11.un1_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_11_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_11_16_7 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_11_LC_11_16_7  (
            .in0(N__37872),
            .in1(N__31988),
            .in2(N__31887),
            .in3(N__31884),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRUGF5_0_5_LC_12_1_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRUGF5_0_5_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRUGF5_0_5_LC_12_1_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst6.count_RNIRUGF5_0_5_LC_12_1_0  (
            .in0(N__32340),
            .in1(_gnd_net_),
            .in2(N__33443),
            .in3(N__32349),
            .lcout(),
            .ltout(\b2v_inst6.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIQ34VA_7_LC_12_1_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIQ34VA_7_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIQ34VA_7_LC_12_1_1 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \b2v_inst6.count_RNIQ34VA_7_LC_12_1_1  (
            .in0(N__32454),
            .in1(N__32448),
            .in2(N__32436),
            .in3(N__33379),
            .lcout(\b2v_inst6.count_1_i_a3_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNICV5H1_1_LC_12_1_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNICV5H1_1_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNICV5H1_1_LC_12_1_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.count_RNICV5H1_1_LC_12_1_2  (
            .in0(N__33186),
            .in1(N__32430),
            .in2(_gnd_net_),
            .in3(N__33588),
            .lcout(\b2v_inst6.count_RNICV5H1Z0Z_1 ),
            .ltout(\b2v_inst6.count_RNICV5H1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNITHKB5_1_LC_12_1_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITHKB5_1_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITHKB5_1_LC_12_1_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNITHKB5_1_LC_12_1_3  (
            .in0(_gnd_net_),
            .in1(N__32384),
            .in2(N__32433),
            .in3(N__33377),
            .lcout(\b2v_inst6.un2_count_1_axb_1 ),
            .ltout(\b2v_inst6.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_1_LC_12_1_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_1_LC_12_1_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_1_LC_12_1_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst6.count_1_LC_12_1_4  (
            .in0(N__33187),
            .in1(_gnd_net_),
            .in2(N__32418),
            .in3(N__33589),
            .lcout(\b2v_inst6.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36968),
            .ce(N__33417),
            .sr(N__33240));
    defparam \b2v_inst6.count_RNITHKB5_0_1_LC_12_1_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITHKB5_0_1_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITHKB5_0_1_LC_12_1_5 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \b2v_inst6.count_RNITHKB5_0_1_LC_12_1_5  (
            .in0(N__32415),
            .in1(N__33383),
            .in2(N__32409),
            .in3(N__32385),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIBT0961_1_LC_12_1_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIBT0961_1_LC_12_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIBT0961_1_LC_12_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNIBT0961_1_LC_12_1_6  (
            .in0(N__32376),
            .in1(N__32367),
            .in2(N__32358),
            .in3(N__32355),
            .lcout(\b2v_inst6.count_1_i_a3_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRUGF5_5_LC_12_1_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRUGF5_5_LC_12_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRUGF5_5_LC_12_1_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIRUGF5_5_LC_12_1_7  (
            .in0(N__32348),
            .in1(N__32339),
            .in2(_gnd_net_),
            .in3(N__33378),
            .lcout(\b2v_inst6.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_2_LC_12_2_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_2_LC_12_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_2_LC_12_2_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst6.count_2_LC_12_2_0  (
            .in0(N__33204),
            .in1(N__32470),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36899),
            .ce(N__33385),
            .sr(N__33222));
    defparam \b2v_inst6.count_RNIH75D5_0_14_LC_12_2_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIH75D5_0_14_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIH75D5_0_14_LC_12_2_1 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst6.count_RNIH75D5_0_14_LC_12_2_1  (
            .in0(N__32535),
            .in1(N__32526),
            .in2(N__33455),
            .in3(N__33223),
            .lcout(\b2v_inst6.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_14_LC_12_2_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_14_LC_12_2_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_14_LC_12_2_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst6.count_14_LC_12_2_2  (
            .in0(N__32525),
            .in1(_gnd_net_),
            .in2(N__33235),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36899),
            .ce(N__33385),
            .sr(N__33222));
    defparam \b2v_inst6.count_RNIH75D5_14_LC_12_2_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIH75D5_14_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIH75D5_14_LC_12_2_3 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst6.count_RNIH75D5_14_LC_12_2_3  (
            .in0(N__32534),
            .in1(N__32524),
            .in2(N__33454),
            .in3(N__33203),
            .lcout(\b2v_inst6.un2_count_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNI32VK1_LC_12_2_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNI32VK1_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNI32VK1_LC_12_2_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_RNI32VK1_LC_12_2_4  (
            .in0(N__33208),
            .in1(N__32474),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI6TISA_2_LC_12_2_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI6TISA_2_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI6TISA_2_LC_12_2_5 .LUT_INIT=16'b0000001100010001;
    LogicCell40 \b2v_inst6.count_RNI6TISA_2_LC_12_2_5  (
            .in0(N__32484),
            .in1(N__32505),
            .in2(N__32499),
            .in3(N__33386),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIANDN72_2_LC_12_2_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIANDN72_2_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIANDN72_2_LC_12_2_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNIANDN72_2_LC_12_2_6  (
            .in0(N__32634),
            .in1(N__32496),
            .in2(N__32487),
            .in3(N__32748),
            .lcout(\b2v_inst6.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNILLDF5_2_LC_12_2_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNILLDF5_2_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNILLDF5_2_LC_12_2_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst6.count_RNILLDF5_2_LC_12_2_7  (
            .in0(N__32483),
            .in1(N__33202),
            .in2(N__32475),
            .in3(N__33384),
            .lcout(\b2v_inst6.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIT1IF5_0_6_LC_12_3_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIT1IF5_0_6_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIT1IF5_0_6_LC_12_3_0 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst6.count_RNIT1IF5_0_6_LC_12_3_0  (
            .in0(N__32628),
            .in1(N__32619),
            .in2(N__33465),
            .in3(N__33157),
            .lcout(),
            .ltout(\b2v_inst6.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI9OO0B_10_LC_12_3_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI9OO0B_10_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI9OO0B_10_LC_12_3_1 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \b2v_inst6.count_RNI9OO0B_10_LC_12_3_1  (
            .in0(N__32547),
            .in1(N__32781),
            .in2(N__32640),
            .in3(N__33446),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI0P8PG_12_LC_12_3_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI0P8PG_12_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI0P8PG_12_LC_12_3_2 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \b2v_inst6.count_RNI0P8PG_12_LC_12_3_2  (
            .in0(N__33445),
            .in1(N__32589),
            .in2(N__32637),
            .in3(N__32582),
            .lcout(\b2v_inst6.count_1_i_a3_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_6_LC_12_3_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_6_LC_12_3_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_6_LC_12_3_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst6.count_6_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__32611),
            .in2(_gnd_net_),
            .in3(N__33159),
            .lcout(\b2v_inst6.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36830),
            .ce(N__33444),
            .sr(N__33160));
    defparam \b2v_inst6.count_RNIT1IF5_6_LC_12_3_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIT1IF5_6_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIT1IF5_6_LC_12_3_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst6.count_RNIT1IF5_6_LC_12_3_4  (
            .in0(N__32627),
            .in1(N__33155),
            .in2(N__32618),
            .in3(N__33387),
            .lcout(\b2v_inst6.un2_count_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIKQGS1_LC_12_3_5 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIKQGS1_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIKQGS1_LC_12_3_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_11_c_RNIKQGS1_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__33161),
            .in2(_gnd_net_),
            .in3(N__32571),
            .lcout(\b2v_inst6.count_rst_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_12_LC_12_3_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_12_LC_12_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_12_LC_12_3_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst6.count_12_LC_12_3_6  (
            .in0(N__32570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33156),
            .lcout(\b2v_inst6.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36830),
            .ce(N__33444),
            .sr(N__33160));
    defparam \b2v_inst6.count_RNIN0GO5_12_LC_12_3_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIN0GO5_12_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIN0GO5_12_LC_12_3_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \b2v_inst6.count_RNIN0GO5_12_LC_12_3_7  (
            .in0(N__33388),
            .in1(N__33158),
            .in2(N__32583),
            .in3(N__32569),
            .lcout(\b2v_inst6.un2_count_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNICM6H5_10_LC_12_4_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNICM6H5_10_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNICM6H5_10_LC_12_4_0 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \b2v_inst6.count_RNICM6H5_10_LC_12_4_0  (
            .in0(N__33341),
            .in1(N__32546),
            .in2(N__32796),
            .in3(N__33217),
            .lcout(\b2v_inst6.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_10_LC_12_4_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_10_LC_12_4_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_10_LC_12_4_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst6.count_10_LC_12_4_1  (
            .in0(N__33218),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32791),
            .lcout(\b2v_inst6.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36890),
            .ce(N__33457),
            .sr(N__33216));
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIBI7L1_LC_12_4_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIBI7L1_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIBI7L1_LC_12_4_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_9_c_RNIBI7L1_LC_12_4_2  (
            .in0(N__32795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33221),
            .lcout(\b2v_inst6.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_13_LC_12_4_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_13_LC_12_4_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_13_LC_12_4_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst6.count_13_LC_12_4_3  (
            .in0(N__33219),
            .in1(_gnd_net_),
            .in2(N__32739),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36890),
            .ce(N__33457),
            .sr(N__33216));
    defparam \b2v_inst6.count_RNIT9JO5_15_LC_12_4_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIT9JO5_15_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIT9JO5_15_LC_12_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst6.count_RNIT9JO5_15_LC_12_4_4  (
            .in0(N__33458),
            .in1(N__33474),
            .in2(_gnd_net_),
            .in3(N__33488),
            .lcout(\b2v_inst6.countZ0Z_15 ),
            .ltout(\b2v_inst6.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIP3HO5_0_13_LC_12_4_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIP3HO5_0_13_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIP3HO5_0_13_LC_12_4_5 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \b2v_inst6.count_RNIP3HO5_0_13_LC_12_4_5  (
            .in0(N__32721),
            .in1(N__32762),
            .in2(N__32751),
            .in3(N__33340),
            .lcout(\b2v_inst6.count_1_i_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNILSHS1_LC_12_4_6 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNILSHS1_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNILSHS1_LC_12_4_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_12_c_RNILSHS1_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(N__32738),
            .in2(_gnd_net_),
            .in3(N__33220),
            .lcout(\b2v_inst6.count_rst_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI1I7Q5_12_LC_12_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI1I7Q5_12_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI1I7Q5_12_LC_12_5_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \b2v_inst11.count_clk_RNI1I7Q5_12_LC_12_5_0  (
            .in0(N__32687),
            .in1(N__32701),
            .in2(N__33825),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_12_LC_12_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_12_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_12_LC_12_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_12_LC_12_5_1  (
            .in0(N__32702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37067),
            .ce(N__33822),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI3L8Q5_13_LC_12_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI3L8Q5_13_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI3L8Q5_13_LC_12_5_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \b2v_inst11.count_clk_RNI3L8Q5_13_LC_12_5_2  (
            .in0(N__32665),
            .in1(N__32652),
            .in2(N__33826),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_13_LC_12_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_13_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_13_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_13_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32666),
            .lcout(\b2v_inst11.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37067),
            .ce(N__33822),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI56PQ5_5_LC_12_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI56PQ5_5_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI56PQ5_5_LC_12_5_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst11.count_clk_RNI56PQ5_5_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__32966),
            .in2(N__33823),
            .in3(N__32956),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_5_LC_12_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_5_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_5_LC_12_5_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_5_LC_12_5_5  (
            .in0(N__32958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37067),
            .ce(N__33822),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI56PQ5_0_5_LC_12_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI56PQ5_0_5_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI56PQ5_0_5_LC_12_5_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst11.count_clk_RNI56PQ5_0_5_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__32967),
            .in2(N__33824),
            .in3(N__32957),
            .lcout(\b2v_inst11.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI9CRQ5_7_LC_12_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI9CRQ5_7_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI9CRQ5_7_LC_12_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI9CRQ5_7_LC_12_5_7  (
            .in0(N__32928),
            .in1(N__33786),
            .in2(_gnd_net_),
            .in3(N__32903),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI33OQ5_4_LC_12_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI33OQ5_4_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI33OQ5_4_LC_12_6_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \b2v_inst11.count_clk_RNI33OQ5_4_LC_12_6_0  (
            .in0(N__32847),
            .in1(_gnd_net_),
            .in2(N__33810),
            .in3(N__32855),
            .lcout(\b2v_inst11.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_4_LC_12_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_4_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_4_LC_12_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_4_LC_12_6_1  (
            .in0(N__32856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37006),
            .ce(N__33767),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVSLQ5_2_LC_12_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVSLQ5_2_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVSLQ5_2_LC_12_6_2 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \b2v_inst11.count_clk_RNIVSLQ5_2_LC_12_6_2  (
            .in0(N__32831),
            .in1(N__32823),
            .in2(N__33809),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_count_clk_2_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_2_LC_12_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_2_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_2_LC_12_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_2_LC_12_6_3  (
            .in0(N__32822),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37006),
            .ce(N__33767),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVSLQ5_0_2_LC_12_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVSLQ5_0_2_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVSLQ5_0_2_LC_12_6_4 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \b2v_inst11.count_clk_RNIVSLQ5_0_2_LC_12_6_4  (
            .in0(N__32832),
            .in1(N__32821),
            .in2(N__33811),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI7RAQ5_15_LC_12_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI7RAQ5_15_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI7RAQ5_15_LC_12_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI7RAQ5_15_LC_12_6_5  (
            .in0(N__33894),
            .in1(N__33885),
            .in2(_gnd_net_),
            .in3(N__33768),
            .lcout(\b2v_inst11.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_15_LC_12_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_15_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_15_LC_12_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_15_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33893),
            .lcout(\b2v_inst11.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37006),
            .ce(N__33767),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI79QQ5_6_LC_12_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI79QQ5_6_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI79QQ5_6_LC_12_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI79QQ5_6_LC_12_6_7  (
            .in0(N__33869),
            .in1(N__33855),
            .in2(_gnd_net_),
            .in3(N__33763),
            .lcout(\b2v_inst11.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIK0DK3_0_LC_12_7_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIK0DK3_0_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIK0DK3_0_LC_12_7_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \b2v_inst6.curr_state_RNIK0DK3_0_LC_12_7_0  (
            .in0(N__33239),
            .in1(N__33612),
            .in2(_gnd_net_),
            .in3(N__35864),
            .lcout(\b2v_inst6.count_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_0_LC_12_7_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_0_LC_12_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.count_RNI_0_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33591),
            .lcout(\b2v_inst6.N_2994_i ),
            .ltout(\b2v_inst6.N_2994_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_0_LC_12_7_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_LC_12_7_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_0_LC_12_7_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst6.count_0_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__33229),
            .in2(N__33534),
            .in3(N__33531),
            .lcout(\b2v_inst6.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37100),
            .ce(N__33407),
            .sr(N__33238));
    defparam \b2v_inst6.count_15_LC_12_7_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_15_LC_12_7_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_15_LC_12_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_15_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33492),
            .lcout(\b2v_inst6.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37100),
            .ce(N__33407),
            .sr(N__33238));
    defparam \b2v_inst11.func_state_RNI_4_1_LC_12_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_4_1_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_4_1_LC_12_7_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.func_state_RNI_4_1_LC_12_7_5  (
            .in0(N__34026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.func_state_RNI_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_5_1_LC_12_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_5_1_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_5_1_LC_12_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNI_5_1_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34025),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_5_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_7_LC_12_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_7_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_7_LC_12_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_7_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34166),
            .lcout(\b2v_inst11.N_200_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITSFK3_6_LC_12_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITSFK3_6_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITSFK3_6_LC_12_8_0 .LUT_INIT=16'b1111111001001110;
    LogicCell40 \b2v_inst11.dutycycle_RNITSFK3_6_LC_12_8_0  (
            .in0(N__38228),
            .in1(N__37178),
            .in2(N__34837),
            .in3(N__34065),
            .lcout(),
            .ltout(\b2v_inst11.N_231_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIJS2L6_6_LC_12_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIJS2L6_6_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIJS2L6_6_LC_12_8_1 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIJS2L6_6_LC_12_8_1  (
            .in0(N__34131),
            .in1(N__34119),
            .in2(N__34110),
            .in3(N__37278),
            .lcout(\b2v_inst11.dutycycle_eena_13 ),
            .ltout(\b2v_inst11.dutycycle_eena_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_6_LC_12_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_6_LC_12_8_2 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_6_LC_12_8_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst11.dutycycle_6_LC_12_8_2  (
            .in0(N__34098),
            .in1(N__34104),
            .in2(N__34107),
            .in3(N__35859),
            .lcout(\b2v_inst11.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37085),
            .ce(),
            .sr(N__36362));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVB4_LC_12_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVB4_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVB4_LC_12_8_3 .LUT_INIT=16'b1111111100110111;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVB4_LC_12_8_3  (
            .in0(N__33941),
            .in1(N__37277),
            .in2(N__34048),
            .in3(N__35244),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4 ),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5IIRB_6_LC_12_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5IIRB_6_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5IIRB_6_LC_12_8_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI5IIRB_6_LC_12_8_4  (
            .in0(N__34097),
            .in1(N__35857),
            .in2(N__34089),
            .in3(N__34086),
            .lcout(\b2v_inst11.dutycycleZ1Z_6 ),
            .ltout(\b2v_inst11.dutycycleZ1Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNILF063_6_LC_12_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNILF063_6_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNILF063_6_LC_12_8_5 .LUT_INIT=16'b0000010011110100;
    LogicCell40 \b2v_inst11.dutycycle_RNILF063_6_LC_12_8_5  (
            .in0(N__34030),
            .in1(N__34080),
            .in2(N__34068),
            .in3(N__37617),
            .lcout(\b2v_inst11.dutycycle_RNILF063Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNI1GBN4_LC_12_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNI1GBN4_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNI1GBN4_LC_12_8_6 .LUT_INIT=16'b1111111100011111;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNI1GBN4_LC_12_8_6  (
            .in0(N__34031),
            .in1(N__33942),
            .in2(N__37316),
            .in3(N__35271),
            .lcout(\b2v_inst11.dutycycle_set_1 ),
            .ltout(\b2v_inst11.dutycycle_set_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_5_LC_12_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_5_LC_12_8_7 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_5_LC_12_8_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst11.dutycycle_5_LC_12_8_7  (
            .in0(N__35858),
            .in1(N__34451),
            .in2(N__34479),
            .in3(N__34476),
            .lcout(\b2v_inst11.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37085),
            .ce(),
            .sr(N__36362));
    defparam \b2v_inst11.dutycycle_RNIOFQO2_3_LC_12_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIOFQO2_3_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIOFQO2_3_LC_12_9_2 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \b2v_inst11.dutycycle_RNIOFQO2_3_LC_12_9_2  (
            .in0(N__37507),
            .in1(N__34322),
            .in2(N__37179),
            .in3(N__37426),
            .lcout(\b2v_inst11.dutycycle_RNIOFQO2Z0Z_3 ),
            .ltout(\b2v_inst11.dutycycle_RNIOFQO2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_3_LC_12_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_3_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_3_LC_12_9_3 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \b2v_inst11.dutycycle_3_LC_12_9_3  (
            .in0(N__34412),
            .in1(N__34422),
            .in2(N__34437),
            .in3(N__37283),
            .lcout(\b2v_inst11.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37070),
            .ce(),
            .sr(N__36368));
    defparam \b2v_inst11.dutycycle_RNIM98E2_3_LC_12_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIM98E2_3_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIM98E2_3_LC_12_9_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNIM98E2_3_LC_12_9_4  (
            .in0(N__35835),
            .in1(N__34434),
            .in2(N__34416),
            .in3(N__36220),
            .lcout(\b2v_inst11.dutycycle_RNIM98E2Z0Z_3 ),
            .ltout(\b2v_inst11.dutycycle_RNIM98E2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI51C57_3_LC_12_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI51C57_3_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI51C57_3_LC_12_9_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \b2v_inst11.dutycycle_RNI51C57_3_LC_12_9_5  (
            .in0(N__34411),
            .in1(N__37282),
            .in2(N__34398),
            .in3(N__34395),
            .lcout(\b2v_inst11.dutycycleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_12_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_12_9_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_12_9_6  (
            .in0(N__39280),
            .in1(N__34266),
            .in2(N__38391),
            .in3(N__34819),
            .lcout(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ),
            .ltout(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIOMFH6_13_LC_12_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIOMFH6_13_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIOMFH6_13_LC_12_9_7 .LUT_INIT=16'b0100111100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIOMFH6_13_LC_12_9_7  (
            .in0(N__37427),
            .in1(N__34497),
            .in2(N__34212),
            .in3(N__35834),
            .lcout(\b2v_inst11.dutycycle_en_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_12_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_12_10_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_12_10_0  (
            .in0(N__36215),
            .in1(N__38813),
            .in2(_gnd_net_),
            .in3(N__37431),
            .lcout(\b2v_inst11.un1_clk_100khz_32_and_i_0_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_12_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_12_10_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_8_LC_12_10_1  (
            .in0(N__37433),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37876),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_32_and_i_0_c_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI484S5_8_LC_12_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI484S5_8_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI484S5_8_LC_12_10_2 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \b2v_inst11.dutycycle_RNI484S5_8_LC_12_10_2  (
            .in0(N__34509),
            .in1(N__37290),
            .in2(N__34512),
            .in3(N__37502),
            .lcout(\b2v_inst11.dutycycle_eena_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_12_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_12_10_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_10_LC_12_10_3  (
            .in0(N__37432),
            .in1(_gnd_net_),
            .in2(N__35461),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_33_and_i_0_c_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI484S5_10_LC_12_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI484S5_10_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI484S5_10_LC_12_10_4 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \b2v_inst11.dutycycle_RNI484S5_10_LC_12_10_4  (
            .in0(N__34508),
            .in1(N__37289),
            .in2(N__34500),
            .in3(N__37501),
            .lcout(\b2v_inst11.dutycycle_eena_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5AV24_13_LC_12_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5AV24_13_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5AV24_13_LC_12_10_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI5AV24_13_LC_12_10_5  (
            .in0(N__38814),
            .in1(N__34607),
            .in2(N__37512),
            .in3(N__36216),
            .lcout(\b2v_inst11.N_153_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5AV24_14_LC_12_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5AV24_14_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5AV24_14_LC_12_10_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI5AV24_14_LC_12_10_6  (
            .in0(N__35205),
            .in1(N__37506),
            .in2(N__36231),
            .in3(N__38815),
            .lcout(),
            .ltout(\b2v_inst11.N_155_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIOMFH6_14_LC_12_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIOMFH6_14_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIOMFH6_14_LC_12_10_7 .LUT_INIT=16'b0100000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIOMFH6_14_LC_12_10_7  (
            .in0(N__37434),
            .in1(N__35788),
            .in2(N__34491),
            .in3(N__37291),
            .lcout(\b2v_inst11.dutycycle_en_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIG6AA9_7_LC_12_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIG6AA9_7_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIG6AA9_7_LC_12_11_0 .LUT_INIT=16'b0000110001001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIG6AA9_7_LC_12_11_0  (
            .in0(N__34485),
            .in1(N__35845),
            .in2(N__37323),
            .in3(N__34716),
            .lcout(\b2v_inst11.g0_0_1_0 ),
            .ltout(\b2v_inst11.g0_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_7_LC_12_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_7_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_7_LC_12_11_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.dutycycle_7_LC_12_11_1  (
            .in0(N__34686),
            .in1(N__34674),
            .in2(N__34488),
            .in3(N__36210),
            .lcout(\b2v_inst11.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37144),
            .ce(),
            .sr(N__36348));
    defparam \b2v_inst11.dutycycle_RNI5AV24_7_LC_12_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5AV24_7_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5AV24_7_LC_12_11_2 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI5AV24_7_LC_12_11_2  (
            .in0(N__36209),
            .in1(N__37981),
            .in2(_gnd_net_),
            .in3(N__37509),
            .lcout(\b2v_inst11.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIG2BA2_0_0_LC_12_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIG2BA2_0_0_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIG2BA2_0_0_LC_12_11_3 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \b2v_inst11.func_state_RNIG2BA2_0_0_LC_12_11_3  (
            .in0(N__35530),
            .in1(N__34854),
            .in2(N__38742),
            .in3(N__38812),
            .lcout(\b2v_inst11.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_7_LC_12_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_7_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_7_LC_12_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_7_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37980),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_7 ),
            .ltout(\b2v_inst11.dutycycle_RNI_7Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIOFQO2_7_LC_12_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIOFQO2_7_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIOFQO2_7_LC_12_11_5 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIOFQO2_7_LC_12_11_5  (
            .in0(N__37428),
            .in1(N__34838),
            .in2(N__34725),
            .in3(N__34722),
            .lcout(\b2v_inst11.un1_clk_100khz_36_and_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNI5V4S_LC_12_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNI5V4S_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNI5V4S_LC_12_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNI5V4S_LC_12_11_6  (
            .in0(N__34710),
            .in1(N__34698),
            .in2(_gnd_net_),
            .in3(N__36050),
            .lcout(\b2v_inst11.un1_dutycycle_94_0_7 ),
            .ltout(\b2v_inst11.un1_dutycycle_94_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIUDOLB_7_LC_12_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIUDOLB_7_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIUDOLB_7_LC_12_11_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNIUDOLB_7_LC_12_11_7  (
            .in0(N__34680),
            .in1(N__34673),
            .in2(N__34665),
            .in3(N__36208),
            .lcout(\b2v_inst11.dutycycleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_13_LC_12_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_13_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_13_LC_12_12_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst11.dutycycle_13_LC_12_12_0  (
            .in0(N__34641),
            .in1(N__34622),
            .in2(N__34635),
            .in3(N__36207),
            .lcout(\b2v_inst11.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37086),
            .ce(),
            .sr(N__36361));
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQ_LC_12_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQ_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQ_LC_12_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQ_LC_12_12_1  (
            .in0(N__36005),
            .in1(N__34662),
            .in2(_gnd_net_),
            .in3(N__34650),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0 ),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDSSV8_13_LC_12_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDSSV8_13_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDSSV8_13_LC_12_12_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNIDSSV8_13_LC_12_12_2  (
            .in0(N__34631),
            .in1(N__34623),
            .in2(N__34611),
            .in3(N__36204),
            .lcout(\b2v_inst11.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIE51T1_LC_12_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIE51T1_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIE51T1_LC_12_12_3 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIE51T1_LC_12_12_3  (
            .in0(N__36203),
            .in1(N__36057),
            .in2(N__35289),
            .in3(N__35280),
            .lcout(\b2v_inst11.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIGFLH1_LC_12_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIGFLH1_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIGFLH1_LC_12_12_4 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIGFLH1_LC_12_12_4  (
            .in0(N__36058),
            .in1(N__35262),
            .in2(N__36221),
            .in3(N__35250),
            .lcout(\b2v_inst11.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IF_LC_12_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IF_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IF_LC_12_12_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IF_LC_12_12_5  (
            .in0(N__35232),
            .in1(_gnd_net_),
            .in2(N__36042),
            .in3(N__35223),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0 ),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIG7HK8_14_LC_12_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIG7HK8_14_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIG7HK8_14_LC_12_12_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNIG7HK8_14_LC_12_12_6  (
            .in0(N__35109),
            .in1(N__35093),
            .in2(N__35214),
            .in3(N__36205),
            .lcout(\b2v_inst11.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_14_LC_12_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_14_LC_12_12_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_14_LC_12_12_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst11.dutycycle_14_LC_12_12_7  (
            .in0(N__36206),
            .in1(N__35115),
            .in2(N__35097),
            .in3(N__35108),
            .lcout(\b2v_inst11.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37086),
            .ce(),
            .sr(N__36361));
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_12_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_12_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_10_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35422),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_10 ),
            .ltout(\b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_12_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_12_13_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_4_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35031),
            .in3(N__35015),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_44_0_3_tz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_12_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_12_13_2 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_8_LC_12_13_2  (
            .in0(N__35537),
            .in1(N__38108),
            .in2(N__34878),
            .in3(N__37881),
            .lcout(\b2v_inst11.un1_dutycycle_53_44_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_10_LC_12_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_10_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_10_LC_12_13_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \b2v_inst11.dutycycle_10_LC_12_13_3  (
            .in0(N__35589),
            .in1(N__35571),
            .in2(N__35583),
            .in3(N__35837),
            .lcout(\b2v_inst11.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37142),
            .ce(),
            .sr(N__36366));
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNION642_LC_12_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNION642_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNION642_LC_12_13_4 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNION642_LC_12_13_4  (
            .in0(N__35607),
            .in1(N__36229),
            .in2(N__36041),
            .in3(N__35595),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642 ),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIM01V8_10_LC_12_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIM01V8_10_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIM01V8_10_LC_12_13_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIM01V8_10_LC_12_13_5  (
            .in0(N__35579),
            .in1(N__35570),
            .in2(N__35559),
            .in3(N__35836),
            .lcout(\b2v_inst11.dutycycleZ0Z_3 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_LC_12_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_12_13_6 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_LC_12_13_6  (
            .in0(N__35536),
            .in1(N__38106),
            .in2(N__35493),
            .in3(N__37877),
            .lcout(\b2v_inst11.un1_dutycycle_53_44_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_10_LC_12_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_10_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_10_LC_12_13_7 .LUT_INIT=16'b0000010111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_10_LC_12_13_7  (
            .in0(N__38107),
            .in1(_gnd_net_),
            .in2(N__37910),
            .in3(N__35423),
            .lcout(\b2v_inst11.g1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI484S5_9_LC_12_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI484S5_9_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI484S5_9_LC_12_14_0 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI484S5_9_LC_12_14_0  (
            .in0(N__37293),
            .in1(N__37511),
            .in2(N__35298),
            .in3(N__37168),
            .lcout(\b2v_inst11.dutycycle_eena_2 ),
            .ltout(\b2v_inst11.dutycycle_eena_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICK668_9_LC_12_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICK668_9_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICK668_9_LC_12_14_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \b2v_inst11.dutycycle_RNICK668_9_LC_12_14_1  (
            .in0(N__35349),
            .in1(N__35830),
            .in2(N__35328),
            .in3(N__35318),
            .lcout(\b2v_inst11.dutycycleZ0Z_0 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_9_LC_12_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_9_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIDQ4A1_9_LC_12_14_2 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \b2v_inst11.dutycycle_RNIDQ4A1_9_LC_12_14_2  (
            .in0(N__38802),
            .in1(N__36225),
            .in2(N__35301),
            .in3(N__37429),
            .lcout(\b2v_inst11.un1_clk_100khz_30_and_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIJI598_15_LC_12_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIJI598_15_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIJI598_15_LC_12_14_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIJI598_15_LC_12_14_3  (
            .in0(N__36228),
            .in1(N__37203),
            .in2(N__37191),
            .in3(N__37209),
            .lcout(\b2v_inst11.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5AV24_15_LC_12_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5AV24_15_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5AV24_15_LC_12_14_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI5AV24_15_LC_12_14_4  (
            .in0(N__38803),
            .in1(N__36227),
            .in2(N__37582),
            .in3(N__37510),
            .lcout(),
            .ltout(\b2v_inst11.N_158_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIOMFH6_15_LC_12_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIOMFH6_15_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIOMFH6_15_LC_12_14_5 .LUT_INIT=16'b0100000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIOMFH6_15_LC_12_14_5  (
            .in0(N__37430),
            .in1(N__35829),
            .in2(N__37365),
            .in3(N__37292),
            .lcout(\b2v_inst11.dutycycle_en_12 ),
            .ltout(\b2v_inst11.dutycycle_en_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_15_LC_12_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_15_LC_12_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_15_LC_12_14_6 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.dutycycle_15_LC_12_14_6  (
            .in0(N__37202),
            .in1(N__37190),
            .in2(N__37194),
            .in3(N__36226),
            .lcout(\b2v_inst11.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37127),
            .ce(),
            .sr(N__36369));
    defparam \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_12_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_12_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__36222),
            .in2(_gnd_net_),
            .in3(N__38801),
            .lcout(\b2v_inst11.N_326_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_8_LC_12_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_8_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_8_LC_12_15_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \b2v_inst11.dutycycle_8_LC_12_15_0  (
            .in0(N__35889),
            .in1(N__35880),
            .in2(N__35865),
            .in3(N__35895),
            .lcout(\b2v_inst11.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37149),
            .ce(),
            .sr(N__36367));
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQ1_LC_12_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQ1_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQ1_LC_12_15_1 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQ1_LC_12_15_1  (
            .in0(N__36246),
            .in1(N__36223),
            .in2(N__36078),
            .in3(N__36037),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1 ),
            .ltout(\b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI99IH8_8_LC_12_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI99IH8_8_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI99IH8_8_LC_12_15_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI99IH8_8_LC_12_15_2  (
            .in0(N__35888),
            .in1(N__35879),
            .in2(N__35868),
            .in3(N__35860),
            .lcout(\b2v_inst11.dutycycleZ0Z_4 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_12_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_12_15_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_7_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35610),
            .in3(N__38030),
            .lcout(\b2v_inst11.un1_i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_12_LC_12_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_12_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_12_LC_12_15_4  (
            .in0(N__37873),
            .in1(N__38121),
            .in2(N__38341),
            .in3(N__37757),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_12_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_12_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_7_LC_12_15_5  (
            .in0(N__38122),
            .in1(N__38031),
            .in2(N__37770),
            .in3(N__37874),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_12_7_LC_12_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_12_7_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_12_7_LC_12_15_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_12_7_LC_12_15_6  (
            .in0(N__37791),
            .in1(N__37785),
            .in2(N__37779),
            .in3(N__37776),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_s_9_sf_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_12_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_12_15_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_12_LC_12_15_7  (
            .in0(N__37761),
            .in1(_gnd_net_),
            .in2(N__37656),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_0_1_LC_12_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_0_1_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_0_1_LC_12_16_0 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_0_1_LC_12_16_0  (
            .in0(N__37602),
            .in1(N__38587),
            .in2(N__38849),
            .in3(N__39182),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_clk_100khz_42_and_i_a2_5_LC_12_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_clk_100khz_42_and_i_a2_5_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_clk_100khz_42_and_i_a2_5_LC_12_16_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.un1_clk_100khz_42_and_i_a2_5_LC_12_16_1  (
            .in0(N__39283),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38526),
            .lcout(),
            .ltout(\b2v_inst11.N_371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_1_1_LC_12_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_1_1_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_1_1_LC_12_16_2 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_1_1_LC_12_16_2  (
            .in0(N__38590),
            .in1(N__39183),
            .in2(N__37623),
            .in3(N__38832),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDUQ02_1_LC_12_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDUQ02_1_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDUQ02_1_LC_12_16_3 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \b2v_inst11.func_state_RNIDUQ02_1_LC_12_16_3  (
            .in0(N__38588),
            .in1(_gnd_net_),
            .in2(N__37620),
            .in3(N__38523),
            .lcout(\b2v_inst11.func_state_RNIDUQ02Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.g2_0_0_0_LC_12_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.g2_0_0_0_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.g2_0_0_0_LC_12_16_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst11.g2_0_0_0_LC_12_16_4  (
            .in0(N__38524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39281),
            .lcout(\b2v_inst11.g2_0_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.g2_3_0_LC_12_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.g2_3_0_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.g2_3_0_LC_12_16_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.g2_3_0_LC_12_16_5  (
            .in0(N__39282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38525),
            .lcout(),
            .ltout(\b2v_inst11.g2_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8H551_1_LC_12_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8H551_1_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8H551_1_LC_12_16_6 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \b2v_inst11.func_state_RNI8H551_1_LC_12_16_6  (
            .in0(N__38591),
            .in1(N__39181),
            .in2(N__38862),
            .in3(N__38831),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_12_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_12_16_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_12_16_7  (
            .in0(N__38589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38527),
            .lcout(\b2v_inst11.N_161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TOP
