// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 9 2022 11:23:42

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    output SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__36183;
    wire N__36182;
    wire N__36181;
    wire N__36174;
    wire N__36173;
    wire N__36172;
    wire N__36165;
    wire N__36164;
    wire N__36163;
    wire N__36156;
    wire N__36155;
    wire N__36154;
    wire N__36147;
    wire N__36146;
    wire N__36145;
    wire N__36138;
    wire N__36137;
    wire N__36136;
    wire N__36129;
    wire N__36128;
    wire N__36127;
    wire N__36120;
    wire N__36119;
    wire N__36118;
    wire N__36111;
    wire N__36110;
    wire N__36109;
    wire N__36102;
    wire N__36101;
    wire N__36100;
    wire N__36093;
    wire N__36092;
    wire N__36091;
    wire N__36084;
    wire N__36083;
    wire N__36082;
    wire N__36075;
    wire N__36074;
    wire N__36073;
    wire N__36066;
    wire N__36065;
    wire N__36064;
    wire N__36057;
    wire N__36056;
    wire N__36055;
    wire N__36048;
    wire N__36047;
    wire N__36046;
    wire N__36039;
    wire N__36038;
    wire N__36037;
    wire N__36030;
    wire N__36029;
    wire N__36028;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36003;
    wire N__36002;
    wire N__36001;
    wire N__35994;
    wire N__35993;
    wire N__35992;
    wire N__35985;
    wire N__35984;
    wire N__35983;
    wire N__35976;
    wire N__35975;
    wire N__35974;
    wire N__35967;
    wire N__35966;
    wire N__35965;
    wire N__35958;
    wire N__35957;
    wire N__35956;
    wire N__35949;
    wire N__35948;
    wire N__35947;
    wire N__35940;
    wire N__35939;
    wire N__35938;
    wire N__35931;
    wire N__35930;
    wire N__35929;
    wire N__35922;
    wire N__35921;
    wire N__35920;
    wire N__35913;
    wire N__35912;
    wire N__35911;
    wire N__35904;
    wire N__35903;
    wire N__35902;
    wire N__35895;
    wire N__35894;
    wire N__35893;
    wire N__35886;
    wire N__35885;
    wire N__35884;
    wire N__35877;
    wire N__35876;
    wire N__35875;
    wire N__35868;
    wire N__35867;
    wire N__35866;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35850;
    wire N__35849;
    wire N__35848;
    wire N__35841;
    wire N__35840;
    wire N__35839;
    wire N__35832;
    wire N__35831;
    wire N__35830;
    wire N__35823;
    wire N__35822;
    wire N__35821;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35805;
    wire N__35804;
    wire N__35803;
    wire N__35796;
    wire N__35795;
    wire N__35794;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35769;
    wire N__35768;
    wire N__35767;
    wire N__35760;
    wire N__35759;
    wire N__35758;
    wire N__35751;
    wire N__35750;
    wire N__35749;
    wire N__35742;
    wire N__35741;
    wire N__35740;
    wire N__35733;
    wire N__35732;
    wire N__35731;
    wire N__35724;
    wire N__35723;
    wire N__35722;
    wire N__35715;
    wire N__35714;
    wire N__35713;
    wire N__35706;
    wire N__35705;
    wire N__35704;
    wire N__35697;
    wire N__35696;
    wire N__35695;
    wire N__35688;
    wire N__35687;
    wire N__35686;
    wire N__35679;
    wire N__35678;
    wire N__35677;
    wire N__35670;
    wire N__35669;
    wire N__35668;
    wire N__35661;
    wire N__35660;
    wire N__35659;
    wire N__35642;
    wire N__35641;
    wire N__35638;
    wire N__35637;
    wire N__35636;
    wire N__35635;
    wire N__35634;
    wire N__35633;
    wire N__35630;
    wire N__35629;
    wire N__35626;
    wire N__35625;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35586;
    wire N__35583;
    wire N__35576;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35561;
    wire N__35558;
    wire N__35557;
    wire N__35552;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35541;
    wire N__35540;
    wire N__35537;
    wire N__35534;
    wire N__35533;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35512;
    wire N__35507;
    wire N__35504;
    wire N__35495;
    wire N__35492;
    wire N__35491;
    wire N__35490;
    wire N__35485;
    wire N__35482;
    wire N__35481;
    wire N__35480;
    wire N__35477;
    wire N__35476;
    wire N__35475;
    wire N__35474;
    wire N__35473;
    wire N__35472;
    wire N__35471;
    wire N__35470;
    wire N__35467;
    wire N__35462;
    wire N__35459;
    wire N__35458;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35450;
    wire N__35449;
    wire N__35448;
    wire N__35447;
    wire N__35446;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35439;
    wire N__35430;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35409;
    wire N__35404;
    wire N__35403;
    wire N__35394;
    wire N__35391;
    wire N__35390;
    wire N__35385;
    wire N__35380;
    wire N__35379;
    wire N__35378;
    wire N__35377;
    wire N__35374;
    wire N__35369;
    wire N__35366;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35351;
    wire N__35346;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35294;
    wire N__35289;
    wire N__35286;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35272;
    wire N__35269;
    wire N__35264;
    wire N__35259;
    wire N__35256;
    wire N__35249;
    wire N__35240;
    wire N__35237;
    wire N__35232;
    wire N__35225;
    wire N__35220;
    wire N__35213;
    wire N__35210;
    wire N__35209;
    wire N__35208;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35195;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35183;
    wire N__35180;
    wire N__35177;
    wire N__35176;
    wire N__35175;
    wire N__35172;
    wire N__35165;
    wire N__35160;
    wire N__35153;
    wire N__35152;
    wire N__35149;
    wire N__35148;
    wire N__35145;
    wire N__35144;
    wire N__35143;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35135;
    wire N__35132;
    wire N__35131;
    wire N__35128;
    wire N__35127;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35119;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35111;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35086;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35050;
    wire N__35049;
    wire N__35044;
    wire N__35041;
    wire N__35036;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35004;
    wire N__34995;
    wire N__34992;
    wire N__34987;
    wire N__34982;
    wire N__34977;
    wire N__34970;
    wire N__34969;
    wire N__34968;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34960;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34937;
    wire N__34936;
    wire N__34935;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34901;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34821;
    wire N__34816;
    wire N__34815;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34811;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34803;
    wire N__34794;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34784;
    wire N__34783;
    wire N__34782;
    wire N__34779;
    wire N__34772;
    wire N__34761;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34741;
    wire N__34740;
    wire N__34739;
    wire N__34738;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34725;
    wire N__34724;
    wire N__34721;
    wire N__34720;
    wire N__34719;
    wire N__34718;
    wire N__34717;
    wire N__34716;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34660;
    wire N__34657;
    wire N__34656;
    wire N__34655;
    wire N__34652;
    wire N__34651;
    wire N__34650;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34622;
    wire N__34621;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34600;
    wire N__34597;
    wire N__34596;
    wire N__34593;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34585;
    wire N__34584;
    wire N__34583;
    wire N__34582;
    wire N__34577;
    wire N__34574;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34557;
    wire N__34554;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34540;
    wire N__34539;
    wire N__34534;
    wire N__34533;
    wire N__34532;
    wire N__34525;
    wire N__34522;
    wire N__34517;
    wire N__34514;
    wire N__34513;
    wire N__34506;
    wire N__34499;
    wire N__34496;
    wire N__34495;
    wire N__34492;
    wire N__34491;
    wire N__34490;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34465;
    wire N__34464;
    wire N__34463;
    wire N__34460;
    wire N__34455;
    wire N__34452;
    wire N__34451;
    wire N__34444;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34416;
    wire N__34409;
    wire N__34406;
    wire N__34405;
    wire N__34404;
    wire N__34403;
    wire N__34400;
    wire N__34399;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34380;
    wire N__34377;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34354;
    wire N__34347;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34326;
    wire N__34323;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34307;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34265;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34254;
    wire N__34251;
    wire N__34246;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34227;
    wire N__34222;
    wire N__34219;
    wire N__34210;
    wire N__34207;
    wire N__34202;
    wire N__34199;
    wire N__34198;
    wire N__34195;
    wire N__34190;
    wire N__34179;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34160;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34138;
    wire N__34135;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34112;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34089;
    wire N__34082;
    wire N__34071;
    wire N__34064;
    wire N__34063;
    wire N__34062;
    wire N__34061;
    wire N__34056;
    wire N__34047;
    wire N__34040;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__33999;
    wire N__33998;
    wire N__33997;
    wire N__33996;
    wire N__33993;
    wire N__33992;
    wire N__33989;
    wire N__33988;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33984;
    wire N__33983;
    wire N__33982;
    wire N__33979;
    wire N__33978;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33957;
    wire N__33956;
    wire N__33955;
    wire N__33948;
    wire N__33945;
    wire N__33944;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33934;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33918;
    wire N__33917;
    wire N__33916;
    wire N__33915;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33865;
    wire N__33858;
    wire N__33841;
    wire N__33824;
    wire N__33821;
    wire N__33820;
    wire N__33819;
    wire N__33818;
    wire N__33817;
    wire N__33812;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33804;
    wire N__33803;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33795;
    wire N__33794;
    wire N__33793;
    wire N__33790;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33776;
    wire N__33773;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33748;
    wire N__33743;
    wire N__33740;
    wire N__33739;
    wire N__33738;
    wire N__33737;
    wire N__33736;
    wire N__33735;
    wire N__33728;
    wire N__33725;
    wire N__33718;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33697;
    wire N__33690;
    wire N__33677;
    wire N__33674;
    wire N__33673;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33667;
    wire N__33666;
    wire N__33663;
    wire N__33662;
    wire N__33661;
    wire N__33660;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33652;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33644;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33635;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33607;
    wire N__33604;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33600;
    wire N__33595;
    wire N__33590;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33571;
    wire N__33566;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33548;
    wire N__33545;
    wire N__33544;
    wire N__33543;
    wire N__33540;
    wire N__33533;
    wire N__33528;
    wire N__33523;
    wire N__33518;
    wire N__33515;
    wire N__33510;
    wire N__33505;
    wire N__33502;
    wire N__33497;
    wire N__33494;
    wire N__33489;
    wire N__33484;
    wire N__33479;
    wire N__33470;
    wire N__33455;
    wire N__33452;
    wire N__33451;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33436;
    wire N__33435;
    wire N__33434;
    wire N__33433;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33404;
    wire N__33403;
    wire N__33402;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33386;
    wire N__33377;
    wire N__33376;
    wire N__33373;
    wire N__33372;
    wire N__33371;
    wire N__33370;
    wire N__33369;
    wire N__33368;
    wire N__33367;
    wire N__33366;
    wire N__33365;
    wire N__33364;
    wire N__33363;
    wire N__33362;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33358;
    wire N__33355;
    wire N__33350;
    wire N__33349;
    wire N__33346;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33330;
    wire N__33327;
    wire N__33318;
    wire N__33313;
    wire N__33308;
    wire N__33303;
    wire N__33302;
    wire N__33301;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33280;
    wire N__33273;
    wire N__33268;
    wire N__33263;
    wire N__33258;
    wire N__33253;
    wire N__33248;
    wire N__33243;
    wire N__33236;
    wire N__33231;
    wire N__33228;
    wire N__33223;
    wire N__33218;
    wire N__33215;
    wire N__33208;
    wire N__33193;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33145;
    wire N__33144;
    wire N__33143;
    wire N__33142;
    wire N__33141;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33134;
    wire N__33133;
    wire N__33132;
    wire N__33129;
    wire N__33128;
    wire N__33125;
    wire N__33124;
    wire N__33123;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33108;
    wire N__33107;
    wire N__33106;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33090;
    wire N__33089;
    wire N__33088;
    wire N__33087;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33065;
    wire N__33062;
    wire N__33057;
    wire N__33056;
    wire N__33053;
    wire N__33052;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33035;
    wire N__33028;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32997;
    wire N__32994;
    wire N__32985;
    wire N__32976;
    wire N__32973;
    wire N__32960;
    wire N__32959;
    wire N__32958;
    wire N__32957;
    wire N__32954;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32946;
    wire N__32943;
    wire N__32942;
    wire N__32941;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32926;
    wire N__32921;
    wire N__32916;
    wire N__32911;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32881;
    wire N__32880;
    wire N__32877;
    wire N__32872;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32847;
    wire N__32846;
    wire N__32845;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32837;
    wire N__32836;
    wire N__32833;
    wire N__32832;
    wire N__32831;
    wire N__32830;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32814;
    wire N__32813;
    wire N__32812;
    wire N__32807;
    wire N__32802;
    wire N__32797;
    wire N__32790;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32773;
    wire N__32772;
    wire N__32771;
    wire N__32770;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32731;
    wire N__32728;
    wire N__32721;
    wire N__32710;
    wire N__32701;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32676;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32659;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32638;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32630;
    wire N__32625;
    wire N__32622;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32602;
    wire N__32599;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32585;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32541;
    wire N__32540;
    wire N__32535;
    wire N__32530;
    wire N__32529;
    wire N__32528;
    wire N__32525;
    wire N__32524;
    wire N__32523;
    wire N__32518;
    wire N__32513;
    wire N__32510;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32484;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32472;
    wire N__32457;
    wire N__32450;
    wire N__32445;
    wire N__32442;
    wire N__32437;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32420;
    wire N__32415;
    wire N__32408;
    wire N__32407;
    wire N__32406;
    wire N__32403;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32395;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32387;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32377;
    wire N__32376;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32361;
    wire N__32356;
    wire N__32353;
    wire N__32352;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32333;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32312;
    wire N__32309;
    wire N__32308;
    wire N__32307;
    wire N__32302;
    wire N__32295;
    wire N__32290;
    wire N__32285;
    wire N__32276;
    wire N__32275;
    wire N__32274;
    wire N__32273;
    wire N__32272;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32262;
    wire N__32259;
    wire N__32258;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32250;
    wire N__32249;
    wire N__32248;
    wire N__32245;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32230;
    wire N__32229;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32197;
    wire N__32194;
    wire N__32193;
    wire N__32192;
    wire N__32187;
    wire N__32182;
    wire N__32179;
    wire N__32172;
    wire N__32169;
    wire N__32164;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32132;
    wire N__32129;
    wire N__32120;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32081;
    wire N__32076;
    wire N__32071;
    wire N__32068;
    wire N__32065;
    wire N__32064;
    wire N__32063;
    wire N__32062;
    wire N__32059;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32041;
    wire N__32030;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32022;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32014;
    wire N__32013;
    wire N__32012;
    wire N__32009;
    wire N__32008;
    wire N__32007;
    wire N__32004;
    wire N__32003;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31991;
    wire N__31988;
    wire N__31987;
    wire N__31984;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31959;
    wire N__31956;
    wire N__31955;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31932;
    wire N__31929;
    wire N__31924;
    wire N__31921;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31903;
    wire N__31892;
    wire N__31891;
    wire N__31888;
    wire N__31887;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31870;
    wire N__31869;
    wire N__31868;
    wire N__31865;
    wire N__31864;
    wire N__31861;
    wire N__31856;
    wire N__31853;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31837;
    wire N__31826;
    wire N__31825;
    wire N__31824;
    wire N__31823;
    wire N__31822;
    wire N__31821;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31813;
    wire N__31812;
    wire N__31811;
    wire N__31810;
    wire N__31809;
    wire N__31808;
    wire N__31807;
    wire N__31804;
    wire N__31799;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31789;
    wire N__31786;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31774;
    wire N__31773;
    wire N__31770;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31756;
    wire N__31753;
    wire N__31752;
    wire N__31751;
    wire N__31750;
    wire N__31747;
    wire N__31746;
    wire N__31743;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31723;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31701;
    wire N__31692;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31665;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31627;
    wire N__31622;
    wire N__31619;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31600;
    wire N__31597;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31585;
    wire N__31582;
    wire N__31581;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31570;
    wire N__31569;
    wire N__31568;
    wire N__31567;
    wire N__31564;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31543;
    wire N__31540;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31494;
    wire N__31491;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31455;
    wire N__31452;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31415;
    wire N__31414;
    wire N__31413;
    wire N__31412;
    wire N__31411;
    wire N__31410;
    wire N__31409;
    wire N__31408;
    wire N__31407;
    wire N__31406;
    wire N__31405;
    wire N__31404;
    wire N__31403;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31395;
    wire N__31388;
    wire N__31387;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31352;
    wire N__31349;
    wire N__31348;
    wire N__31347;
    wire N__31346;
    wire N__31345;
    wire N__31342;
    wire N__31341;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31329;
    wire N__31326;
    wire N__31319;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31303;
    wire N__31298;
    wire N__31295;
    wire N__31290;
    wire N__31283;
    wire N__31276;
    wire N__31259;
    wire N__31258;
    wire N__31257;
    wire N__31256;
    wire N__31255;
    wire N__31254;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31245;
    wire N__31244;
    wire N__31243;
    wire N__31242;
    wire N__31235;
    wire N__31234;
    wire N__31231;
    wire N__31230;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31224;
    wire N__31221;
    wire N__31220;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31216;
    wire N__31215;
    wire N__31212;
    wire N__31207;
    wire N__31204;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31188;
    wire N__31183;
    wire N__31176;
    wire N__31173;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31147;
    wire N__31144;
    wire N__31121;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31109;
    wire N__31108;
    wire N__31107;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31090;
    wire N__31087;
    wire N__31086;
    wire N__31085;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31061;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31045;
    wire N__31044;
    wire N__31041;
    wire N__31036;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31028;
    wire N__31027;
    wire N__31026;
    wire N__31025;
    wire N__31024;
    wire N__31021;
    wire N__31020;
    wire N__31019;
    wire N__31018;
    wire N__31017;
    wire N__31016;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__30998;
    wire N__30997;
    wire N__30996;
    wire N__30993;
    wire N__30988;
    wire N__30985;
    wire N__30984;
    wire N__30979;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30955;
    wire N__30952;
    wire N__30943;
    wire N__30940;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30882;
    wire N__30879;
    wire N__30874;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30858;
    wire N__30855;
    wire N__30854;
    wire N__30853;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30833;
    wire N__30832;
    wire N__30829;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30810;
    wire N__30809;
    wire N__30804;
    wire N__30801;
    wire N__30800;
    wire N__30799;
    wire N__30798;
    wire N__30797;
    wire N__30796;
    wire N__30795;
    wire N__30794;
    wire N__30791;
    wire N__30790;
    wire N__30787;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30742;
    wire N__30739;
    wire N__30730;
    wire N__30729;
    wire N__30724;
    wire N__30721;
    wire N__30716;
    wire N__30713;
    wire N__30712;
    wire N__30711;
    wire N__30710;
    wire N__30709;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30691;
    wire N__30688;
    wire N__30681;
    wire N__30676;
    wire N__30665;
    wire N__30664;
    wire N__30663;
    wire N__30662;
    wire N__30661;
    wire N__30660;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30644;
    wire N__30641;
    wire N__30640;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30632;
    wire N__30631;
    wire N__30630;
    wire N__30629;
    wire N__30626;
    wire N__30625;
    wire N__30622;
    wire N__30617;
    wire N__30616;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30591;
    wire N__30586;
    wire N__30581;
    wire N__30578;
    wire N__30577;
    wire N__30576;
    wire N__30575;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30561;
    wire N__30560;
    wire N__30559;
    wire N__30552;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30540;
    wire N__30539;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30503;
    wire N__30500;
    wire N__30495;
    wire N__30488;
    wire N__30467;
    wire N__30466;
    wire N__30465;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30424;
    wire N__30421;
    wire N__30420;
    wire N__30419;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30401;
    wire N__30400;
    wire N__30397;
    wire N__30396;
    wire N__30395;
    wire N__30394;
    wire N__30391;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30364;
    wire N__30359;
    wire N__30358;
    wire N__30355;
    wire N__30350;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30332;
    wire N__30329;
    wire N__30324;
    wire N__30311;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30299;
    wire N__30296;
    wire N__30295;
    wire N__30292;
    wire N__30291;
    wire N__30290;
    wire N__30289;
    wire N__30284;
    wire N__30283;
    wire N__30278;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30272;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30257;
    wire N__30252;
    wire N__30249;
    wire N__30246;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30224;
    wire N__30219;
    wire N__30206;
    wire N__30205;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30197;
    wire N__30196;
    wire N__30195;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30150;
    wire N__30141;
    wire N__30140;
    wire N__30135;
    wire N__30132;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30071;
    wire N__30070;
    wire N__30069;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30055;
    wire N__30054;
    wire N__30053;
    wire N__30052;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30034;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29961;
    wire N__29960;
    wire N__29959;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29945;
    wire N__29940;
    wire N__29939;
    wire N__29934;
    wire N__29929;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29908;
    wire N__29897;
    wire N__29894;
    wire N__29893;
    wire N__29890;
    wire N__29889;
    wire N__29888;
    wire N__29887;
    wire N__29886;
    wire N__29885;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29853;
    wire N__29850;
    wire N__29849;
    wire N__29848;
    wire N__29847;
    wire N__29846;
    wire N__29845;
    wire N__29844;
    wire N__29843;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29827;
    wire N__29820;
    wire N__29817;
    wire N__29812;
    wire N__29803;
    wire N__29798;
    wire N__29793;
    wire N__29790;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29703;
    wire N__29698;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29672;
    wire N__29669;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29653;
    wire N__29650;
    wire N__29645;
    wire N__29642;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29623;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29569;
    wire N__29568;
    wire N__29567;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29559;
    wire N__29556;
    wire N__29555;
    wire N__29552;
    wire N__29547;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29531;
    wire N__29530;
    wire N__29525;
    wire N__29522;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29510;
    wire N__29509;
    wire N__29508;
    wire N__29503;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29487;
    wire N__29478;
    wire N__29465;
    wire N__29462;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29453;
    wire N__29452;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29436;
    wire N__29435;
    wire N__29432;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29413;
    wire N__29412;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29406;
    wire N__29403;
    wire N__29402;
    wire N__29397;
    wire N__29390;
    wire N__29389;
    wire N__29386;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29370;
    wire N__29369;
    wire N__29368;
    wire N__29367;
    wire N__29364;
    wire N__29359;
    wire N__29352;
    wire N__29345;
    wire N__29338;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29314;
    wire N__29311;
    wire N__29310;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29298;
    wire N__29295;
    wire N__29294;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29263;
    wire N__29262;
    wire N__29261;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29247;
    wire N__29246;
    wire N__29245;
    wire N__29242;
    wire N__29241;
    wire N__29240;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29221;
    wire N__29216;
    wire N__29213;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29189;
    wire N__29188;
    wire N__29187;
    wire N__29186;
    wire N__29185;
    wire N__29182;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29131;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29123;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29115;
    wire N__29112;
    wire N__29103;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29012;
    wire N__29009;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28963;
    wire N__28962;
    wire N__28961;
    wire N__28958;
    wire N__28951;
    wire N__28948;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28932;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28927;
    wire N__28926;
    wire N__28925;
    wire N__28924;
    wire N__28923;
    wire N__28922;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28918;
    wire N__28917;
    wire N__28916;
    wire N__28915;
    wire N__28912;
    wire N__28905;
    wire N__28900;
    wire N__28893;
    wire N__28884;
    wire N__28875;
    wire N__28866;
    wire N__28859;
    wire N__28854;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28837;
    wire N__28834;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28817;
    wire N__28816;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28801;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28780;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28748;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28700;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28675;
    wire N__28674;
    wire N__28671;
    wire N__28666;
    wire N__28665;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28528;
    wire N__28527;
    wire N__28526;
    wire N__28525;
    wire N__28522;
    wire N__28515;
    wire N__28512;
    wire N__28511;
    wire N__28510;
    wire N__28509;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28495;
    wire N__28492;
    wire N__28491;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28463;
    wire N__28460;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28435;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28352;
    wire N__28349;
    wire N__28348;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28324;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28305;
    wire N__28304;
    wire N__28303;
    wire N__28302;
    wire N__28299;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28285;
    wire N__28284;
    wire N__28281;
    wire N__28280;
    wire N__28279;
    wire N__28278;
    wire N__28275;
    wire N__28274;
    wire N__28273;
    wire N__28272;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28251;
    wire N__28246;
    wire N__28241;
    wire N__28236;
    wire N__28233;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28201;
    wire N__28200;
    wire N__28199;
    wire N__28198;
    wire N__28195;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28183;
    wire N__28182;
    wire N__28181;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28171;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28163;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28151;
    wire N__28148;
    wire N__28141;
    wire N__28136;
    wire N__28131;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28087;
    wire N__28084;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27985;
    wire N__27982;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27944;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27910;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27895;
    wire N__27892;
    wire N__27891;
    wire N__27890;
    wire N__27887;
    wire N__27886;
    wire N__27883;
    wire N__27878;
    wire N__27875;
    wire N__27874;
    wire N__27873;
    wire N__27870;
    wire N__27869;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27854;
    wire N__27851;
    wire N__27846;
    wire N__27843;
    wire N__27838;
    wire N__27833;
    wire N__27830;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27807;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27799;
    wire N__27798;
    wire N__27797;
    wire N__27792;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27767;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27682;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27662;
    wire N__27661;
    wire N__27660;
    wire N__27657;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27647;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27629;
    wire N__27626;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27550;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27532;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27499;
    wire N__27494;
    wire N__27491;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27452;
    wire N__27449;
    wire N__27448;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27425;
    wire N__27422;
    wire N__27421;
    wire N__27420;
    wire N__27417;
    wire N__27416;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27389;
    wire N__27386;
    wire N__27381;
    wire N__27378;
    wire N__27373;
    wire N__27370;
    wire N__27365;
    wire N__27362;
    wire N__27353;
    wire N__27352;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27342;
    wire N__27341;
    wire N__27340;
    wire N__27339;
    wire N__27338;
    wire N__27333;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27321;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27289;
    wire N__27284;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27061;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27043;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27025;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26966;
    wire N__26965;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26893;
    wire N__26890;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26845;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26813;
    wire N__26812;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26764;
    wire N__26763;
    wire N__26758;
    wire N__26755;
    wire N__26750;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26728;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26692;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26672;
    wire N__26669;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26651;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26599;
    wire N__26594;
    wire N__26591;
    wire N__26590;
    wire N__26589;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26572;
    wire N__26571;
    wire N__26566;
    wire N__26563;
    wire N__26558;
    wire N__26557;
    wire N__26552;
    wire N__26549;
    wire N__26548;
    wire N__26543;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26531;
    wire N__26530;
    wire N__26529;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26510;
    wire N__26507;
    wire N__26506;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26488;
    wire N__26485;
    wire N__26480;
    wire N__26477;
    wire N__26476;
    wire N__26475;
    wire N__26472;
    wire N__26467;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26449;
    wire N__26444;
    wire N__26441;
    wire N__26440;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26416;
    wire N__26411;
    wire N__26408;
    wire N__26407;
    wire N__26406;
    wire N__26401;
    wire N__26398;
    wire N__26393;
    wire N__26392;
    wire N__26387;
    wire N__26384;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26328;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26285;
    wire N__26284;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26269;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26242;
    wire N__26239;
    wire N__26238;
    wire N__26237;
    wire N__26234;
    wire N__26233;
    wire N__26232;
    wire N__26229;
    wire N__26228;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26196;
    wire N__26193;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26137;
    wire N__26134;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26050;
    wire N__26047;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26035;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26020;
    wire N__26019;
    wire N__26012;
    wire N__26011;
    wire N__26010;
    wire N__26009;
    wire N__26008;
    wire N__26007;
    wire N__26006;
    wire N__26005;
    wire N__26002;
    wire N__25993;
    wire N__25990;
    wire N__25989;
    wire N__25988;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25967;
    wire N__25958;
    wire N__25949;
    wire N__25948;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25930;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25918;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25900;
    wire N__25899;
    wire N__25896;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25880;
    wire N__25877;
    wire N__25876;
    wire N__25875;
    wire N__25874;
    wire N__25873;
    wire N__25872;
    wire N__25871;
    wire N__25870;
    wire N__25869;
    wire N__25868;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25856;
    wire N__25853;
    wire N__25852;
    wire N__25849;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25837;
    wire N__25836;
    wire N__25835;
    wire N__25832;
    wire N__25823;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25806;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25732;
    wire N__25729;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25711;
    wire N__25710;
    wire N__25709;
    wire N__25708;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25696;
    wire N__25691;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25665;
    wire N__25664;
    wire N__25663;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25610;
    wire N__25607;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25577;
    wire N__25574;
    wire N__25573;
    wire N__25572;
    wire N__25571;
    wire N__25570;
    wire N__25567;
    wire N__25566;
    wire N__25563;
    wire N__25562;
    wire N__25561;
    wire N__25560;
    wire N__25557;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25548;
    wire N__25545;
    wire N__25544;
    wire N__25543;
    wire N__25542;
    wire N__25541;
    wire N__25540;
    wire N__25539;
    wire N__25538;
    wire N__25537;
    wire N__25536;
    wire N__25535;
    wire N__25534;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25512;
    wire N__25507;
    wire N__25498;
    wire N__25491;
    wire N__25484;
    wire N__25479;
    wire N__25470;
    wire N__25469;
    wire N__25468;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25452;
    wire N__25447;
    wire N__25438;
    wire N__25431;
    wire N__25428;
    wire N__25417;
    wire N__25412;
    wire N__25411;
    wire N__25410;
    wire N__25409;
    wire N__25408;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25401;
    wire N__25400;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25390;
    wire N__25387;
    wire N__25386;
    wire N__25385;
    wire N__25384;
    wire N__25381;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25373;
    wire N__25368;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25360;
    wire N__25351;
    wire N__25344;
    wire N__25335;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25311;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25300;
    wire N__25299;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25295;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25270;
    wire N__25267;
    wire N__25262;
    wire N__25255;
    wire N__25252;
    wire N__25247;
    wire N__25240;
    wire N__25231;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25174;
    wire N__25169;
    wire N__25166;
    wire N__25165;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25152;
    wire N__25147;
    wire N__25140;
    wire N__25137;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25107;
    wire N__25106;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25088;
    wire N__25085;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25036;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24976;
    wire N__24973;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24944;
    wire N__24941;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24924;
    wire N__24923;
    wire N__24922;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24891;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24844;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24752;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24740;
    wire N__24737;
    wire N__24736;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24718;
    wire N__24717;
    wire N__24714;
    wire N__24709;
    wire N__24706;
    wire N__24701;
    wire N__24698;
    wire N__24697;
    wire N__24696;
    wire N__24695;
    wire N__24694;
    wire N__24693;
    wire N__24692;
    wire N__24691;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24687;
    wire N__24684;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24676;
    wire N__24675;
    wire N__24670;
    wire N__24669;
    wire N__24668;
    wire N__24667;
    wire N__24666;
    wire N__24665;
    wire N__24664;
    wire N__24663;
    wire N__24662;
    wire N__24661;
    wire N__24656;
    wire N__24655;
    wire N__24654;
    wire N__24653;
    wire N__24650;
    wire N__24649;
    wire N__24648;
    wire N__24645;
    wire N__24644;
    wire N__24643;
    wire N__24642;
    wire N__24641;
    wire N__24640;
    wire N__24639;
    wire N__24632;
    wire N__24631;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24620;
    wire N__24617;
    wire N__24616;
    wire N__24615;
    wire N__24612;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24588;
    wire N__24581;
    wire N__24578;
    wire N__24565;
    wire N__24556;
    wire N__24555;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24506;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24486;
    wire N__24483;
    wire N__24476;
    wire N__24471;
    wire N__24466;
    wire N__24461;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24439;
    wire N__24434;
    wire N__24427;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24350;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24308;
    wire N__24307;
    wire N__24306;
    wire N__24305;
    wire N__24304;
    wire N__24303;
    wire N__24302;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24271;
    wire N__24268;
    wire N__24263;
    wire N__24262;
    wire N__24261;
    wire N__24260;
    wire N__24251;
    wire N__24248;
    wire N__24247;
    wire N__24246;
    wire N__24245;
    wire N__24244;
    wire N__24243;
    wire N__24242;
    wire N__24239;
    wire N__24226;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24197;
    wire N__24194;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24170;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24160;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24153;
    wire N__24152;
    wire N__24149;
    wire N__24148;
    wire N__24147;
    wire N__24146;
    wire N__24145;
    wire N__24144;
    wire N__24143;
    wire N__24142;
    wire N__24141;
    wire N__24140;
    wire N__24139;
    wire N__24138;
    wire N__24137;
    wire N__24136;
    wire N__24135;
    wire N__24134;
    wire N__24133;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24121;
    wire N__24114;
    wire N__24105;
    wire N__24096;
    wire N__24093;
    wire N__24084;
    wire N__24077;
    wire N__24068;
    wire N__24059;
    wire N__24054;
    wire N__24049;
    wire N__24048;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24037;
    wire N__24036;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23944;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23908;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23887;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23860;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23789;
    wire N__23784;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23761;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23650;
    wire N__23645;
    wire N__23642;
    wire N__23641;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23572;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23560;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23473;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23461;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23449;
    wire N__23448;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23409;
    wire N__23404;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23368;
    wire N__23363;
    wire N__23360;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23338;
    wire N__23333;
    wire N__23330;
    wire N__23329;
    wire N__23328;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23276;
    wire N__23273;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23246;
    wire N__23243;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23231;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23216;
    wire N__23213;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23201;
    wire N__23198;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23186;
    wire N__23183;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23171;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23163;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23148;
    wire N__23147;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23135;
    wire N__23134;
    wire N__23131;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23063;
    wire N__23060;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22933;
    wire N__22932;
    wire N__22927;
    wire N__22924;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22900;
    wire N__22899;
    wire N__22898;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22882;
    wire N__22877;
    wire N__22874;
    wire N__22873;
    wire N__22872;
    wire N__22871;
    wire N__22864;
    wire N__22861;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22843;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22801;
    wire N__22798;
    wire N__22797;
    wire N__22794;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22768;
    wire N__22763;
    wire N__22760;
    wire N__22759;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22532;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22490;
    wire N__22487;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22292;
    wire N__22289;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22240;
    wire N__22237;
    wire N__22236;
    wire N__22233;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22221;
    wire N__22218;
    wire N__22213;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22183;
    wire N__22180;
    wire N__22179;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22122;
    wire N__22121;
    wire N__22120;
    wire N__22117;
    wire N__22110;
    wire N__22107;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22054;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21958;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21928;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21887;
    wire N__21884;
    wire N__21883;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21866;
    wire N__21865;
    wire N__21862;
    wire N__21861;
    wire N__21854;
    wire N__21851;
    wire N__21850;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21716;
    wire N__21715;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21707;
    wire N__21706;
    wire N__21705;
    wire N__21704;
    wire N__21703;
    wire N__21702;
    wire N__21699;
    wire N__21698;
    wire N__21695;
    wire N__21694;
    wire N__21693;
    wire N__21682;
    wire N__21673;
    wire N__21670;
    wire N__21661;
    wire N__21652;
    wire N__21649;
    wire N__21648;
    wire N__21647;
    wire N__21646;
    wire N__21645;
    wire N__21644;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21632;
    wire N__21629;
    wire N__21624;
    wire N__21621;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21593;
    wire N__21584;
    wire N__21577;
    wire N__21574;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21548;
    wire N__21547;
    wire N__21546;
    wire N__21545;
    wire N__21544;
    wire N__21543;
    wire N__21542;
    wire N__21541;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21537;
    wire N__21536;
    wire N__21533;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21519;
    wire N__21518;
    wire N__21517;
    wire N__21516;
    wire N__21513;
    wire N__21504;
    wire N__21497;
    wire N__21492;
    wire N__21491;
    wire N__21490;
    wire N__21489;
    wire N__21488;
    wire N__21487;
    wire N__21486;
    wire N__21485;
    wire N__21484;
    wire N__21483;
    wire N__21482;
    wire N__21481;
    wire N__21480;
    wire N__21475;
    wire N__21466;
    wire N__21461;
    wire N__21456;
    wire N__21451;
    wire N__21440;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21414;
    wire N__21409;
    wire N__21402;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21374;
    wire N__21373;
    wire N__21372;
    wire N__21371;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21350;
    wire N__21349;
    wire N__21348;
    wire N__21345;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21337;
    wire N__21336;
    wire N__21329;
    wire N__21322;
    wire N__21317;
    wire N__21314;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21306;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21247;
    wire N__21246;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21053;
    wire N__21052;
    wire N__21051;
    wire N__21050;
    wire N__21049;
    wire N__21048;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21008;
    wire N__21005;
    wire N__21004;
    wire N__21001;
    wire N__21000;
    wire N__20999;
    wire N__20998;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20987;
    wire N__20986;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20970;
    wire N__20961;
    wire N__20958;
    wire N__20957;
    wire N__20954;
    wire N__20947;
    wire N__20936;
    wire N__20927;
    wire N__20924;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20899;
    wire N__20896;
    wire N__20895;
    wire N__20890;
    wire N__20885;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20865;
    wire N__20858;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20842;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20824;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20807;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20736;
    wire N__20733;
    wire N__20726;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20680;
    wire N__20677;
    wire N__20676;
    wire N__20673;
    wire N__20672;
    wire N__20669;
    wire N__20664;
    wire N__20661;
    wire N__20654;
    wire N__20651;
    wire N__20650;
    wire N__20647;
    wire N__20646;
    wire N__20643;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20590;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20561;
    wire N__20560;
    wire N__20559;
    wire N__20554;
    wire N__20551;
    wire N__20546;
    wire N__20543;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20535;
    wire N__20534;
    wire N__20527;
    wire N__20524;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20494;
    wire N__20489;
    wire N__20486;
    wire N__20485;
    wire N__20484;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20422;
    wire N__20421;
    wire N__20418;
    wire N__20417;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20329;
    wire N__20326;
    wire N__20325;
    wire N__20322;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20294;
    wire N__20287;
    wire N__20284;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20152;
    wire N__20149;
    wire N__20148;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20047;
    wire N__20046;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20039;
    wire N__20036;
    wire N__20035;
    wire N__20034;
    wire N__20031;
    wire N__20030;
    wire N__20029;
    wire N__20028;
    wire N__20027;
    wire N__20026;
    wire N__20025;
    wire N__20024;
    wire N__20023;
    wire N__20018;
    wire N__20013;
    wire N__20010;
    wire N__20009;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19989;
    wire N__19984;
    wire N__19981;
    wire N__19980;
    wire N__19979;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19961;
    wire N__19960;
    wire N__19959;
    wire N__19954;
    wire N__19953;
    wire N__19952;
    wire N__19949;
    wire N__19940;
    wire N__19935;
    wire N__19934;
    wire N__19931;
    wire N__19924;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19903;
    wire N__19900;
    wire N__19893;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19840;
    wire N__19835;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19823;
    wire N__19820;
    wire N__19819;
    wire N__19816;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19670;
    wire N__19669;
    wire N__19666;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19600;
    wire N__19599;
    wire N__19596;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19584;
    wire N__19581;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19561;
    wire N__19556;
    wire N__19553;
    wire N__19552;
    wire N__19547;
    wire N__19544;
    wire N__19543;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19492;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19471;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19456;
    wire N__19453;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19435;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19411;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19384;
    wire N__19379;
    wire N__19378;
    wire N__19377;
    wire N__19374;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19348;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19330;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19276;
    wire N__19273;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19246;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19226;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19218;
    wire N__19215;
    wire N__19210;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19192;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19176;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19172;
    wire N__19167;
    wire N__19164;
    wire N__19163;
    wire N__19162;
    wire N__19161;
    wire N__19160;
    wire N__19151;
    wire N__19148;
    wire N__19147;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19143;
    wire N__19142;
    wire N__19141;
    wire N__19138;
    wire N__19131;
    wire N__19128;
    wire N__19123;
    wire N__19114;
    wire N__19107;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19058;
    wire N__19057;
    wire N__19054;
    wire N__19047;
    wire N__19044;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19012;
    wire N__19011;
    wire N__19010;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18994;
    wire N__18991;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18971;
    wire N__18970;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18946;
    wire N__18945;
    wire N__18944;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18916;
    wire N__18915;
    wire N__18912;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18766;
    wire N__18763;
    wire N__18762;
    wire N__18755;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18732;
    wire N__18731;
    wire N__18730;
    wire N__18727;
    wire N__18720;
    wire N__18717;
    wire N__18710;
    wire N__18709;
    wire N__18706;
    wire N__18705;
    wire N__18698;
    wire N__18695;
    wire N__18694;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18683;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18671;
    wire N__18668;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18622;
    wire N__18619;
    wire N__18618;
    wire N__18611;
    wire N__18608;
    wire N__18607;
    wire N__18604;
    wire N__18603;
    wire N__18596;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18584;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18572;
    wire N__18571;
    wire N__18568;
    wire N__18567;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18476;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18464;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18449;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18346;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18314;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18302;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18287;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18275;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18263;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18236;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18224;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18212;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18200;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18185;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18173;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18162;
    wire N__18161;
    wire N__18156;
    wire N__18151;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18125;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18104;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18092;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18080;
    wire N__18079;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18065;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18034;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17989;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17977;
    wire N__17974;
    wire N__17973;
    wire N__17970;
    wire N__17965;
    wire N__17960;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17948;
    wire N__17947;
    wire N__17944;
    wire N__17943;
    wire N__17940;
    wire N__17935;
    wire N__17930;
    wire N__17929;
    wire N__17928;
    wire N__17925;
    wire N__17920;
    wire N__17915;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17900;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17866;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17773;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17761;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17735;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17716;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17671;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17629;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17614;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17588;
    wire N__17585;
    wire N__17584;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17482;
    wire N__17479;
    wire N__17478;
    wire N__17475;
    wire N__17470;
    wire N__17465;
    wire N__17462;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17444;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17423;
    wire N__17422;
    wire N__17421;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17365;
    wire N__17362;
    wire N__17361;
    wire N__17360;
    wire N__17351;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17317;
    wire N__17314;
    wire N__17313;
    wire N__17310;
    wire N__17309;
    wire N__17308;
    wire N__17305;
    wire N__17298;
    wire N__17295;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17249;
    wire N__17246;
    wire N__17245;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17233;
    wire N__17232;
    wire N__17229;
    wire N__17224;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17137;
    wire N__17134;
    wire N__17133;
    wire N__17130;
    wire N__17129;
    wire N__17128;
    wire N__17125;
    wire N__17118;
    wire N__17115;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17079;
    wire N__17078;
    wire N__17077;
    wire N__17074;
    wire N__17067;
    wire N__17064;
    wire N__17057;
    wire N__17054;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17046;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17034;
    wire N__17031;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16933;
    wire N__16928;
    wire N__16925;
    wire N__16924;
    wire N__16919;
    wire N__16916;
    wire N__16915;
    wire N__16912;
    wire N__16907;
    wire N__16904;
    wire N__16903;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16771;
    wire N__16770;
    wire N__16769;
    wire N__16768;
    wire N__16765;
    wire N__16756;
    wire N__16751;
    wire N__16750;
    wire N__16745;
    wire N__16742;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16734;
    wire N__16733;
    wire N__16732;
    wire N__16731;
    wire N__16728;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16699;
    wire N__16698;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16686;
    wire N__16679;
    wire N__16678;
    wire N__16677;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16637;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16613;
    wire N__16610;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16531;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16513;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16469;
    wire N__16466;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16454;
    wire N__16451;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16439;
    wire N__16436;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16421;
    wire N__16418;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16403;
    wire N__16400;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16388;
    wire N__16385;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16366;
    wire N__16365;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16352;
    wire N__16349;
    wire N__16344;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16310;
    wire N__16307;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16295;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16280;
    wire N__16277;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16265;
    wire N__16262;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16250;
    wire N__16247;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16235;
    wire N__16232;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16205;
    wire N__16202;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16171;
    wire N__16170;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16156;
    wire N__16155;
    wire N__16150;
    wire N__16147;
    wire N__16142;
    wire N__16139;
    wire N__16138;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16084;
    wire N__16081;
    wire N__16080;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15991;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15931;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15865;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15831;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15819;
    wire N__15812;
    wire N__15811;
    wire N__15806;
    wire N__15805;
    wire N__15804;
    wire N__15803;
    wire N__15802;
    wire N__15801;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15797;
    wire N__15796;
    wire N__15795;
    wire N__15794;
    wire N__15793;
    wire N__15792;
    wire N__15789;
    wire N__15784;
    wire N__15781;
    wire N__15780;
    wire N__15777;
    wire N__15770;
    wire N__15763;
    wire N__15754;
    wire N__15747;
    wire N__15744;
    wire N__15731;
    wire N__15730;
    wire N__15729;
    wire N__15728;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15707;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15689;
    wire N__15686;
    wire N__15685;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15614;
    wire N__15613;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15593;
    wire N__15592;
    wire N__15591;
    wire N__15584;
    wire N__15581;
    wire N__15580;
    wire N__15575;
    wire N__15572;
    wire N__15571;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15496;
    wire N__15495;
    wire N__15492;
    wire N__15487;
    wire N__15482;
    wire N__15481;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15463;
    wire N__15462;
    wire N__15455;
    wire N__15452;
    wire N__15451;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15394;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15377;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15365;
    wire N__15362;
    wire N__15361;
    wire N__15360;
    wire N__15357;
    wire N__15352;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15333;
    wire N__15330;
    wire N__15329;
    wire N__15326;
    wire N__15321;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15289;
    wire N__15284;
    wire N__15281;
    wire N__15272;
    wire N__15271;
    wire N__15270;
    wire N__15267;
    wire N__15266;
    wire N__15263;
    wire N__15262;
    wire N__15261;
    wire N__15260;
    wire N__15259;
    wire N__15258;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15236;
    wire N__15233;
    wire N__15224;
    wire N__15221;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15209;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15187;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15170;
    wire N__15167;
    wire N__15166;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15145;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15129;
    wire N__15124;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15080;
    wire N__15077;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15065;
    wire N__15062;
    wire N__15061;
    wire N__15060;
    wire N__15057;
    wire N__15052;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14992;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14951;
    wire N__14948;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14936;
    wire N__14933;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14896;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14878;
    wire N__14873;
    wire N__14870;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14858;
    wire N__14855;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14840;
    wire N__14837;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14801;
    wire N__14798;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14783;
    wire N__14780;
    wire N__14779;
    wire N__14776;
    wire N__14775;
    wire N__14770;
    wire N__14767;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14734;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14701;
    wire N__14698;
    wire N__14697;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14662;
    wire N__14659;
    wire N__14658;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14620;
    wire N__14617;
    wire N__14616;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14508;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14449;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14437;
    wire N__14436;
    wire N__14433;
    wire N__14428;
    wire N__14423;
    wire N__14422;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14368;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14339;
    wire N__14338;
    wire N__14335;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14323;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14299;
    wire N__14298;
    wire N__14295;
    wire N__14290;
    wire N__14285;
    wire N__14284;
    wire N__14281;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14252;
    wire N__14251;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14209;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14174;
    wire N__14173;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14083;
    wire N__14082;
    wire N__14081;
    wire N__14080;
    wire N__14069;
    wire N__14066;
    wire N__14065;
    wire N__14064;
    wire N__14063;
    wire N__14060;
    wire N__14059;
    wire N__14056;
    wire N__14047;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire VCCG0;
    wire N_428_cascade_;
    wire \PCH_PWRGD.delayed_vccin_okZ0 ;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.m14_i_0 ;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_ ;
    wire hda_sdo_atp;
    wire \HDA_STRAP.N_16_cascade_ ;
    wire \HDA_STRAP.HDA_SDO_ATP_3_0 ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire \HDA_STRAP.un4_count_9_cascade_ ;
    wire \HDA_STRAP.un4_count_12 ;
    wire \HDA_STRAP.un4_count_11 ;
    wire \HDA_STRAP.un4_count_13_cascade_ ;
    wire \HDA_STRAP.un4_count_10 ;
    wire \HDA_STRAP.un4_count_cascade_ ;
    wire \PCH_PWRGD.count_rst_5 ;
    wire \PCH_PWRGD.count_rst_5_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_9_cascade_ ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_8_cascade_ ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.count_rst_9_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_5_cascade_ ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.count_rst_10_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_4_cascade_ ;
    wire \PCH_PWRGD.count_rst_10 ;
    wire \PCH_PWRGD.count_0_4 ;
    wire bfn_1_6_0_;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.un2_count_1_axb_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.countZ0Z_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire \PCH_PWRGD.un2_count_1_axb_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire bfn_1_7_0_;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.un2_count_1_axb_13 ;
    wire \PCH_PWRGD.count_0_15 ;
    wire \PCH_PWRGD.count_rst ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \PCH_PWRGD.countZ0Z_15_cascade_ ;
    wire \PCH_PWRGD.count_rst_1 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.count_0_12 ;
    wire bfn_1_9_0_;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire bfn_1_10_0_;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire bfn_1_11_0_;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire bfn_1_12_0_;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \POWERLED.g1_i_a4_0_1_cascade_ ;
    wire \POWERLED.N_12 ;
    wire \POWERLED.N_5_cascade_ ;
    wire \POWERLED.pwm_out_en_cascade_ ;
    wire pwrbtn_led;
    wire \POWERLED.N_11 ;
    wire \POWERLED.g0_2_1 ;
    wire \POWERLED.pwm_outZ0 ;
    wire \POWERLED.N_2360_i_cascade_ ;
    wire \VPP_VDDQ.un6_count_11_cascade_ ;
    wire \VPP_VDDQ.un6_count_9 ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \VPP_VDDQ.un6_count_8 ;
    wire vpp_ok;
    wire vddq_en;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire bfn_2_1_0_;
    wire \HDA_STRAP.countZ0Z_1 ;
    wire \HDA_STRAP.un1_count_1_cry_0 ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.un1_count_1_cry_1 ;
    wire \HDA_STRAP.countZ0Z_3 ;
    wire \HDA_STRAP.un1_count_1_cry_2 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.un1_count_1_cry_3 ;
    wire \HDA_STRAP.countZ0Z_5 ;
    wire \HDA_STRAP.un1_count_1_cry_4 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.un1_count_1_cry_5_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_5 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un1_count_1_cry_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7 ;
    wire \HDA_STRAP.countZ0Z_8 ;
    wire \HDA_STRAP.un1_count_1_cry_7_THRU_CO ;
    wire bfn_2_2_0_;
    wire \HDA_STRAP.countZ0Z_9 ;
    wire \HDA_STRAP.un1_count_1_cry_8 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.un1_count_1_cry_9_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_9 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.un1_count_1_cry_10_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_10 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.un1_count_1_cry_11 ;
    wire \HDA_STRAP.countZ0Z_13 ;
    wire \HDA_STRAP.un1_count_1_cry_12 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.un1_count_1_cry_13 ;
    wire \HDA_STRAP.countZ0Z_15 ;
    wire \HDA_STRAP.un1_count_1_cry_14 ;
    wire \HDA_STRAP.un1_count_1_cry_15 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.un1_count_1_cry_15_THRU_CO ;
    wire bfn_2_3_0_;
    wire \HDA_STRAP.curr_state_RNIH91AZ0Z_0 ;
    wire \HDA_STRAP.un4_count ;
    wire \HDA_STRAP.un1_count_1_cry_16 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.count_rst_7_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.count_rst_7 ;
    wire \PCH_PWRGD.count_0_7 ;
    wire \PCH_PWRGD.un2_count_1_axb_7 ;
    wire \PCH_PWRGD.count_rst_3 ;
    wire \PCH_PWRGD.count_0_11 ;
    wire \PCH_PWRGD.countZ0Z_11 ;
    wire \PCH_PWRGD.countZ0Z_11_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_4_0 ;
    wire \PCH_PWRGD.count_1_i_a2_5_0 ;
    wire \PCH_PWRGD.count_1_i_a2_3_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_6_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_2226_i_cascade_ ;
    wire \PCH_PWRGD.curr_state_7_0 ;
    wire \PCH_PWRGD.N_386_cascade_ ;
    wire \PCH_PWRGD.count_rst_11_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_3_cascade_ ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.countZ0Z_14_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.count_1_i_a2_1_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_2_0 ;
    wire \PCH_PWRGD.count_1_i_a2_11_0 ;
    wire \PCH_PWRGD.count_1_i_a2_11_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_12_0 ;
    wire \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.count_rst_12 ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.un2_count_1_axb_2 ;
    wire \PCH_PWRGD.count_rst_14 ;
    wire \PCH_PWRGD.count_0_0 ;
    wire \PCH_PWRGD.count_0_sqmuxa_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.countZ0Z_6_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_0_0 ;
    wire \PCH_PWRGD.un2_count_1_axb_1_cascade_ ;
    wire \PCH_PWRGD.count_rst_13 ;
    wire \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.un2_count_1_axb_10 ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.curr_state_0_0 ;
    wire \PCH_PWRGD.N_2244_i ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.N_2244_i_cascade_ ;
    wire \PCH_PWRGD.N_655_cascade_ ;
    wire \PCH_PWRGD.m6_i_i_a2 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.N_386 ;
    wire \PCH_PWRGD.N_2226_i ;
    wire \PCH_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.N_655 ;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire N_626_cascade_;
    wire \POWERLED.G_30Z0Z_0_cascade_ ;
    wire VPP_VDDQ_un6_count;
    wire G_30_cascade_;
    wire bfn_2_10_0_;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_axb_4_l_fx ;
    wire bfn_2_11_0_;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire bfn_2_12_0_;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.count_1_5_cascade_ ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.count_1_5 ;
    wire \POWERLED.un79_clk_100khzlto6_0_cascade_ ;
    wire \POWERLED.un79_clk_100khz ;
    wire \POWERLED.un79_clk_100khz_cascade_ ;
    wire \POWERLED.N_2360_i ;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \VPP_VDDQ.N_64_i ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire bfn_2_14_0_;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire bfn_2_15_0_;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_2_16_0_;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.N_92_0 ;
    wire G_30;
    wire \VPP_VDDQ.count_2_1_8_cascade_ ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.count_2_1_9_cascade_ ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.count_2_1_14_cascade_ ;
    wire \VPP_VDDQ.count_2_1_4_cascade_ ;
    wire \VPP_VDDQ.count_2_0_4 ;
    wire \VPP_VDDQ.count_2_0_5 ;
    wire \VPP_VDDQ.count_2_1_5_cascade_ ;
    wire \VPP_VDDQ.count_2_1_12_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_12_cascade_ ;
    wire \VPP_VDDQ.count_2_0_12 ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.count_2_0_14 ;
    wire VPP_VDDQ_curr_state_0;
    wire VPP_VDDQ_curr_state_1;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ;
    wire N_626;
    wire \PCH_PWRGD.curr_state_0_sqmuxa ;
    wire \PCH_PWRGD.N_38_f0 ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \VPP_VDDQ.count_2_0_10 ;
    wire \VPP_VDDQ.count_2_1_10_cascade_ ;
    wire bfn_4_5_0_;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_4_6_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_4_7_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_4_8_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \POWERLED.N_4842_i ;
    wire bfn_4_9_0_;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.count_i_3 ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.count_RNIGTVS_1Z0Z_5 ;
    wire \POWERLED.mult1_un131_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.count_i_6 ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.N_4841_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.count_i_8 ;
    wire bfn_4_10_0_;
    wire \POWERLED.N_4849_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.count_i_10 ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.count_i_11 ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.N_4851_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.N_4855_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.N_4856_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_4_11_0_;
    wire \POWERLED.mult1_un117_sum_i_8 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_i_8 ;
    wire \POWERLED.mult1_un89_sum_i_8 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_i_8 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_i_8 ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.N_437_cascade_ ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.curr_stateZ0Z_0_cascade_ ;
    wire \POWERLED.curr_state_1_0 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.mult1_un152_sum_i_8 ;
    wire \POWERLED.count_RNIAKSS_0Z0Z_2 ;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.un79_clk_100khzlto4_0_cascade_ ;
    wire \POWERLED.un79_clk_100khzlt6 ;
    wire \POWERLED.mult1_un138_sum_i_8 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.count_RNIJEFE_0Z0Z_4 ;
    wire \POWERLED.mult1_un159_sum_i_8 ;
    wire \POWERLED.count_RNIUGSJ_0Z0Z_1 ;
    wire \POWERLED.N_660 ;
    wire \POWERLED.count_0_sqmuxa_cascade_ ;
    wire \POWERLED.count_1_0_cascade_ ;
    wire \POWERLED.countZ0Z_0_cascade_ ;
    wire \POWERLED.count_1_1 ;
    wire \POWERLED.count_1_1_cascade_ ;
    wire \POWERLED.un1_count_axb_1_cascade_ ;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.count_0_0 ;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.countZ0Z_14_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_5 ;
    wire \POWERLED.g1_i_o4_4 ;
    wire \POWERLED.count_0_15 ;
    wire \VPP_VDDQ.count_2_0_2 ;
    wire \VPP_VDDQ.count_2_1_2_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_2_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire bfn_5_2_0_;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ;
    wire bfn_5_3_0_;
    wire \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ;
    wire \VPP_VDDQ.count_2_1_13 ;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire \VPP_VDDQ.un9_clk_100khz_10 ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.un9_clk_100khz_7 ;
    wire \VPP_VDDQ.count_2_1_7 ;
    wire \VPP_VDDQ.count_2_1_7_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.count_2_1_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \PCH_PWRGD.N_670 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire bfn_5_8_0_;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire vccst_en;
    wire G_12;
    wire \POWERLED.mult1_un68_sum_i_8 ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un124_sum_i_8 ;
    wire bfn_5_11_0_;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire bfn_5_12_0_;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.un1_count_axb_1 ;
    wire bfn_5_13_0_;
    wire \POWERLED.un1_count_axb_2 ;
    wire \POWERLED.count_1_2 ;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.un1_count_cry_2_c_RNICZ0Z419 ;
    wire \POWERLED.un1_count_cry_2 ;
    wire \POWERLED.un1_count_axb_4 ;
    wire \POWERLED.count_1_4 ;
    wire \POWERLED.un1_count_cry_3 ;
    wire \POWERLED.un1_count_axb_5 ;
    wire \POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ;
    wire \POWERLED.un1_count_cry_4 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire bfn_5_14_0_;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.count_1_11 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.un1_count_cry_11 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.count_1_14 ;
    wire \POWERLED.un1_count_cry_13 ;
    wire \POWERLED.count_0_sqmuxa ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ;
    wire \POWERLED.un1_count_axb_12 ;
    wire \POWERLED.count_1_9 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.count_1_10 ;
    wire \POWERLED.count_0_10 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.count_1_6 ;
    wire \POWERLED.count_0_6 ;
    wire \POWERLED.count_1_8 ;
    wire \POWERLED.count_0_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire \VPP_VDDQ.count_2_1_3_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.delayed_vddq_okZ0 ;
    wire VPP_VDDQ_delayed_vddq_ok_cascade_;
    wire vccst_pwrgd;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \VPP_VDDQ.un9_clk_100khz_9 ;
    wire \VPP_VDDQ.un9_clk_100khz_0_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ;
    wire \VPP_VDDQ.N_1_i_cascade_ ;
    wire \VPP_VDDQ.count_2_1_6 ;
    wire \VPP_VDDQ.count_2_1_6_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_6 ;
    wire v1p8a_ok;
    wire v5a_ok;
    wire v33a_ok;
    wire slp_susn;
    wire v33a_enn;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2_1_1_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1 ;
    wire \VPP_VDDQ.count_2_1_1 ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.un9_clk_100khz_1 ;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1 ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ;
    wire \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ;
    wire \VPP_VDDQ.count_2_1_11_cascade_ ;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire \VPP_VDDQ.N_60_i ;
    wire \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.N_60 ;
    wire \VPP_VDDQ.N_60_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_ok_en ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_6_5_0_;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire COUNTER_un4_counter_7;
    wire bfn_6_6_0_;
    wire bfn_6_7_0_;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_2161;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.mult1_un166_sum_i_8 ;
    wire \POWERLED.mult1_un145_sum_i_8 ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire bfn_6_10_0_;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un75_sum_i_8 ;
    wire bfn_6_11_0_;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire bfn_6_12_0_;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un82_sum_i_8 ;
    wire \POWERLED.count_RNICOIT_0Z0Z_12 ;
    wire \POWERLED.count_0_13 ;
    wire \POWERLED.count_1_13 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.countZ0Z_13_cascade_ ;
    wire \POWERLED.count_1_12 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.un79_clk_100khzlto15_3_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_6 ;
    wire \POWERLED.un79_clk_100khzlto15_3 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.g1_i_o4_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.count_1_7 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.N_6 ;
    wire \POWERLED.count_clk_0_6 ;
    wire bfn_6_15_0_;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire \VPP_VDDQ.N_53_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1 ;
    wire \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.N_664_cascade_ ;
    wire \VPP_VDDQ.m4_0_0_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire \VPP_VDDQ.curr_state_2_RNIZ0Z_1 ;
    wire vddq_ok;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.N_664 ;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire \VPP_VDDQ.N_53 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire N_557_g;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_ ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10 ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12_cascade_ ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9 ;
    wire bfn_7_3_0_;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire \POWERLED.dutycycleZ0Z_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_3_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_3_cascade_ ;
    wire \POWERLED.dutycycle_cascade_ ;
    wire \POWERLED.dutycycle_1_0_0 ;
    wire \POWERLED.dutycycle_1_0_0_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.dutycycle_1_0_1_cascade_ ;
    wire dutycycle_RNII6848_0_1_cascade_;
    wire \POWERLED.dutycycle_eena_0 ;
    wire \POWERLED.dutycycle_1_0_1 ;
    wire \POWERLED.dutycycle_eena_0_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.N_15 ;
    wire \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_ ;
    wire \POWERLED.N_672_cascade_ ;
    wire dutycycle_RNI_1_5;
    wire POWERLED_un1_dutycycle_172_m1;
    wire dutycycle_RNI_3_1_cascade_;
    wire bfn_7_7_0_;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.un1_dutycycle_53_axb_4_1 ;
    wire \POWERLED.g0_7_a2_2 ;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_0 ;
    wire \POWERLED.un2_count_clk_17_0_0_a2_0_4_cascade_ ;
    wire \POWERLED.N_604 ;
    wire \POWERLED.func_state_RNI1O2V5Z0Z_1 ;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.N_9_i_1_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_8_cascade_ ;
    wire \POWERLED.un1_clk_100khz_32_and_i_0_a2_0_0_0 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_6_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_0_a2_0_3 ;
    wire \POWERLED.un1_dutycycle_53_axb_0 ;
    wire bfn_7_11_0_;
    wire \POWERLED.dutycycle_RNI_2Z0Z_0 ;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_2 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_1 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_2 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_2 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_3 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_3 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_3 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_4 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_5 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_6 ;
    wire \POWERLED.un1_dutycycle_53_cry_7 ;
    wire \POWERLED.dutycycle_RNIZ0Z_11 ;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_7_12_0_;
    wire \POWERLED.dutycycle_RNIZ0Z_12 ;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_9 ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire bfn_7_13_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.un1_dutycycle_53_i_28 ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_14 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ;
    wire bfn_7_15_0_;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_axb_4 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_5 ;
    wire \POWERLED.mult1_un47_sum_cry_6_s ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire bfn_8_1_0_;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire bfn_8_2_0_;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_3_0_;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \POWERLED.N_413_N_cascade_ ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.N_413_N ;
    wire \POWERLED.N_430_cascade_ ;
    wire \POWERLED.dutycycle_eena_1 ;
    wire SUSWARN_N_fast;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m0 ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m1_ns_1_cascade_ ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m1 ;
    wire \COUNTER.tmp_0_fast_RNI0RLUZ0Z1 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_10Z0Z_0_cascade_ ;
    wire \POWERLED.N_676_cascade_ ;
    wire G_11_i_a10_0_1_cascade_;
    wire G_11_i_2;
    wire N_9_2_cascade_;
    wire N_8_3;
    wire G_11_i_a10_0_1;
    wire N_8_3_cascade_;
    wire \POWERLED.N_10_1 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_1 ;
    wire \POWERLED.dutycycle_0_5 ;
    wire \POWERLED.g0_i_o4_2 ;
    wire \POWERLED.dutycycleZ1Z_5_cascade_ ;
    wire \POWERLED.N_546 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_5 ;
    wire \POWERLED.N_612 ;
    wire N_16_0;
    wire \POWERLED.g0_0_1 ;
    wire \POWERLED.N_598_cascade_ ;
    wire \POWERLED.N_450_cascade_ ;
    wire \POWERLED.dutycycle_RNI5FJ65Z0Z_13 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.dutycycle_RNI5FJ65Z0Z_13_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_11_cascade_ ;
    wire \POWERLED.N_2336_i ;
    wire \POWERLED.N_449 ;
    wire \POWERLED.un1_m2_e_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.dutycycleZ0Z_7_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_56_a1_2_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_8 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \POWERLED.dutycycle_RNIT70K5Z0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_8_cascade_ ;
    wire \POWERLED.N_6_3_cascade_ ;
    wire \POWERLED.g0_9_1_0 ;
    wire \POWERLED.N_9_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_15Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_15 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_10 ;
    wire \POWERLED.N_4_0 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_13 ;
    wire \POWERLED.un1_dutycycle_53_12_1_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_6 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_8 ;
    wire \POWERLED.dutycycleZ1Z_14 ;
    wire \POWERLED.dutycycleZ0Z_10_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_13 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_15 ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.N_492 ;
    wire \POWERLED.count_clk_en_cascade_ ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.count_clk_0_4 ;
    wire bfn_8_15_0_;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_7_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire bfn_8_16_0_;
    wire \POWERLED.un1_count_clk_2_axb_10 ;
    wire \POWERLED.un1_count_clk_2_cry_9_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_10 ;
    wire \POWERLED.un1_count_clk_2_cry_11 ;
    wire \POWERLED.count_clk_1_13 ;
    wire \POWERLED.un1_count_clk_2_cry_12_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_13 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.count_clk_1_15 ;
    wire \POWERLED.un1_count_clk_2_axb_14 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11 ;
    wire \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ;
    wire \RSMRST_PWRGD.N_264_i ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0 ;
    wire \RSMRST_PWRGD.N_662 ;
    wire \RSMRST_PWRGD.N_555_cascade_ ;
    wire \RSMRST_PWRGD.G_14 ;
    wire N_92_g;
    wire \RSMRST_PWRGD.G_14_cascade_ ;
    wire \RSMRST_PWRGD.N_92_1 ;
    wire \POWERLED.N_423_0_cascade_ ;
    wire \POWERLED.g1_cascade_ ;
    wire \POWERLED.g0_0_0 ;
    wire \POWERLED.N_8_0_0 ;
    wire \POWERLED.g0_0_2_cascade_ ;
    wire \POWERLED.N_541_cascade_ ;
    wire \POWERLED.N_542 ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \POWERLED.g2 ;
    wire \POWERLED.g0_0_5 ;
    wire \POWERLED.g2_0 ;
    wire \POWERLED.g2_cascade_ ;
    wire \POWERLED.N_13_0_0_0 ;
    wire \POWERLED.func_stateZ0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_0 ;
    wire suswarn_n;
    wire \POWERLED.N_8_0_cascade_ ;
    wire \POWERLED.N_16_2 ;
    wire \POWERLED.dutycycle_e_N_3L4_0_1_cascade_ ;
    wire \POWERLED.g0_8Z0Z_0 ;
    wire \POWERLED.N_435_cascade_ ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_0 ;
    wire \POWERLED.func_state_1_m2s2_i_0_0 ;
    wire \POWERLED.N_423_cascade_ ;
    wire \POWERLED.dutycycle_RNI_10Z0Z_0 ;
    wire \POWERLED.N_613 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_3_1_cascade_ ;
    wire \POWERLED.N_252_N ;
    wire \POWERLED.dutycycle_eena_13_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_13_cascade_ ;
    wire \POWERLED.N_452 ;
    wire \POWERLED.dutycycle_set_1 ;
    wire \POWERLED.func_state_RNI12ASZ0Z_1 ;
    wire \POWERLED.func_state_RNI12ASZ0Z_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3 ;
    wire \POWERLED.dutycycle_eena_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3_cascade_ ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.dutycycle_RNI_13Z0Z_0 ;
    wire \POWERLED.N_2363_0_cascade_ ;
    wire \POWERLED.N_12_3_0 ;
    wire G_11_i_a10_2_1_cascade_;
    wire \POWERLED.g2_3 ;
    wire N_28;
    wire N_7;
    wire N_50;
    wire N_7_cascade_;
    wire \POWERLED.N_2363_0 ;
    wire \POWERLED.g1_0_1_cascade_ ;
    wire N_43;
    wire \POWERLED.g2_1 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire \PCH_PWRGD.un2_count_1_axb_1 ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0 ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_axb_7_l_fx ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire N_428;
    wire pch_pwrok;
    wire bfn_9_9_0_;
    wire dutycycle_RNII6848_0_1;
    wire \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ;
    wire bfn_9_10_0_;
    wire \POWERLED.un1_dutycycle_94_cry_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_cZ0 ;
    wire \POWERLED.N_435_i ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ;
    wire \POWERLED.un1_dutycycle_53_2_1 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_11 ;
    wire \POWERLED.un1_dutycycle_53_59_a0_0 ;
    wire \POWERLED.dutycycleZ1Z_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_56_a1_2 ;
    wire \POWERLED.un1_dutycycle_53_8_2 ;
    wire \POWERLED.un1_dutycycle_53_8_0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.G_7_i_a5_1_1_cascade_ ;
    wire \POWERLED.N_11_1 ;
    wire \POWERLED.N_16_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_2_cascade_ ;
    wire \POWERLED.g0_9_1 ;
    wire \POWERLED.g0_9_1_1_0 ;
    wire \POWERLED.dutycycle_RNIHDMC5Z0Z_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \POWERLED.dutycycle_RNI6SKJ1Z0Z_9 ;
    wire \POWERLED.dutycycle_RNIHDMC5Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.un1_dutycycle_53_7_0 ;
    wire \POWERLED.un1_dutycycle_53_41_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_13 ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ;
    wire \POWERLED.dutycycle_RNIHDMC5Z0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \POWERLED.N_17_cascade_ ;
    wire \POWERLED.N_8_2 ;
    wire \POWERLED.G_7_i_0 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.count_clkZ0Z_3_cascade_ ;
    wire \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.N_625 ;
    wire \POWERLED.N_625_cascade_ ;
    wire \POWERLED.count_clkZ0Z_9_cascade_ ;
    wire \POWERLED.count_clk_RNINSEUC_0Z0Z_10 ;
    wire \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ;
    wire \POWERLED.count_clk_0_9 ;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.count_clkZ0Z_7_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.count_clk_0_7 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.count_clk_1_10 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_0 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_2_cascade_ ;
    wire \POWERLED.count_clk_RNINSEUCZ0Z_10 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_1 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.count_clk_1_12 ;
    wire \POWERLED.un1_count_clk_2_axb_12 ;
    wire \POWERLED.count_clk_1_14 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.count_off_0_9 ;
    wire \POWERLED.count_offZ0Z_9_cascade_ ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_off_0_12 ;
    wire bfn_11_3_0_;
    wire \POWERLED.un3_count_off_1_cry_1 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_off_1_9 ;
    wire bfn_11_4_0_;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_off_1_10 ;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.count_off_1_12 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.N_627 ;
    wire \POWERLED.N_688 ;
    wire \POWERLED.N_74 ;
    wire \POWERLED.N_6_1_cascade_ ;
    wire \POWERLED.func_state_1_m2_1_cascade_ ;
    wire \POWERLED.func_state_cascade_ ;
    wire \POWERLED.N_426_i ;
    wire \POWERLED.N_562 ;
    wire \POWERLED.func_state_enZ0 ;
    wire \POWERLED.func_state_1_m2_1 ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ;
    wire \POWERLED.count_off_0_3 ;
    wire \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_offZ0Z_3_cascade_ ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.un34_clk_100khz_11 ;
    wire \POWERLED.un34_clk_100khz_8_cascade_ ;
    wire \POWERLED.count_off_RNI_0Z0Z_10_cascade_ ;
    wire \POWERLED.count_off_RNI8AQHZ0Z_10_cascade_ ;
    wire \POWERLED.func_state_1_m2_ns_1_1 ;
    wire \POWERLED.N_494 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ;
    wire \POWERLED.dutycycle_1_0_iv_i_i_m2_1_6_cascade_ ;
    wire \POWERLED.N_453 ;
    wire \POWERLED.N_133 ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0 ;
    wire \POWERLED.N_490 ;
    wire \POWERLED.g1_0_2 ;
    wire \POWERLED.func_state_RNI2MQDZ0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_eena_13_1_0 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6 ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_a2_d ;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ;
    wire \POWERLED.dutycycle_e_1_4 ;
    wire \POWERLED.dutycycle_e_1_4_cascade_ ;
    wire \POWERLED.func_state_RNIJ17U4Z0Z_1 ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ;
    wire \POWERLED.dutycycle_e_1_7 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.dutycycle_e_1_7_cascade_ ;
    wire \POWERLED.func_state_RNI9S7D5Z0Z_1 ;
    wire \POWERLED.dutycycleZ1Z_6_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_25_0_tz_1_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_4 ;
    wire \POWERLED.func_state_RNI_0Z0Z_1 ;
    wire \POWERLED.func_state_RNI2MQDZ0Z_1 ;
    wire \POWERLED.func_state_RNI2MQDZ0Z_1_cascade_ ;
    wire \POWERLED.func_state_RNI_8Z0Z_1_cascade_ ;
    wire \POWERLED.func_state_RNIMQ0F_0Z0Z_1 ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d ;
    wire \POWERLED.func_state_RNIMQ0F_0Z0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI2MQDZ0Z_7 ;
    wire \POWERLED.dutycycle_RNIEBSB1Z0Z_7 ;
    wire \POWERLED.N_545 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ;
    wire \POWERLED.N_71 ;
    wire \POWERLED.N_2075_tz_tz ;
    wire \POWERLED.N_600 ;
    wire \POWERLED.count_clk_en_0 ;
    wire \POWERLED.N_443 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_1 ;
    wire \POWERLED.N_443_cascade_ ;
    wire \POWERLED.count_clk_RNINSEUCZ0Z_7 ;
    wire \POWERLED.N_668 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_2 ;
    wire N_247;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_0 ;
    wire RSMRSTn_rep1;
    wire \POWERLED.N_506_cascade_ ;
    wire \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_10 ;
    wire \POWERLED.g0_i_0_1 ;
    wire \POWERLED.N_514_cascade_ ;
    wire \POWERLED.dutycycle_RNIHDMC5Z0Z_11 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.N_508 ;
    wire \POWERLED.N_512_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_11 ;
    wire \POWERLED.N_526_cascade_ ;
    wire \POWERLED.un1_clk_100khz_47_and_i_1 ;
    wire \POWERLED.dutycycle_en_11 ;
    wire \POWERLED.N_518_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.dutycycle_RNIE3861_0Z0Z_12 ;
    wire \POWERLED.N_520_cascade_ ;
    wire \POWERLED.dutycycle_RNIPK9V4Z0Z_12 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNIN405GZ0 ;
    wire \POWERLED.count_off_0_15 ;
    wire \POWERLED.count_off_RNI8AQHZ0Z_10 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_5 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_0_cascade_ ;
    wire \POWERLED.count_clk_RNIZ0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.count_clkZ0Z_1_cascade_ ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.count_off_1_14 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.count_off_0_7 ;
    wire \POWERLED.count_off_1_8 ;
    wire \POWERLED.count_off_0_8 ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.count_off_0_2 ;
    wire \POWERLED.count_off_1_5 ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_0_6 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_offZ0Z_6_cascade_ ;
    wire \POWERLED.un34_clk_100khz_9 ;
    wire \POWERLED.count_off_0_11 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_off_1_13 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_offZ0Z_13_cascade_ ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.un34_clk_100khz_10 ;
    wire \POWERLED.count_off_0_0 ;
    wire \POWERLED.count_off_1_0_cascade_ ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_offZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_RNIZ0Z_1 ;
    wire \POWERLED.N_123 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.count_off_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.un1_func_state25_6_0_0_a6_1_0_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_o_N_4 ;
    wire \POWERLED.un1_func_state25_6_0_0_0_2_1 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_5_cascade_ ;
    wire \POWERLED.N_421 ;
    wire \POWERLED.un1_func_state25_6_0_0_0_2_cascade_ ;
    wire \POWERLED.func_state_RNI31IBHZ0Z_0 ;
    wire \POWERLED.N_6_2 ;
    wire \POWERLED.func_state_RNI_0Z0Z_0 ;
    wire \POWERLED.func_state_RNIBVNSZ0Z_0 ;
    wire \POWERLED.count_off_RNI_0Z0Z_10 ;
    wire \POWERLED.func_state_RNI_3Z0Z_1 ;
    wire \POWERLED.func_state_RNIBVNSZ0Z_0_cascade_ ;
    wire \POWERLED.func_state_1_m0_1_1 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_7_2 ;
    wire rsmrst_pwrgd_signal;
    wire v5s_ok;
    wire vccst_cpu_ok;
    wire \VCCIN_PWRGD.un10_outputZ0Z_1_cascade_ ;
    wire v33s_ok;
    wire vccin_en;
    wire \POWERLED.N_253 ;
    wire \POWERLED.func_state_RNI_6Z0Z_1 ;
    wire \POWERLED.g1_1 ;
    wire \POWERLED.func_state_RNI_6Z0Z_1_cascade_ ;
    wire \POWERLED.N_2361_0_cascade_ ;
    wire N_6_0;
    wire \POWERLED.dutycycle_e_N_6L11_1 ;
    wire \POWERLED.dutycycle_RNI2MQDZ0Z_4_cascade_ ;
    wire \POWERLED.dutycycle_RNIOGRSZ0Z_4 ;
    wire \POWERLED.G_11_i_o10_1_0 ;
    wire \POWERLED.dutycycle ;
    wire N_9_0;
    wire RSMRSTn_rep2;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.N_488 ;
    wire \POWERLED.N_540_1 ;
    wire POWERLED_un1_dutycycle_172_m0_0;
    wire \POWERLED.N_435 ;
    wire \POWERLED.func_state_RNI_4Z0Z_1 ;
    wire \POWERLED.un1_dutycycle_172_m0_ns_1_0 ;
    wire \POWERLED.func_state_RNI_4Z0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI5DLRZ0Z_5 ;
    wire SUSWARN_N_rep1;
    wire \POWERLED.dutycycle_RNI7ABC3Z0Z_5_cascade_ ;
    wire COUNTER_un4_counter_7_THRU_CO;
    wire \POWERLED.g2_1_1 ;
    wire \POWERLED.g1_1cf0 ;
    wire \POWERLED.dutycycleZ1Z_5 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_5 ;
    wire \POWERLED.un1_clk_100khz_32_and_i_0cf0_cascade_ ;
    wire RSMRSTn_fast;
    wire \POWERLED.un1_clk_100khz_32_and_i_0 ;
    wire v5s_enn;
    wire \POWERLED.N_2291_i ;
    wire \POWERLED.N_676 ;
    wire \POWERLED.dutycycle_RNI6SKJ1Z0Z_3 ;
    wire \POWERLED.func_state_RNILP0FZ0Z_1_cascade_ ;
    wire \POWERLED.N_523 ;
    wire \POWERLED.dutycycleZ0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNIHDMC5Z0Z_3 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ;
    wire \POWERLED.dutycycleZ1Z_3 ;
    wire \POWERLED.N_430_iZ0 ;
    wire \POWERLED.N_5_0_cascade_ ;
    wire \POWERLED.N_12_2 ;
    wire \POWERLED.g0_7_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_4 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.i2_mux ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.N_2341_i_cascade_ ;
    wire \POWERLED.N_430 ;
    wire \POWERLED.N_529_cascade_ ;
    wire G_141;
    wire \POWERLED.dutycycle_en_12 ;
    wire \POWERLED.func_state_RNILP0FZ0Z_1 ;
    wire \POWERLED.func_state ;
    wire \POWERLED.N_527 ;
    wire \POWERLED.N_2341_i ;
    wire \POWERLED.un1_clk_100khz_48_and_i_1 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_8 ;
    wire \POWERLED.g0_i_0_0_0 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire vpp_en;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.G_7_i_o5_0 ;
    wire slp_s4n;
    wire gpio_fpga_soc_4;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycle_e_N_3L4_1 ;
    wire \POWERLED.func_state_RNI_8Z0Z_1 ;
    wire VCCST_EN_i_1;
    wire \POWERLED.N_203 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.N_505 ;
    wire count_clk_RNINSEUC_0_6;
    wire \POWERLED.N_412_i ;
    wire slp_s3n;
    wire \POWERLED.N_251 ;
    wire rsmrstn;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.N_524 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.func_state_RNIUQMRH_0_1 ;
    wire \POWERLED.count_clk_0_0 ;
    wire fpga_osc;
    wire \POWERLED.count_clk_en ;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__36183),
            .DIN(N__36182),
            .DOUT(N__36181),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__36183),
            .PADOUT(N__36182),
            .PADIN(N__36181),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__36174),
            .DIN(N__36173),
            .DOUT(N__36172),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__36174),
            .PADOUT(N__36173),
            .PADIN(N__36172),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19646),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__36165),
            .DIN(N__36164),
            .DOUT(N__36163),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__36165),
            .PADOUT(N__36164),
            .PADIN(N__36163),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19710),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__36156),
            .DIN(N__36155),
            .DOUT(N__36154),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__36156),
            .PADOUT(N__36155),
            .PADIN(N__36154),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14906),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__36147),
            .DIN(N__36146),
            .DOUT(N__36145),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__36147),
            .PADOUT(N__36146),
            .PADIN(N__36145),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__36138),
            .DIN(N__36137),
            .DOUT(N__36136),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__36138),
            .PADOUT(N__36137),
            .PADIN(N__36136),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__36129),
            .DIN(N__36128),
            .DOUT(N__36127),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__36129),
            .PADOUT(N__36128),
            .PADIN(N__36127),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__36120),
            .DIN(N__36119),
            .DOUT(N__36118),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__36120),
            .PADOUT(N__36119),
            .PADIN(N__36118),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__36111),
            .DIN(N__36110),
            .DOUT(N__36109),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__36111),
            .PADOUT(N__36110),
            .PADIN(N__36109),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30817),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__36102),
            .DIN(N__36101),
            .DOUT(N__36100),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__36102),
            .PADOUT(N__36101),
            .PADIN(N__36100),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__36093),
            .DIN(N__36092),
            .DOUT(N__36091),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__36093),
            .PADOUT(N__36092),
            .PADIN(N__36091),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__36084),
            .DIN(N__36083),
            .DOUT(N__36082),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__36084),
            .PADOUT(N__36083),
            .PADIN(N__36082),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14630),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__36075),
            .DIN(N__36074),
            .DOUT(N__36073),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__36075),
            .PADOUT(N__36074),
            .PADIN(N__36073),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__36066),
            .DIN(N__36065),
            .DOUT(N__36064),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__36066),
            .PADOUT(N__36065),
            .PADIN(N__36064),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_SLP_SUSn_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__36057),
            .DIN(N__36056),
            .DOUT(N__36055),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__36057),
            .PADOUT(N__36056),
            .PADIN(N__36055),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__36048),
            .DIN(N__36047),
            .DOUT(N__36046),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__36048),
            .PADOUT(N__36047),
            .PADIN(N__36046),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__36039),
            .DIN(N__36038),
            .DOUT(N__36037),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__36039),
            .PADOUT(N__36038),
            .PADIN(N__36037),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18557),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__36030),
            .DIN(N__36029),
            .DOUT(N__36028),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__36030),
            .PADOUT(N__36029),
            .PADIN(N__36028),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__36021),
            .DIN(N__36020),
            .DOUT(N__36019),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__36021),
            .PADOUT(N__36020),
            .PADIN(N__36019),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__36012),
            .DIN(N__36011),
            .DOUT(N__36010),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__36012),
            .PADOUT(N__36011),
            .PADIN(N__36010),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24697),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__36003),
            .DIN(N__36002),
            .DOUT(N__36001),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__36003),
            .PADOUT(N__36002),
            .PADIN(N__36001),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__35994),
            .DIN(N__35993),
            .DOUT(N__35992),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__35994),
            .PADOUT(N__35993),
            .PADIN(N__35992),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__35985),
            .DIN(N__35984),
            .DOUT(N__35983),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__35985),
            .PADOUT(N__35984),
            .PADIN(N__35983),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__35976),
            .DIN(N__35975),
            .DOUT(N__35974),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__35976),
            .PADOUT(N__35975),
            .PADIN(N__35974),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__35967),
            .DIN(N__35966),
            .DOUT(N__35965),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__35967),
            .PADOUT(N__35966),
            .PADIN(N__35965),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__35152),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__35958),
            .DIN(N__35957),
            .DOUT(N__35956),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__35958),
            .PADOUT(N__35957),
            .PADIN(N__35956),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__35949),
            .DIN(N__35948),
            .DOUT(N__35947),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__35949),
            .PADOUT(N__35948),
            .PADIN(N__35947),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19532),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__35940),
            .DIN(N__35939),
            .DOUT(N__35938),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__35940),
            .PADOUT(N__35939),
            .PADIN(N__35938),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25084),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__35931),
            .DIN(N__35930),
            .DOUT(N__35929),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__35931),
            .PADOUT(N__35930),
            .PADIN(N__35929),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__35922),
            .DIN(N__35921),
            .DOUT(N__35920),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__35922),
            .PADOUT(N__35921),
            .PADIN(N__35920),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__35913),
            .DIN(N__35912),
            .DOUT(N__35911),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__35913),
            .PADOUT(N__35912),
            .PADIN(N__35911),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__35904),
            .DIN(N__35903),
            .DOUT(N__35902),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__35904),
            .PADOUT(N__35903),
            .PADIN(N__35902),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__35895),
            .DIN(N__35894),
            .DOUT(N__35893),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__35895),
            .PADOUT(N__35894),
            .PADIN(N__35893),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__35886),
            .DIN(N__35885),
            .DOUT(N__35884),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__35886),
            .PADOUT(N__35885),
            .PADIN(N__35884),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14039),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__35877),
            .DIN(N__35876),
            .DOUT(N__35875),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__35877),
            .PADOUT(N__35876),
            .PADIN(N__35875),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__35868),
            .DIN(N__35867),
            .DOUT(N__35866),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__35868),
            .PADOUT(N__35867),
            .PADIN(N__35866),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32867),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__35859),
            .DIN(N__35858),
            .DOUT(N__35857),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__35859),
            .PADOUT(N__35858),
            .PADIN(N__35857),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__35850),
            .DIN(N__35849),
            .DOUT(N__35848),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__35850),
            .PADOUT(N__35849),
            .PADIN(N__35848),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__35841),
            .DIN(N__35840),
            .DOUT(N__35839),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__35841),
            .PADOUT(N__35840),
            .PADIN(N__35839),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__35832),
            .DIN(N__35831),
            .DOUT(N__35830),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__35832),
            .PADOUT(N__35831),
            .PADIN(N__35830),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__35823),
            .DIN(N__35822),
            .DOUT(N__35821),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__35823),
            .PADOUT(N__35822),
            .PADIN(N__35821),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19769),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__35814),
            .DIN(N__35813),
            .DOUT(N__35812),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__35814),
            .PADOUT(N__35813),
            .PADIN(N__35812),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__35805),
            .DIN(N__35804),
            .DOUT(N__35803),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__35805),
            .PADOUT(N__35804),
            .PADIN(N__35803),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30818),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__35796),
            .DIN(N__35795),
            .DOUT(N__35794),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__35796),
            .PADOUT(N__35795),
            .PADIN(N__35794),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    defparam ipInertedIOPad_DSW_PWROK_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__35787),
            .DIN(N__35786),
            .DOUT(N__35785),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__35787),
            .PADOUT(N__35786),
            .PADIN(N__35785),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23135),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__35778),
            .DIN(N__35777),
            .DOUT(N__35776),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__35778),
            .PADOUT(N__35777),
            .PADIN(N__35776),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19724),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__35769),
            .DIN(N__35768),
            .DOUT(N__35767),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__35769),
            .PADOUT(N__35768),
            .PADIN(N__35767),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__35760),
            .DIN(N__35759),
            .DOUT(N__35758),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__35760),
            .PADOUT(N__35759),
            .PADIN(N__35758),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__35751),
            .DIN(N__35750),
            .DOUT(N__35749),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__35751),
            .PADOUT(N__35750),
            .PADIN(N__35749),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__35742),
            .DIN(N__35741),
            .DOUT(N__35740),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__35742),
            .PADOUT(N__35741),
            .PADIN(N__35740),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__35733),
            .DIN(N__35732),
            .DOUT(N__35731),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__35733),
            .PADOUT(N__35732),
            .PADIN(N__35731),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29732),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__35724),
            .DIN(N__35723),
            .DOUT(N__35722),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__35724),
            .PADOUT(N__35723),
            .PADIN(N__35722),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__35715),
            .DIN(N__35714),
            .DOUT(N__35713),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__35715),
            .PADOUT(N__35714),
            .PADIN(N__35713),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__35706),
            .DIN(N__35705),
            .DOUT(N__35704),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__35706),
            .PADOUT(N__35705),
            .PADIN(N__35704),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__35697),
            .DIN(N__35696),
            .DOUT(N__35695),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__35697),
            .PADOUT(N__35696),
            .PADIN(N__35695),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__35688),
            .DIN(N__35687),
            .DOUT(N__35686),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__35688),
            .PADOUT(N__35687),
            .PADIN(N__35686),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__35679),
            .DIN(N__35678),
            .DOUT(N__35677),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__35679),
            .PADOUT(N__35678),
            .PADIN(N__35677),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__35670),
            .DIN(N__35669),
            .DOUT(N__35668),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__35670),
            .PADOUT(N__35669),
            .PADIN(N__35668),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25088),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__35661),
            .DIN(N__35660),
            .DOUT(N__35659),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__35661),
            .PADOUT(N__35660),
            .PADIN(N__35659),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__8387 (
            .O(N__35642),
            .I(N__35638));
    CascadeMux I__8386 (
            .O(N__35641),
            .I(N__35630));
    LocalMux I__8385 (
            .O(N__35638),
            .I(N__35626));
    InMux I__8384 (
            .O(N__35637),
            .I(N__35614));
    InMux I__8383 (
            .O(N__35636),
            .I(N__35614));
    InMux I__8382 (
            .O(N__35635),
            .I(N__35614));
    InMux I__8381 (
            .O(N__35634),
            .I(N__35614));
    InMux I__8380 (
            .O(N__35633),
            .I(N__35614));
    InMux I__8379 (
            .O(N__35630),
            .I(N__35611));
    InMux I__8378 (
            .O(N__35629),
            .I(N__35608));
    Span4Mux_v I__8377 (
            .O(N__35626),
            .I(N__35605));
    InMux I__8376 (
            .O(N__35625),
            .I(N__35602));
    LocalMux I__8375 (
            .O(N__35614),
            .I(N__35597));
    LocalMux I__8374 (
            .O(N__35611),
            .I(N__35597));
    LocalMux I__8373 (
            .O(N__35608),
            .I(N__35594));
    Span4Mux_v I__8372 (
            .O(N__35605),
            .I(N__35591));
    LocalMux I__8371 (
            .O(N__35602),
            .I(N__35586));
    Sp12to4 I__8370 (
            .O(N__35597),
            .I(N__35586));
    Span4Mux_s2_h I__8369 (
            .O(N__35594),
            .I(N__35583));
    Odrv4 I__8368 (
            .O(N__35591),
            .I(count_clk_RNINSEUC_0_6));
    Odrv12 I__8367 (
            .O(N__35586),
            .I(count_clk_RNINSEUC_0_6));
    Odrv4 I__8366 (
            .O(N__35583),
            .I(count_clk_RNINSEUC_0_6));
    InMux I__8365 (
            .O(N__35576),
            .I(N__35572));
    CascadeMux I__8364 (
            .O(N__35575),
            .I(N__35569));
    LocalMux I__8363 (
            .O(N__35572),
            .I(N__35565));
    InMux I__8362 (
            .O(N__35569),
            .I(N__35562));
    CascadeMux I__8361 (
            .O(N__35568),
            .I(N__35558));
    Span4Mux_v I__8360 (
            .O(N__35565),
            .I(N__35552));
    LocalMux I__8359 (
            .O(N__35562),
            .I(N__35552));
    InMux I__8358 (
            .O(N__35561),
            .I(N__35548));
    InMux I__8357 (
            .O(N__35558),
            .I(N__35545));
    InMux I__8356 (
            .O(N__35557),
            .I(N__35542));
    Span4Mux_h I__8355 (
            .O(N__35552),
            .I(N__35537));
    CascadeMux I__8354 (
            .O(N__35551),
            .I(N__35534));
    LocalMux I__8353 (
            .O(N__35548),
            .I(N__35526));
    LocalMux I__8352 (
            .O(N__35545),
            .I(N__35526));
    LocalMux I__8351 (
            .O(N__35542),
            .I(N__35526));
    InMux I__8350 (
            .O(N__35541),
            .I(N__35523));
    InMux I__8349 (
            .O(N__35540),
            .I(N__35520));
    Span4Mux_v I__8348 (
            .O(N__35537),
            .I(N__35517));
    InMux I__8347 (
            .O(N__35534),
            .I(N__35512));
    InMux I__8346 (
            .O(N__35533),
            .I(N__35512));
    Span4Mux_v I__8345 (
            .O(N__35526),
            .I(N__35507));
    LocalMux I__8344 (
            .O(N__35523),
            .I(N__35507));
    LocalMux I__8343 (
            .O(N__35520),
            .I(N__35504));
    Odrv4 I__8342 (
            .O(N__35517),
            .I(\POWERLED.N_412_i ));
    LocalMux I__8341 (
            .O(N__35512),
            .I(\POWERLED.N_412_i ));
    Odrv4 I__8340 (
            .O(N__35507),
            .I(\POWERLED.N_412_i ));
    Odrv12 I__8339 (
            .O(N__35504),
            .I(\POWERLED.N_412_i ));
    CascadeMux I__8338 (
            .O(N__35495),
            .I(N__35492));
    InMux I__8337 (
            .O(N__35492),
            .I(N__35485));
    InMux I__8336 (
            .O(N__35491),
            .I(N__35485));
    CascadeMux I__8335 (
            .O(N__35490),
            .I(N__35482));
    LocalMux I__8334 (
            .O(N__35485),
            .I(N__35477));
    InMux I__8333 (
            .O(N__35482),
            .I(N__35467));
    InMux I__8332 (
            .O(N__35481),
            .I(N__35462));
    InMux I__8331 (
            .O(N__35480),
            .I(N__35462));
    Span4Mux_v I__8330 (
            .O(N__35477),
            .I(N__35459));
    CascadeMux I__8329 (
            .O(N__35476),
            .I(N__35454));
    CascadeMux I__8328 (
            .O(N__35475),
            .I(N__35451));
    InMux I__8327 (
            .O(N__35474),
            .I(N__35439));
    InMux I__8326 (
            .O(N__35473),
            .I(N__35430));
    InMux I__8325 (
            .O(N__35472),
            .I(N__35430));
    InMux I__8324 (
            .O(N__35471),
            .I(N__35430));
    InMux I__8323 (
            .O(N__35470),
            .I(N__35430));
    LocalMux I__8322 (
            .O(N__35467),
            .I(N__35425));
    LocalMux I__8321 (
            .O(N__35462),
            .I(N__35425));
    Span4Mux_v I__8320 (
            .O(N__35459),
            .I(N__35422));
    InMux I__8319 (
            .O(N__35458),
            .I(N__35419));
    InMux I__8318 (
            .O(N__35457),
            .I(N__35416));
    InMux I__8317 (
            .O(N__35454),
            .I(N__35413));
    InMux I__8316 (
            .O(N__35451),
            .I(N__35410));
    InMux I__8315 (
            .O(N__35450),
            .I(N__35404));
    InMux I__8314 (
            .O(N__35449),
            .I(N__35404));
    InMux I__8313 (
            .O(N__35448),
            .I(N__35394));
    InMux I__8312 (
            .O(N__35447),
            .I(N__35394));
    InMux I__8311 (
            .O(N__35446),
            .I(N__35394));
    InMux I__8310 (
            .O(N__35445),
            .I(N__35394));
    InMux I__8309 (
            .O(N__35444),
            .I(N__35391));
    InMux I__8308 (
            .O(N__35443),
            .I(N__35385));
    InMux I__8307 (
            .O(N__35442),
            .I(N__35385));
    LocalMux I__8306 (
            .O(N__35439),
            .I(N__35380));
    LocalMux I__8305 (
            .O(N__35430),
            .I(N__35380));
    Span4Mux_v I__8304 (
            .O(N__35425),
            .I(N__35374));
    Span4Mux_h I__8303 (
            .O(N__35422),
            .I(N__35369));
    LocalMux I__8302 (
            .O(N__35419),
            .I(N__35369));
    LocalMux I__8301 (
            .O(N__35416),
            .I(N__35366));
    LocalMux I__8300 (
            .O(N__35413),
            .I(N__35361));
    LocalMux I__8299 (
            .O(N__35410),
            .I(N__35361));
    InMux I__8298 (
            .O(N__35409),
            .I(N__35358));
    LocalMux I__8297 (
            .O(N__35404),
            .I(N__35355));
    InMux I__8296 (
            .O(N__35403),
            .I(N__35352));
    LocalMux I__8295 (
            .O(N__35394),
            .I(N__35346));
    LocalMux I__8294 (
            .O(N__35391),
            .I(N__35346));
    CascadeMux I__8293 (
            .O(N__35390),
            .I(N__35341));
    LocalMux I__8292 (
            .O(N__35385),
            .I(N__35337));
    Span4Mux_h I__8291 (
            .O(N__35380),
            .I(N__35334));
    InMux I__8290 (
            .O(N__35379),
            .I(N__35331));
    InMux I__8289 (
            .O(N__35378),
            .I(N__35326));
    InMux I__8288 (
            .O(N__35377),
            .I(N__35326));
    IoSpan4Mux I__8287 (
            .O(N__35374),
            .I(N__35321));
    Span4Mux_v I__8286 (
            .O(N__35369),
            .I(N__35318));
    Span4Mux_v I__8285 (
            .O(N__35366),
            .I(N__35311));
    Span4Mux_v I__8284 (
            .O(N__35361),
            .I(N__35311));
    LocalMux I__8283 (
            .O(N__35358),
            .I(N__35311));
    Span4Mux_h I__8282 (
            .O(N__35355),
            .I(N__35308));
    LocalMux I__8281 (
            .O(N__35352),
            .I(N__35305));
    InMux I__8280 (
            .O(N__35351),
            .I(N__35302));
    Span4Mux_s1_h I__8279 (
            .O(N__35346),
            .I(N__35299));
    InMux I__8278 (
            .O(N__35345),
            .I(N__35294));
    InMux I__8277 (
            .O(N__35344),
            .I(N__35294));
    InMux I__8276 (
            .O(N__35341),
            .I(N__35289));
    InMux I__8275 (
            .O(N__35340),
            .I(N__35289));
    Span4Mux_v I__8274 (
            .O(N__35337),
            .I(N__35286));
    Span4Mux_v I__8273 (
            .O(N__35334),
            .I(N__35279));
    LocalMux I__8272 (
            .O(N__35331),
            .I(N__35279));
    LocalMux I__8271 (
            .O(N__35326),
            .I(N__35279));
    InMux I__8270 (
            .O(N__35325),
            .I(N__35276));
    InMux I__8269 (
            .O(N__35324),
            .I(N__35273));
    IoSpan4Mux I__8268 (
            .O(N__35321),
            .I(N__35269));
    Span4Mux_s2_v I__8267 (
            .O(N__35318),
            .I(N__35264));
    Span4Mux_v I__8266 (
            .O(N__35311),
            .I(N__35264));
    Span4Mux_v I__8265 (
            .O(N__35308),
            .I(N__35259));
    Span4Mux_s1_h I__8264 (
            .O(N__35305),
            .I(N__35259));
    LocalMux I__8263 (
            .O(N__35302),
            .I(N__35256));
    Span4Mux_v I__8262 (
            .O(N__35299),
            .I(N__35249));
    LocalMux I__8261 (
            .O(N__35294),
            .I(N__35249));
    LocalMux I__8260 (
            .O(N__35289),
            .I(N__35249));
    Span4Mux_h I__8259 (
            .O(N__35286),
            .I(N__35240));
    Span4Mux_v I__8258 (
            .O(N__35279),
            .I(N__35240));
    LocalMux I__8257 (
            .O(N__35276),
            .I(N__35240));
    LocalMux I__8256 (
            .O(N__35273),
            .I(N__35240));
    InMux I__8255 (
            .O(N__35272),
            .I(N__35237));
    IoSpan4Mux I__8254 (
            .O(N__35269),
            .I(N__35232));
    IoSpan4Mux I__8253 (
            .O(N__35264),
            .I(N__35232));
    Span4Mux_v I__8252 (
            .O(N__35259),
            .I(N__35225));
    Span4Mux_s1_h I__8251 (
            .O(N__35256),
            .I(N__35225));
    Span4Mux_v I__8250 (
            .O(N__35249),
            .I(N__35225));
    Span4Mux_v I__8249 (
            .O(N__35240),
            .I(N__35220));
    LocalMux I__8248 (
            .O(N__35237),
            .I(N__35220));
    Odrv4 I__8247 (
            .O(N__35232),
            .I(slp_s3n));
    Odrv4 I__8246 (
            .O(N__35225),
            .I(slp_s3n));
    Odrv4 I__8245 (
            .O(N__35220),
            .I(slp_s3n));
    InMux I__8244 (
            .O(N__35213),
            .I(N__35210));
    LocalMux I__8243 (
            .O(N__35210),
            .I(N__35203));
    InMux I__8242 (
            .O(N__35209),
            .I(N__35200));
    InMux I__8241 (
            .O(N__35208),
            .I(N__35195));
    InMux I__8240 (
            .O(N__35207),
            .I(N__35195));
    CascadeMux I__8239 (
            .O(N__35206),
            .I(N__35191));
    Span4Mux_v I__8238 (
            .O(N__35203),
            .I(N__35188));
    LocalMux I__8237 (
            .O(N__35200),
            .I(N__35183));
    LocalMux I__8236 (
            .O(N__35195),
            .I(N__35183));
    InMux I__8235 (
            .O(N__35194),
            .I(N__35180));
    InMux I__8234 (
            .O(N__35191),
            .I(N__35177));
    Span4Mux_v I__8233 (
            .O(N__35188),
            .I(N__35172));
    Sp12to4 I__8232 (
            .O(N__35183),
            .I(N__35165));
    LocalMux I__8231 (
            .O(N__35180),
            .I(N__35165));
    LocalMux I__8230 (
            .O(N__35177),
            .I(N__35165));
    InMux I__8229 (
            .O(N__35176),
            .I(N__35160));
    InMux I__8228 (
            .O(N__35175),
            .I(N__35160));
    Odrv4 I__8227 (
            .O(N__35172),
            .I(\POWERLED.N_251 ));
    Odrv12 I__8226 (
            .O(N__35165),
            .I(\POWERLED.N_251 ));
    LocalMux I__8225 (
            .O(N__35160),
            .I(\POWERLED.N_251 ));
    CascadeMux I__8224 (
            .O(N__35153),
            .I(N__35149));
    IoInMux I__8223 (
            .O(N__35152),
            .I(N__35145));
    InMux I__8222 (
            .O(N__35149),
            .I(N__35139));
    CascadeMux I__8221 (
            .O(N__35148),
            .I(N__35136));
    LocalMux I__8220 (
            .O(N__35145),
            .I(N__35132));
    CascadeMux I__8219 (
            .O(N__35144),
            .I(N__35128));
    InMux I__8218 (
            .O(N__35143),
            .I(N__35123));
    InMux I__8217 (
            .O(N__35142),
            .I(N__35120));
    LocalMux I__8216 (
            .O(N__35139),
            .I(N__35115));
    InMux I__8215 (
            .O(N__35136),
            .I(N__35112));
    CascadeMux I__8214 (
            .O(N__35135),
            .I(N__35107));
    Span4Mux_s3_v I__8213 (
            .O(N__35132),
            .I(N__35104));
    InMux I__8212 (
            .O(N__35131),
            .I(N__35101));
    InMux I__8211 (
            .O(N__35128),
            .I(N__35098));
    InMux I__8210 (
            .O(N__35127),
            .I(N__35094));
    InMux I__8209 (
            .O(N__35126),
            .I(N__35091));
    LocalMux I__8208 (
            .O(N__35123),
            .I(N__35086));
    LocalMux I__8207 (
            .O(N__35120),
            .I(N__35086));
    InMux I__8206 (
            .O(N__35119),
            .I(N__35082));
    InMux I__8205 (
            .O(N__35118),
            .I(N__35079));
    Span4Mux_s1_h I__8204 (
            .O(N__35115),
            .I(N__35074));
    LocalMux I__8203 (
            .O(N__35112),
            .I(N__35074));
    InMux I__8202 (
            .O(N__35111),
            .I(N__35071));
    InMux I__8201 (
            .O(N__35110),
            .I(N__35068));
    InMux I__8200 (
            .O(N__35107),
            .I(N__35065));
    Span4Mux_v I__8199 (
            .O(N__35104),
            .I(N__35060));
    LocalMux I__8198 (
            .O(N__35101),
            .I(N__35060));
    LocalMux I__8197 (
            .O(N__35098),
            .I(N__35057));
    InMux I__8196 (
            .O(N__35097),
            .I(N__35054));
    LocalMux I__8195 (
            .O(N__35094),
            .I(N__35051));
    LocalMux I__8194 (
            .O(N__35091),
            .I(N__35044));
    Span4Mux_s3_h I__8193 (
            .O(N__35086),
            .I(N__35044));
    InMux I__8192 (
            .O(N__35085),
            .I(N__35041));
    LocalMux I__8191 (
            .O(N__35082),
            .I(N__35036));
    LocalMux I__8190 (
            .O(N__35079),
            .I(N__35036));
    Span4Mux_v I__8189 (
            .O(N__35074),
            .I(N__35031));
    LocalMux I__8188 (
            .O(N__35071),
            .I(N__35031));
    LocalMux I__8187 (
            .O(N__35068),
            .I(N__35028));
    LocalMux I__8186 (
            .O(N__35065),
            .I(N__35025));
    Span4Mux_h I__8185 (
            .O(N__35060),
            .I(N__35018));
    Span4Mux_h I__8184 (
            .O(N__35057),
            .I(N__35018));
    LocalMux I__8183 (
            .O(N__35054),
            .I(N__35018));
    Span4Mux_s3_h I__8182 (
            .O(N__35051),
            .I(N__35015));
    InMux I__8181 (
            .O(N__35050),
            .I(N__35012));
    InMux I__8180 (
            .O(N__35049),
            .I(N__35009));
    Span4Mux_v I__8179 (
            .O(N__35044),
            .I(N__35004));
    LocalMux I__8178 (
            .O(N__35041),
            .I(N__35004));
    Span4Mux_v I__8177 (
            .O(N__35036),
            .I(N__34995));
    Span4Mux_v I__8176 (
            .O(N__35031),
            .I(N__34995));
    Span4Mux_s1_h I__8175 (
            .O(N__35028),
            .I(N__34995));
    Span4Mux_s1_h I__8174 (
            .O(N__35025),
            .I(N__34995));
    Span4Mux_v I__8173 (
            .O(N__35018),
            .I(N__34992));
    Span4Mux_v I__8172 (
            .O(N__35015),
            .I(N__34987));
    LocalMux I__8171 (
            .O(N__35012),
            .I(N__34987));
    LocalMux I__8170 (
            .O(N__35009),
            .I(N__34982));
    Span4Mux_v I__8169 (
            .O(N__35004),
            .I(N__34982));
    Span4Mux_v I__8168 (
            .O(N__34995),
            .I(N__34977));
    Span4Mux_v I__8167 (
            .O(N__34992),
            .I(N__34977));
    Odrv4 I__8166 (
            .O(N__34987),
            .I(rsmrstn));
    Odrv4 I__8165 (
            .O(N__34982),
            .I(rsmrstn));
    Odrv4 I__8164 (
            .O(N__34977),
            .I(rsmrstn));
    CascadeMux I__8163 (
            .O(N__34970),
            .I(N__34964));
    InMux I__8162 (
            .O(N__34969),
            .I(N__34961));
    CascadeMux I__8161 (
            .O(N__34968),
            .I(N__34956));
    CascadeMux I__8160 (
            .O(N__34967),
            .I(N__34953));
    InMux I__8159 (
            .O(N__34964),
            .I(N__34950));
    LocalMux I__8158 (
            .O(N__34961),
            .I(N__34947));
    InMux I__8157 (
            .O(N__34960),
            .I(N__34944));
    InMux I__8156 (
            .O(N__34959),
            .I(N__34941));
    InMux I__8155 (
            .O(N__34956),
            .I(N__34938));
    InMux I__8154 (
            .O(N__34953),
            .I(N__34931));
    LocalMux I__8153 (
            .O(N__34950),
            .I(N__34928));
    Span4Mux_v I__8152 (
            .O(N__34947),
            .I(N__34925));
    LocalMux I__8151 (
            .O(N__34944),
            .I(N__34918));
    LocalMux I__8150 (
            .O(N__34941),
            .I(N__34918));
    LocalMux I__8149 (
            .O(N__34938),
            .I(N__34918));
    InMux I__8148 (
            .O(N__34937),
            .I(N__34915));
    InMux I__8147 (
            .O(N__34936),
            .I(N__34912));
    InMux I__8146 (
            .O(N__34935),
            .I(N__34909));
    InMux I__8145 (
            .O(N__34934),
            .I(N__34906));
    LocalMux I__8144 (
            .O(N__34931),
            .I(N__34901));
    Span4Mux_s3_h I__8143 (
            .O(N__34928),
            .I(N__34901));
    Odrv4 I__8142 (
            .O(N__34925),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv12 I__8141 (
            .O(N__34918),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__8140 (
            .O(N__34915),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__8139 (
            .O(N__34912),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__8138 (
            .O(N__34909),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__8137 (
            .O(N__34906),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__8136 (
            .O(N__34901),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    InMux I__8135 (
            .O(N__34886),
            .I(N__34883));
    LocalMux I__8134 (
            .O(N__34883),
            .I(\POWERLED.N_524 ));
    CascadeMux I__8133 (
            .O(N__34880),
            .I(N__34876));
    CascadeMux I__8132 (
            .O(N__34879),
            .I(N__34873));
    InMux I__8131 (
            .O(N__34876),
            .I(N__34869));
    InMux I__8130 (
            .O(N__34873),
            .I(N__34866));
    InMux I__8129 (
            .O(N__34872),
            .I(N__34861));
    LocalMux I__8128 (
            .O(N__34869),
            .I(N__34858));
    LocalMux I__8127 (
            .O(N__34866),
            .I(N__34855));
    InMux I__8126 (
            .O(N__34865),
            .I(N__34850));
    InMux I__8125 (
            .O(N__34864),
            .I(N__34850));
    LocalMux I__8124 (
            .O(N__34861),
            .I(N__34847));
    Span4Mux_h I__8123 (
            .O(N__34858),
            .I(N__34844));
    Odrv4 I__8122 (
            .O(N__34855),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__8121 (
            .O(N__34850),
            .I(\POWERLED.count_clkZ0Z_0 ));
    Odrv4 I__8120 (
            .O(N__34847),
            .I(\POWERLED.count_clkZ0Z_0 ));
    Odrv4 I__8119 (
            .O(N__34844),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__8118 (
            .O(N__34835),
            .I(N__34821));
    InMux I__8117 (
            .O(N__34834),
            .I(N__34821));
    InMux I__8116 (
            .O(N__34833),
            .I(N__34821));
    InMux I__8115 (
            .O(N__34832),
            .I(N__34821));
    InMux I__8114 (
            .O(N__34831),
            .I(N__34816));
    InMux I__8113 (
            .O(N__34830),
            .I(N__34816));
    LocalMux I__8112 (
            .O(N__34821),
            .I(N__34803));
    LocalMux I__8111 (
            .O(N__34816),
            .I(N__34803));
    InMux I__8110 (
            .O(N__34815),
            .I(N__34794));
    InMux I__8109 (
            .O(N__34814),
            .I(N__34794));
    InMux I__8108 (
            .O(N__34813),
            .I(N__34794));
    InMux I__8107 (
            .O(N__34812),
            .I(N__34794));
    InMux I__8106 (
            .O(N__34811),
            .I(N__34787));
    InMux I__8105 (
            .O(N__34810),
            .I(N__34787));
    InMux I__8104 (
            .O(N__34809),
            .I(N__34787));
    InMux I__8103 (
            .O(N__34808),
            .I(N__34779));
    Span4Mux_s1_v I__8102 (
            .O(N__34803),
            .I(N__34772));
    LocalMux I__8101 (
            .O(N__34794),
            .I(N__34772));
    LocalMux I__8100 (
            .O(N__34787),
            .I(N__34772));
    InMux I__8099 (
            .O(N__34786),
            .I(N__34761));
    InMux I__8098 (
            .O(N__34785),
            .I(N__34761));
    InMux I__8097 (
            .O(N__34784),
            .I(N__34761));
    InMux I__8096 (
            .O(N__34783),
            .I(N__34761));
    InMux I__8095 (
            .O(N__34782),
            .I(N__34761));
    LocalMux I__8094 (
            .O(N__34779),
            .I(\POWERLED.func_state_RNIUQMRH_0_1 ));
    Odrv4 I__8093 (
            .O(N__34772),
            .I(\POWERLED.func_state_RNIUQMRH_0_1 ));
    LocalMux I__8092 (
            .O(N__34761),
            .I(\POWERLED.func_state_RNIUQMRH_0_1 ));
    InMux I__8091 (
            .O(N__34754),
            .I(N__34751));
    LocalMux I__8090 (
            .O(N__34751),
            .I(N__34748));
    Span4Mux_s2_v I__8089 (
            .O(N__34748),
            .I(N__34745));
    Odrv4 I__8088 (
            .O(N__34745),
            .I(\POWERLED.count_clk_0_0 ));
    ClkMux I__8087 (
            .O(N__34742),
            .I(N__34734));
    ClkMux I__8086 (
            .O(N__34741),
            .I(N__34731));
    ClkMux I__8085 (
            .O(N__34740),
            .I(N__34728));
    ClkMux I__8084 (
            .O(N__34739),
            .I(N__34721));
    ClkMux I__8083 (
            .O(N__34738),
            .I(N__34712));
    ClkMux I__8082 (
            .O(N__34737),
            .I(N__34709));
    LocalMux I__8081 (
            .O(N__34734),
            .I(N__34705));
    LocalMux I__8080 (
            .O(N__34731),
            .I(N__34702));
    LocalMux I__8079 (
            .O(N__34728),
            .I(N__34696));
    ClkMux I__8078 (
            .O(N__34727),
            .I(N__34693));
    ClkMux I__8077 (
            .O(N__34726),
            .I(N__34690));
    ClkMux I__8076 (
            .O(N__34725),
            .I(N__34687));
    ClkMux I__8075 (
            .O(N__34724),
            .I(N__34682));
    LocalMux I__8074 (
            .O(N__34721),
            .I(N__34673));
    ClkMux I__8073 (
            .O(N__34720),
            .I(N__34670));
    ClkMux I__8072 (
            .O(N__34719),
            .I(N__34667));
    ClkMux I__8071 (
            .O(N__34718),
            .I(N__34664));
    ClkMux I__8070 (
            .O(N__34717),
            .I(N__34661));
    ClkMux I__8069 (
            .O(N__34716),
            .I(N__34657));
    ClkMux I__8068 (
            .O(N__34715),
            .I(N__34652));
    LocalMux I__8067 (
            .O(N__34712),
            .I(N__34645));
    LocalMux I__8066 (
            .O(N__34709),
            .I(N__34645));
    ClkMux I__8065 (
            .O(N__34708),
            .I(N__34642));
    Span4Mux_v I__8064 (
            .O(N__34705),
            .I(N__34639));
    Span4Mux_s3_h I__8063 (
            .O(N__34702),
            .I(N__34636));
    ClkMux I__8062 (
            .O(N__34701),
            .I(N__34633));
    ClkMux I__8061 (
            .O(N__34700),
            .I(N__34630));
    ClkMux I__8060 (
            .O(N__34699),
            .I(N__34627));
    Span4Mux_v I__8059 (
            .O(N__34696),
            .I(N__34622));
    LocalMux I__8058 (
            .O(N__34693),
            .I(N__34622));
    LocalMux I__8057 (
            .O(N__34690),
            .I(N__34616));
    LocalMux I__8056 (
            .O(N__34687),
            .I(N__34616));
    ClkMux I__8055 (
            .O(N__34686),
            .I(N__34613));
    ClkMux I__8054 (
            .O(N__34685),
            .I(N__34610));
    LocalMux I__8053 (
            .O(N__34682),
            .I(N__34607));
    ClkMux I__8052 (
            .O(N__34681),
            .I(N__34604));
    ClkMux I__8051 (
            .O(N__34680),
            .I(N__34601));
    ClkMux I__8050 (
            .O(N__34679),
            .I(N__34597));
    ClkMux I__8049 (
            .O(N__34678),
            .I(N__34593));
    ClkMux I__8048 (
            .O(N__34677),
            .I(N__34589));
    ClkMux I__8047 (
            .O(N__34676),
            .I(N__34586));
    Span4Mux_s2_v I__8046 (
            .O(N__34673),
            .I(N__34577));
    LocalMux I__8045 (
            .O(N__34670),
            .I(N__34577));
    LocalMux I__8044 (
            .O(N__34667),
            .I(N__34574));
    LocalMux I__8043 (
            .O(N__34664),
            .I(N__34570));
    LocalMux I__8042 (
            .O(N__34661),
            .I(N__34567));
    ClkMux I__8041 (
            .O(N__34660),
            .I(N__34564));
    LocalMux I__8040 (
            .O(N__34657),
            .I(N__34561));
    ClkMux I__8039 (
            .O(N__34656),
            .I(N__34558));
    ClkMux I__8038 (
            .O(N__34655),
            .I(N__34554));
    LocalMux I__8037 (
            .O(N__34652),
            .I(N__34547));
    ClkMux I__8036 (
            .O(N__34651),
            .I(N__34544));
    ClkMux I__8035 (
            .O(N__34650),
            .I(N__34541));
    Span4Mux_s3_v I__8034 (
            .O(N__34645),
            .I(N__34534));
    LocalMux I__8033 (
            .O(N__34642),
            .I(N__34534));
    Span4Mux_h I__8032 (
            .O(N__34639),
            .I(N__34525));
    Span4Mux_h I__8031 (
            .O(N__34636),
            .I(N__34525));
    LocalMux I__8030 (
            .O(N__34633),
            .I(N__34525));
    LocalMux I__8029 (
            .O(N__34630),
            .I(N__34522));
    LocalMux I__8028 (
            .O(N__34627),
            .I(N__34517));
    Span4Mux_v I__8027 (
            .O(N__34622),
            .I(N__34517));
    ClkMux I__8026 (
            .O(N__34621),
            .I(N__34514));
    Span4Mux_h I__8025 (
            .O(N__34616),
            .I(N__34506));
    LocalMux I__8024 (
            .O(N__34613),
            .I(N__34506));
    LocalMux I__8023 (
            .O(N__34610),
            .I(N__34506));
    Span4Mux_s1_v I__8022 (
            .O(N__34607),
            .I(N__34499));
    LocalMux I__8021 (
            .O(N__34604),
            .I(N__34499));
    LocalMux I__8020 (
            .O(N__34601),
            .I(N__34499));
    ClkMux I__8019 (
            .O(N__34600),
            .I(N__34496));
    LocalMux I__8018 (
            .O(N__34597),
            .I(N__34492));
    ClkMux I__8017 (
            .O(N__34596),
            .I(N__34486));
    LocalMux I__8016 (
            .O(N__34593),
            .I(N__34483));
    ClkMux I__8015 (
            .O(N__34592),
            .I(N__34480));
    LocalMux I__8014 (
            .O(N__34589),
            .I(N__34475));
    LocalMux I__8013 (
            .O(N__34586),
            .I(N__34475));
    ClkMux I__8012 (
            .O(N__34585),
            .I(N__34472));
    ClkMux I__8011 (
            .O(N__34584),
            .I(N__34469));
    ClkMux I__8010 (
            .O(N__34583),
            .I(N__34466));
    ClkMux I__8009 (
            .O(N__34582),
            .I(N__34460));
    Span4Mux_v I__8008 (
            .O(N__34577),
            .I(N__34455));
    Span4Mux_s1_h I__8007 (
            .O(N__34574),
            .I(N__34455));
    ClkMux I__8006 (
            .O(N__34573),
            .I(N__34452));
    Span4Mux_s2_v I__8005 (
            .O(N__34570),
            .I(N__34444));
    Span4Mux_s2_h I__8004 (
            .O(N__34567),
            .I(N__34444));
    LocalMux I__8003 (
            .O(N__34564),
            .I(N__34444));
    Span4Mux_s1_h I__8002 (
            .O(N__34561),
            .I(N__34439));
    LocalMux I__8001 (
            .O(N__34558),
            .I(N__34439));
    ClkMux I__8000 (
            .O(N__34557),
            .I(N__34436));
    LocalMux I__7999 (
            .O(N__34554),
            .I(N__34433));
    ClkMux I__7998 (
            .O(N__34553),
            .I(N__34430));
    ClkMux I__7997 (
            .O(N__34552),
            .I(N__34427));
    ClkMux I__7996 (
            .O(N__34551),
            .I(N__34420));
    ClkMux I__7995 (
            .O(N__34550),
            .I(N__34417));
    Span4Mux_v I__7994 (
            .O(N__34547),
            .I(N__34409));
    LocalMux I__7993 (
            .O(N__34544),
            .I(N__34409));
    LocalMux I__7992 (
            .O(N__34541),
            .I(N__34409));
    ClkMux I__7991 (
            .O(N__34540),
            .I(N__34406));
    ClkMux I__7990 (
            .O(N__34539),
            .I(N__34400));
    Span4Mux_v I__7989 (
            .O(N__34534),
            .I(N__34395));
    ClkMux I__7988 (
            .O(N__34533),
            .I(N__34392));
    ClkMux I__7987 (
            .O(N__34532),
            .I(N__34389));
    Span4Mux_v I__7986 (
            .O(N__34525),
            .I(N__34380));
    Span4Mux_h I__7985 (
            .O(N__34522),
            .I(N__34380));
    Span4Mux_h I__7984 (
            .O(N__34517),
            .I(N__34380));
    LocalMux I__7983 (
            .O(N__34514),
            .I(N__34380));
    ClkMux I__7982 (
            .O(N__34513),
            .I(N__34377));
    Span4Mux_v I__7981 (
            .O(N__34506),
            .I(N__34370));
    Span4Mux_v I__7980 (
            .O(N__34499),
            .I(N__34370));
    LocalMux I__7979 (
            .O(N__34496),
            .I(N__34370));
    ClkMux I__7978 (
            .O(N__34495),
            .I(N__34367));
    Span4Mux_v I__7977 (
            .O(N__34492),
            .I(N__34364));
    ClkMux I__7976 (
            .O(N__34491),
            .I(N__34361));
    ClkMux I__7975 (
            .O(N__34490),
            .I(N__34358));
    ClkMux I__7974 (
            .O(N__34489),
            .I(N__34355));
    LocalMux I__7973 (
            .O(N__34486),
            .I(N__34347));
    Span4Mux_h I__7972 (
            .O(N__34483),
            .I(N__34347));
    LocalMux I__7971 (
            .O(N__34480),
            .I(N__34347));
    Span4Mux_v I__7970 (
            .O(N__34475),
            .I(N__34340));
    LocalMux I__7969 (
            .O(N__34472),
            .I(N__34340));
    LocalMux I__7968 (
            .O(N__34469),
            .I(N__34340));
    LocalMux I__7967 (
            .O(N__34466),
            .I(N__34337));
    ClkMux I__7966 (
            .O(N__34465),
            .I(N__34334));
    ClkMux I__7965 (
            .O(N__34464),
            .I(N__34330));
    ClkMux I__7964 (
            .O(N__34463),
            .I(N__34327));
    LocalMux I__7963 (
            .O(N__34460),
            .I(N__34323));
    Span4Mux_v I__7962 (
            .O(N__34455),
            .I(N__34318));
    LocalMux I__7961 (
            .O(N__34452),
            .I(N__34318));
    ClkMux I__7960 (
            .O(N__34451),
            .I(N__34315));
    Span4Mux_v I__7959 (
            .O(N__34444),
            .I(N__34312));
    Span4Mux_h I__7958 (
            .O(N__34439),
            .I(N__34307));
    LocalMux I__7957 (
            .O(N__34436),
            .I(N__34307));
    Span4Mux_s2_v I__7956 (
            .O(N__34433),
            .I(N__34300));
    LocalMux I__7955 (
            .O(N__34430),
            .I(N__34300));
    LocalMux I__7954 (
            .O(N__34427),
            .I(N__34300));
    ClkMux I__7953 (
            .O(N__34426),
            .I(N__34297));
    ClkMux I__7952 (
            .O(N__34425),
            .I(N__34294));
    ClkMux I__7951 (
            .O(N__34424),
            .I(N__34290));
    ClkMux I__7950 (
            .O(N__34423),
            .I(N__34287));
    LocalMux I__7949 (
            .O(N__34420),
            .I(N__34283));
    LocalMux I__7948 (
            .O(N__34417),
            .I(N__34280));
    ClkMux I__7947 (
            .O(N__34416),
            .I(N__34277));
    Span4Mux_v I__7946 (
            .O(N__34409),
            .I(N__34272));
    LocalMux I__7945 (
            .O(N__34406),
            .I(N__34272));
    ClkMux I__7944 (
            .O(N__34405),
            .I(N__34269));
    ClkMux I__7943 (
            .O(N__34404),
            .I(N__34266));
    ClkMux I__7942 (
            .O(N__34403),
            .I(N__34261));
    LocalMux I__7941 (
            .O(N__34400),
            .I(N__34258));
    ClkMux I__7940 (
            .O(N__34399),
            .I(N__34255));
    ClkMux I__7939 (
            .O(N__34398),
            .I(N__34251));
    Span4Mux_v I__7938 (
            .O(N__34395),
            .I(N__34246));
    LocalMux I__7937 (
            .O(N__34392),
            .I(N__34246));
    LocalMux I__7936 (
            .O(N__34389),
            .I(N__34242));
    Span4Mux_v I__7935 (
            .O(N__34380),
            .I(N__34239));
    LocalMux I__7934 (
            .O(N__34377),
            .I(N__34236));
    Span4Mux_v I__7933 (
            .O(N__34370),
            .I(N__34227));
    LocalMux I__7932 (
            .O(N__34367),
            .I(N__34227));
    Span4Mux_s2_v I__7931 (
            .O(N__34364),
            .I(N__34227));
    LocalMux I__7930 (
            .O(N__34361),
            .I(N__34227));
    LocalMux I__7929 (
            .O(N__34358),
            .I(N__34222));
    LocalMux I__7928 (
            .O(N__34355),
            .I(N__34222));
    ClkMux I__7927 (
            .O(N__34354),
            .I(N__34219));
    Span4Mux_v I__7926 (
            .O(N__34347),
            .I(N__34210));
    Span4Mux_v I__7925 (
            .O(N__34340),
            .I(N__34210));
    Span4Mux_s3_h I__7924 (
            .O(N__34337),
            .I(N__34210));
    LocalMux I__7923 (
            .O(N__34334),
            .I(N__34210));
    ClkMux I__7922 (
            .O(N__34333),
            .I(N__34207));
    LocalMux I__7921 (
            .O(N__34330),
            .I(N__34202));
    LocalMux I__7920 (
            .O(N__34327),
            .I(N__34202));
    ClkMux I__7919 (
            .O(N__34326),
            .I(N__34199));
    Span4Mux_h I__7918 (
            .O(N__34323),
            .I(N__34195));
    Span4Mux_v I__7917 (
            .O(N__34318),
            .I(N__34190));
    LocalMux I__7916 (
            .O(N__34315),
            .I(N__34190));
    Span4Mux_h I__7915 (
            .O(N__34312),
            .I(N__34179));
    Span4Mux_v I__7914 (
            .O(N__34307),
            .I(N__34179));
    Span4Mux_v I__7913 (
            .O(N__34300),
            .I(N__34179));
    LocalMux I__7912 (
            .O(N__34297),
            .I(N__34179));
    LocalMux I__7911 (
            .O(N__34294),
            .I(N__34179));
    ClkMux I__7910 (
            .O(N__34293),
            .I(N__34176));
    LocalMux I__7909 (
            .O(N__34290),
            .I(N__34173));
    LocalMux I__7908 (
            .O(N__34287),
            .I(N__34170));
    ClkMux I__7907 (
            .O(N__34286),
            .I(N__34167));
    Span4Mux_v I__7906 (
            .O(N__34283),
            .I(N__34160));
    Span4Mux_h I__7905 (
            .O(N__34280),
            .I(N__34160));
    LocalMux I__7904 (
            .O(N__34277),
            .I(N__34160));
    Span4Mux_v I__7903 (
            .O(N__34272),
            .I(N__34155));
    LocalMux I__7902 (
            .O(N__34269),
            .I(N__34155));
    LocalMux I__7901 (
            .O(N__34266),
            .I(N__34152));
    ClkMux I__7900 (
            .O(N__34265),
            .I(N__34149));
    ClkMux I__7899 (
            .O(N__34264),
            .I(N__34146));
    LocalMux I__7898 (
            .O(N__34261),
            .I(N__34143));
    Span4Mux_h I__7897 (
            .O(N__34258),
            .I(N__34138));
    LocalMux I__7896 (
            .O(N__34255),
            .I(N__34138));
    ClkMux I__7895 (
            .O(N__34254),
            .I(N__34135));
    LocalMux I__7894 (
            .O(N__34251),
            .I(N__34130));
    Sp12to4 I__7893 (
            .O(N__34246),
            .I(N__34130));
    ClkMux I__7892 (
            .O(N__34245),
            .I(N__34127));
    IoSpan4Mux I__7891 (
            .O(N__34242),
            .I(N__34124));
    Span4Mux_h I__7890 (
            .O(N__34239),
            .I(N__34121));
    Span4Mux_h I__7889 (
            .O(N__34236),
            .I(N__34112));
    Span4Mux_v I__7888 (
            .O(N__34227),
            .I(N__34112));
    Span4Mux_v I__7887 (
            .O(N__34222),
            .I(N__34112));
    LocalMux I__7886 (
            .O(N__34219),
            .I(N__34112));
    Span4Mux_v I__7885 (
            .O(N__34210),
            .I(N__34107));
    LocalMux I__7884 (
            .O(N__34207),
            .I(N__34107));
    Span4Mux_s2_v I__7883 (
            .O(N__34202),
            .I(N__34104));
    LocalMux I__7882 (
            .O(N__34199),
            .I(N__34101));
    ClkMux I__7881 (
            .O(N__34198),
            .I(N__34098));
    Span4Mux_v I__7880 (
            .O(N__34195),
            .I(N__34089));
    Span4Mux_h I__7879 (
            .O(N__34190),
            .I(N__34089));
    Span4Mux_v I__7878 (
            .O(N__34179),
            .I(N__34089));
    LocalMux I__7877 (
            .O(N__34176),
            .I(N__34089));
    Span4Mux_s1_h I__7876 (
            .O(N__34173),
            .I(N__34082));
    Span4Mux_s1_h I__7875 (
            .O(N__34170),
            .I(N__34082));
    LocalMux I__7874 (
            .O(N__34167),
            .I(N__34082));
    Span4Mux_v I__7873 (
            .O(N__34160),
            .I(N__34071));
    Span4Mux_s2_h I__7872 (
            .O(N__34155),
            .I(N__34071));
    Span4Mux_s2_h I__7871 (
            .O(N__34152),
            .I(N__34071));
    LocalMux I__7870 (
            .O(N__34149),
            .I(N__34071));
    LocalMux I__7869 (
            .O(N__34146),
            .I(N__34071));
    Span4Mux_s2_h I__7868 (
            .O(N__34143),
            .I(N__34064));
    Span4Mux_h I__7867 (
            .O(N__34138),
            .I(N__34064));
    LocalMux I__7866 (
            .O(N__34135),
            .I(N__34064));
    Span12Mux_s5_h I__7865 (
            .O(N__34130),
            .I(N__34056));
    LocalMux I__7864 (
            .O(N__34127),
            .I(N__34056));
    IoSpan4Mux I__7863 (
            .O(N__34124),
            .I(N__34047));
    IoSpan4Mux I__7862 (
            .O(N__34121),
            .I(N__34047));
    IoSpan4Mux I__7861 (
            .O(N__34112),
            .I(N__34047));
    IoSpan4Mux I__7860 (
            .O(N__34107),
            .I(N__34047));
    Span4Mux_h I__7859 (
            .O(N__34104),
            .I(N__34040));
    Span4Mux_h I__7858 (
            .O(N__34101),
            .I(N__34040));
    LocalMux I__7857 (
            .O(N__34098),
            .I(N__34040));
    Span4Mux_v I__7856 (
            .O(N__34089),
            .I(N__34033));
    Span4Mux_h I__7855 (
            .O(N__34082),
            .I(N__34033));
    Span4Mux_h I__7854 (
            .O(N__34071),
            .I(N__34033));
    Span4Mux_h I__7853 (
            .O(N__34064),
            .I(N__34030));
    ClkMux I__7852 (
            .O(N__34063),
            .I(N__34027));
    ClkMux I__7851 (
            .O(N__34062),
            .I(N__34024));
    ClkMux I__7850 (
            .O(N__34061),
            .I(N__34021));
    Odrv12 I__7849 (
            .O(N__34056),
            .I(fpga_osc));
    Odrv4 I__7848 (
            .O(N__34047),
            .I(fpga_osc));
    Odrv4 I__7847 (
            .O(N__34040),
            .I(fpga_osc));
    Odrv4 I__7846 (
            .O(N__34033),
            .I(fpga_osc));
    Odrv4 I__7845 (
            .O(N__34030),
            .I(fpga_osc));
    LocalMux I__7844 (
            .O(N__34027),
            .I(fpga_osc));
    LocalMux I__7843 (
            .O(N__34024),
            .I(fpga_osc));
    LocalMux I__7842 (
            .O(N__34021),
            .I(fpga_osc));
    CEMux I__7841 (
            .O(N__34004),
            .I(N__33999));
    CEMux I__7840 (
            .O(N__34003),
            .I(N__33993));
    CEMux I__7839 (
            .O(N__34002),
            .I(N__33989));
    LocalMux I__7838 (
            .O(N__33999),
            .I(N__33979));
    CascadeMux I__7837 (
            .O(N__33998),
            .I(N__33974));
    CascadeMux I__7836 (
            .O(N__33997),
            .I(N__33971));
    CEMux I__7835 (
            .O(N__33996),
            .I(N__33967));
    LocalMux I__7834 (
            .O(N__33993),
            .I(N__33964));
    CEMux I__7833 (
            .O(N__33992),
            .I(N__33961));
    LocalMux I__7832 (
            .O(N__33989),
            .I(N__33958));
    InMux I__7831 (
            .O(N__33988),
            .I(N__33948));
    InMux I__7830 (
            .O(N__33987),
            .I(N__33948));
    InMux I__7829 (
            .O(N__33986),
            .I(N__33948));
    CascadeMux I__7828 (
            .O(N__33985),
            .I(N__33945));
    InMux I__7827 (
            .O(N__33984),
            .I(N__33937));
    InMux I__7826 (
            .O(N__33983),
            .I(N__33937));
    InMux I__7825 (
            .O(N__33982),
            .I(N__33937));
    Span4Mux_s2_v I__7824 (
            .O(N__33979),
            .I(N__33930));
    InMux I__7823 (
            .O(N__33978),
            .I(N__33927));
    InMux I__7822 (
            .O(N__33977),
            .I(N__33918));
    InMux I__7821 (
            .O(N__33974),
            .I(N__33918));
    InMux I__7820 (
            .O(N__33971),
            .I(N__33918));
    InMux I__7819 (
            .O(N__33970),
            .I(N__33918));
    LocalMux I__7818 (
            .O(N__33967),
            .I(N__33910));
    Span4Mux_s1_h I__7817 (
            .O(N__33964),
            .I(N__33910));
    LocalMux I__7816 (
            .O(N__33961),
            .I(N__33907));
    Span4Mux_v I__7815 (
            .O(N__33958),
            .I(N__33904));
    InMux I__7814 (
            .O(N__33957),
            .I(N__33899));
    InMux I__7813 (
            .O(N__33956),
            .I(N__33899));
    InMux I__7812 (
            .O(N__33955),
            .I(N__33896));
    LocalMux I__7811 (
            .O(N__33948),
            .I(N__33893));
    InMux I__7810 (
            .O(N__33945),
            .I(N__33888));
    InMux I__7809 (
            .O(N__33944),
            .I(N__33888));
    LocalMux I__7808 (
            .O(N__33937),
            .I(N__33885));
    CEMux I__7807 (
            .O(N__33936),
            .I(N__33882));
    CEMux I__7806 (
            .O(N__33935),
            .I(N__33879));
    CEMux I__7805 (
            .O(N__33934),
            .I(N__33876));
    CEMux I__7804 (
            .O(N__33933),
            .I(N__33873));
    Span4Mux_s3_h I__7803 (
            .O(N__33930),
            .I(N__33870));
    LocalMux I__7802 (
            .O(N__33927),
            .I(N__33865));
    LocalMux I__7801 (
            .O(N__33918),
            .I(N__33865));
    InMux I__7800 (
            .O(N__33917),
            .I(N__33858));
    InMux I__7799 (
            .O(N__33916),
            .I(N__33858));
    InMux I__7798 (
            .O(N__33915),
            .I(N__33858));
    Span4Mux_s2_v I__7797 (
            .O(N__33910),
            .I(N__33841));
    Span4Mux_s2_v I__7796 (
            .O(N__33907),
            .I(N__33841));
    Span4Mux_v I__7795 (
            .O(N__33904),
            .I(N__33841));
    LocalMux I__7794 (
            .O(N__33899),
            .I(N__33841));
    LocalMux I__7793 (
            .O(N__33896),
            .I(N__33841));
    Span4Mux_h I__7792 (
            .O(N__33893),
            .I(N__33841));
    LocalMux I__7791 (
            .O(N__33888),
            .I(N__33841));
    Span4Mux_s2_v I__7790 (
            .O(N__33885),
            .I(N__33841));
    LocalMux I__7789 (
            .O(N__33882),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7788 (
            .O(N__33879),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7787 (
            .O(N__33876),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7786 (
            .O(N__33873),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__7785 (
            .O(N__33870),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__7784 (
            .O(N__33865),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7783 (
            .O(N__33858),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__7782 (
            .O(N__33841),
            .I(\POWERLED.count_clk_en ));
    CascadeMux I__7781 (
            .O(N__33824),
            .I(\POWERLED.N_2341_i_cascade_ ));
    InMux I__7780 (
            .O(N__33821),
            .I(N__33812));
    InMux I__7779 (
            .O(N__33820),
            .I(N__33812));
    InMux I__7778 (
            .O(N__33819),
            .I(N__33808));
    InMux I__7777 (
            .O(N__33818),
            .I(N__33805));
    InMux I__7776 (
            .O(N__33817),
            .I(N__33799));
    LocalMux I__7775 (
            .O(N__33812),
            .I(N__33796));
    InMux I__7774 (
            .O(N__33811),
            .I(N__33790));
    LocalMux I__7773 (
            .O(N__33808),
            .I(N__33786));
    LocalMux I__7772 (
            .O(N__33805),
            .I(N__33783));
    InMux I__7771 (
            .O(N__33804),
            .I(N__33780));
    InMux I__7770 (
            .O(N__33803),
            .I(N__33777));
    InMux I__7769 (
            .O(N__33802),
            .I(N__33773));
    LocalMux I__7768 (
            .O(N__33799),
            .I(N__33768));
    Span4Mux_h I__7767 (
            .O(N__33796),
            .I(N__33768));
    InMux I__7766 (
            .O(N__33795),
            .I(N__33765));
    InMux I__7765 (
            .O(N__33794),
            .I(N__33762));
    InMux I__7764 (
            .O(N__33793),
            .I(N__33759));
    LocalMux I__7763 (
            .O(N__33790),
            .I(N__33756));
    InMux I__7762 (
            .O(N__33789),
            .I(N__33753));
    Span4Mux_s3_h I__7761 (
            .O(N__33786),
            .I(N__33748));
    Span4Mux_v I__7760 (
            .O(N__33783),
            .I(N__33748));
    LocalMux I__7759 (
            .O(N__33780),
            .I(N__33743));
    LocalMux I__7758 (
            .O(N__33777),
            .I(N__33743));
    InMux I__7757 (
            .O(N__33776),
            .I(N__33740));
    LocalMux I__7756 (
            .O(N__33773),
            .I(N__33728));
    Span4Mux_v I__7755 (
            .O(N__33768),
            .I(N__33728));
    LocalMux I__7754 (
            .O(N__33765),
            .I(N__33728));
    LocalMux I__7753 (
            .O(N__33762),
            .I(N__33725));
    LocalMux I__7752 (
            .O(N__33759),
            .I(N__33718));
    Span4Mux_v I__7751 (
            .O(N__33756),
            .I(N__33718));
    LocalMux I__7750 (
            .O(N__33753),
            .I(N__33718));
    Span4Mux_v I__7749 (
            .O(N__33748),
            .I(N__33713));
    Span4Mux_s3_h I__7748 (
            .O(N__33743),
            .I(N__33713));
    LocalMux I__7747 (
            .O(N__33740),
            .I(N__33710));
    InMux I__7746 (
            .O(N__33739),
            .I(N__33707));
    InMux I__7745 (
            .O(N__33738),
            .I(N__33704));
    InMux I__7744 (
            .O(N__33737),
            .I(N__33697));
    InMux I__7743 (
            .O(N__33736),
            .I(N__33697));
    InMux I__7742 (
            .O(N__33735),
            .I(N__33697));
    Span4Mux_v I__7741 (
            .O(N__33728),
            .I(N__33690));
    Span4Mux_s0_h I__7740 (
            .O(N__33725),
            .I(N__33690));
    Span4Mux_v I__7739 (
            .O(N__33718),
            .I(N__33690));
    Odrv4 I__7738 (
            .O(N__33713),
            .I(\POWERLED.N_430 ));
    Odrv4 I__7737 (
            .O(N__33710),
            .I(\POWERLED.N_430 ));
    LocalMux I__7736 (
            .O(N__33707),
            .I(\POWERLED.N_430 ));
    LocalMux I__7735 (
            .O(N__33704),
            .I(\POWERLED.N_430 ));
    LocalMux I__7734 (
            .O(N__33697),
            .I(\POWERLED.N_430 ));
    Odrv4 I__7733 (
            .O(N__33690),
            .I(\POWERLED.N_430 ));
    CascadeMux I__7732 (
            .O(N__33677),
            .I(\POWERLED.N_529_cascade_ ));
    CascadeMux I__7731 (
            .O(N__33674),
            .I(N__33663));
    InMux I__7730 (
            .O(N__33673),
            .I(N__33652));
    InMux I__7729 (
            .O(N__33672),
            .I(N__33652));
    CascadeMux I__7728 (
            .O(N__33671),
            .I(N__33648));
    CascadeMux I__7727 (
            .O(N__33670),
            .I(N__33645));
    CascadeMux I__7726 (
            .O(N__33669),
            .I(N__33639));
    InMux I__7725 (
            .O(N__33668),
            .I(N__33636));
    InMux I__7724 (
            .O(N__33667),
            .I(N__33631));
    InMux I__7723 (
            .O(N__33666),
            .I(N__33628));
    InMux I__7722 (
            .O(N__33663),
            .I(N__33625));
    InMux I__7721 (
            .O(N__33662),
            .I(N__33622));
    InMux I__7720 (
            .O(N__33661),
            .I(N__33618));
    InMux I__7719 (
            .O(N__33660),
            .I(N__33615));
    InMux I__7718 (
            .O(N__33659),
            .I(N__33612));
    InMux I__7717 (
            .O(N__33658),
            .I(N__33607));
    InMux I__7716 (
            .O(N__33657),
            .I(N__33607));
    LocalMux I__7715 (
            .O(N__33652),
            .I(N__33604));
    InMux I__7714 (
            .O(N__33651),
            .I(N__33595));
    InMux I__7713 (
            .O(N__33648),
            .I(N__33595));
    InMux I__7712 (
            .O(N__33645),
            .I(N__33590));
    InMux I__7711 (
            .O(N__33644),
            .I(N__33590));
    CascadeMux I__7710 (
            .O(N__33643),
            .I(N__33586));
    CascadeMux I__7709 (
            .O(N__33642),
            .I(N__33583));
    InMux I__7708 (
            .O(N__33639),
            .I(N__33579));
    LocalMux I__7707 (
            .O(N__33636),
            .I(N__33576));
    InMux I__7706 (
            .O(N__33635),
            .I(N__33571));
    InMux I__7705 (
            .O(N__33634),
            .I(N__33571));
    LocalMux I__7704 (
            .O(N__33631),
            .I(N__33566));
    LocalMux I__7703 (
            .O(N__33628),
            .I(N__33566));
    LocalMux I__7702 (
            .O(N__33625),
            .I(N__33561));
    LocalMux I__7701 (
            .O(N__33622),
            .I(N__33561));
    IoInMux I__7700 (
            .O(N__33621),
            .I(N__33558));
    LocalMux I__7699 (
            .O(N__33618),
            .I(N__33555));
    LocalMux I__7698 (
            .O(N__33615),
            .I(N__33548));
    LocalMux I__7697 (
            .O(N__33612),
            .I(N__33548));
    LocalMux I__7696 (
            .O(N__33607),
            .I(N__33548));
    Span4Mux_h I__7695 (
            .O(N__33604),
            .I(N__33545));
    InMux I__7694 (
            .O(N__33603),
            .I(N__33540));
    InMux I__7693 (
            .O(N__33602),
            .I(N__33533));
    InMux I__7692 (
            .O(N__33601),
            .I(N__33533));
    InMux I__7691 (
            .O(N__33600),
            .I(N__33533));
    LocalMux I__7690 (
            .O(N__33595),
            .I(N__33528));
    LocalMux I__7689 (
            .O(N__33590),
            .I(N__33528));
    InMux I__7688 (
            .O(N__33589),
            .I(N__33523));
    InMux I__7687 (
            .O(N__33586),
            .I(N__33523));
    InMux I__7686 (
            .O(N__33583),
            .I(N__33518));
    InMux I__7685 (
            .O(N__33582),
            .I(N__33518));
    LocalMux I__7684 (
            .O(N__33579),
            .I(N__33515));
    Span4Mux_v I__7683 (
            .O(N__33576),
            .I(N__33510));
    LocalMux I__7682 (
            .O(N__33571),
            .I(N__33510));
    Span4Mux_v I__7681 (
            .O(N__33566),
            .I(N__33505));
    Span4Mux_s0_h I__7680 (
            .O(N__33561),
            .I(N__33505));
    LocalMux I__7679 (
            .O(N__33558),
            .I(N__33502));
    Span4Mux_v I__7678 (
            .O(N__33555),
            .I(N__33497));
    Span4Mux_v I__7677 (
            .O(N__33548),
            .I(N__33497));
    Span4Mux_v I__7676 (
            .O(N__33545),
            .I(N__33494));
    InMux I__7675 (
            .O(N__33544),
            .I(N__33489));
    InMux I__7674 (
            .O(N__33543),
            .I(N__33489));
    LocalMux I__7673 (
            .O(N__33540),
            .I(N__33484));
    LocalMux I__7672 (
            .O(N__33533),
            .I(N__33484));
    Span12Mux_s5_h I__7671 (
            .O(N__33528),
            .I(N__33479));
    LocalMux I__7670 (
            .O(N__33523),
            .I(N__33479));
    LocalMux I__7669 (
            .O(N__33518),
            .I(N__33470));
    Span4Mux_v I__7668 (
            .O(N__33515),
            .I(N__33470));
    Span4Mux_h I__7667 (
            .O(N__33510),
            .I(N__33470));
    Span4Mux_h I__7666 (
            .O(N__33505),
            .I(N__33470));
    Odrv12 I__7665 (
            .O(N__33502),
            .I(G_141));
    Odrv4 I__7664 (
            .O(N__33497),
            .I(G_141));
    Odrv4 I__7663 (
            .O(N__33494),
            .I(G_141));
    LocalMux I__7662 (
            .O(N__33489),
            .I(G_141));
    Odrv4 I__7661 (
            .O(N__33484),
            .I(G_141));
    Odrv12 I__7660 (
            .O(N__33479),
            .I(G_141));
    Odrv4 I__7659 (
            .O(N__33470),
            .I(G_141));
    CascadeMux I__7658 (
            .O(N__33455),
            .I(N__33452));
    InMux I__7657 (
            .O(N__33452),
            .I(N__33446));
    InMux I__7656 (
            .O(N__33451),
            .I(N__33446));
    LocalMux I__7655 (
            .O(N__33446),
            .I(N__33443));
    Span4Mux_h I__7654 (
            .O(N__33443),
            .I(N__33440));
    Odrv4 I__7653 (
            .O(N__33440),
            .I(\POWERLED.dutycycle_en_12 ));
    InMux I__7652 (
            .O(N__33437),
            .I(N__33429));
    InMux I__7651 (
            .O(N__33436),
            .I(N__33426));
    InMux I__7650 (
            .O(N__33435),
            .I(N__33423));
    InMux I__7649 (
            .O(N__33434),
            .I(N__33418));
    InMux I__7648 (
            .O(N__33433),
            .I(N__33418));
    InMux I__7647 (
            .O(N__33432),
            .I(N__33415));
    LocalMux I__7646 (
            .O(N__33429),
            .I(N__33412));
    LocalMux I__7645 (
            .O(N__33426),
            .I(N__33409));
    LocalMux I__7644 (
            .O(N__33423),
            .I(N__33404));
    LocalMux I__7643 (
            .O(N__33418),
            .I(N__33404));
    LocalMux I__7642 (
            .O(N__33415),
            .I(N__33397));
    Span4Mux_h I__7641 (
            .O(N__33412),
            .I(N__33397));
    Span4Mux_v I__7640 (
            .O(N__33409),
            .I(N__33394));
    Span4Mux_v I__7639 (
            .O(N__33404),
            .I(N__33391));
    InMux I__7638 (
            .O(N__33403),
            .I(N__33386));
    InMux I__7637 (
            .O(N__33402),
            .I(N__33386));
    Odrv4 I__7636 (
            .O(N__33397),
            .I(\POWERLED.func_state_RNILP0FZ0Z_1 ));
    Odrv4 I__7635 (
            .O(N__33394),
            .I(\POWERLED.func_state_RNILP0FZ0Z_1 ));
    Odrv4 I__7634 (
            .O(N__33391),
            .I(\POWERLED.func_state_RNILP0FZ0Z_1 ));
    LocalMux I__7633 (
            .O(N__33386),
            .I(\POWERLED.func_state_RNILP0FZ0Z_1 ));
    CascadeMux I__7632 (
            .O(N__33377),
            .I(N__33373));
    InMux I__7631 (
            .O(N__33376),
            .I(N__33355));
    InMux I__7630 (
            .O(N__33373),
            .I(N__33350));
    InMux I__7629 (
            .O(N__33372),
            .I(N__33350));
    CascadeMux I__7628 (
            .O(N__33371),
            .I(N__33346));
    InMux I__7627 (
            .O(N__33370),
            .I(N__33342));
    InMux I__7626 (
            .O(N__33369),
            .I(N__33339));
    InMux I__7625 (
            .O(N__33368),
            .I(N__33330));
    InMux I__7624 (
            .O(N__33367),
            .I(N__33330));
    InMux I__7623 (
            .O(N__33366),
            .I(N__33330));
    InMux I__7622 (
            .O(N__33365),
            .I(N__33330));
    InMux I__7621 (
            .O(N__33364),
            .I(N__33327));
    InMux I__7620 (
            .O(N__33363),
            .I(N__33318));
    InMux I__7619 (
            .O(N__33362),
            .I(N__33318));
    InMux I__7618 (
            .O(N__33361),
            .I(N__33318));
    InMux I__7617 (
            .O(N__33360),
            .I(N__33318));
    InMux I__7616 (
            .O(N__33359),
            .I(N__33313));
    InMux I__7615 (
            .O(N__33358),
            .I(N__33313));
    LocalMux I__7614 (
            .O(N__33355),
            .I(N__33308));
    LocalMux I__7613 (
            .O(N__33350),
            .I(N__33308));
    InMux I__7612 (
            .O(N__33349),
            .I(N__33303));
    InMux I__7611 (
            .O(N__33346),
            .I(N__33303));
    InMux I__7610 (
            .O(N__33345),
            .I(N__33284));
    LocalMux I__7609 (
            .O(N__33342),
            .I(N__33281));
    LocalMux I__7608 (
            .O(N__33339),
            .I(N__33273));
    LocalMux I__7607 (
            .O(N__33330),
            .I(N__33273));
    LocalMux I__7606 (
            .O(N__33327),
            .I(N__33273));
    LocalMux I__7605 (
            .O(N__33318),
            .I(N__33268));
    LocalMux I__7604 (
            .O(N__33313),
            .I(N__33268));
    Span4Mux_s2_h I__7603 (
            .O(N__33308),
            .I(N__33263));
    LocalMux I__7602 (
            .O(N__33303),
            .I(N__33263));
    InMux I__7601 (
            .O(N__33302),
            .I(N__33258));
    InMux I__7600 (
            .O(N__33301),
            .I(N__33258));
    InMux I__7599 (
            .O(N__33300),
            .I(N__33253));
    InMux I__7598 (
            .O(N__33299),
            .I(N__33253));
    InMux I__7597 (
            .O(N__33298),
            .I(N__33248));
    InMux I__7596 (
            .O(N__33297),
            .I(N__33248));
    InMux I__7595 (
            .O(N__33296),
            .I(N__33243));
    InMux I__7594 (
            .O(N__33295),
            .I(N__33243));
    InMux I__7593 (
            .O(N__33294),
            .I(N__33236));
    InMux I__7592 (
            .O(N__33293),
            .I(N__33236));
    InMux I__7591 (
            .O(N__33292),
            .I(N__33236));
    InMux I__7590 (
            .O(N__33291),
            .I(N__33231));
    InMux I__7589 (
            .O(N__33290),
            .I(N__33231));
    InMux I__7588 (
            .O(N__33289),
            .I(N__33228));
    InMux I__7587 (
            .O(N__33288),
            .I(N__33223));
    InMux I__7586 (
            .O(N__33287),
            .I(N__33223));
    LocalMux I__7585 (
            .O(N__33284),
            .I(N__33218));
    Span4Mux_v I__7584 (
            .O(N__33281),
            .I(N__33218));
    InMux I__7583 (
            .O(N__33280),
            .I(N__33215));
    Span4Mux_v I__7582 (
            .O(N__33273),
            .I(N__33208));
    Span4Mux_h I__7581 (
            .O(N__33268),
            .I(N__33208));
    Span4Mux_v I__7580 (
            .O(N__33263),
            .I(N__33208));
    LocalMux I__7579 (
            .O(N__33258),
            .I(N__33193));
    LocalMux I__7578 (
            .O(N__33253),
            .I(N__33193));
    LocalMux I__7577 (
            .O(N__33248),
            .I(N__33193));
    LocalMux I__7576 (
            .O(N__33243),
            .I(N__33193));
    LocalMux I__7575 (
            .O(N__33236),
            .I(N__33193));
    LocalMux I__7574 (
            .O(N__33231),
            .I(N__33193));
    LocalMux I__7573 (
            .O(N__33228),
            .I(N__33193));
    LocalMux I__7572 (
            .O(N__33223),
            .I(\POWERLED.func_state ));
    Odrv4 I__7571 (
            .O(N__33218),
            .I(\POWERLED.func_state ));
    LocalMux I__7570 (
            .O(N__33215),
            .I(\POWERLED.func_state ));
    Odrv4 I__7569 (
            .O(N__33208),
            .I(\POWERLED.func_state ));
    Odrv12 I__7568 (
            .O(N__33193),
            .I(\POWERLED.func_state ));
    CascadeMux I__7567 (
            .O(N__33182),
            .I(N__33179));
    InMux I__7566 (
            .O(N__33179),
            .I(N__33176));
    LocalMux I__7565 (
            .O(N__33176),
            .I(\POWERLED.N_527 ));
    InMux I__7564 (
            .O(N__33173),
            .I(N__33170));
    LocalMux I__7563 (
            .O(N__33170),
            .I(N__33166));
    InMux I__7562 (
            .O(N__33169),
            .I(N__33163));
    Span4Mux_v I__7561 (
            .O(N__33166),
            .I(N__33160));
    LocalMux I__7560 (
            .O(N__33163),
            .I(N__33155));
    Span4Mux_h I__7559 (
            .O(N__33160),
            .I(N__33155));
    Odrv4 I__7558 (
            .O(N__33155),
            .I(\POWERLED.N_2341_i ));
    InMux I__7557 (
            .O(N__33152),
            .I(N__33149));
    LocalMux I__7556 (
            .O(N__33149),
            .I(\POWERLED.un1_clk_100khz_48_and_i_1 ));
    CascadeMux I__7555 (
            .O(N__33146),
            .I(N__33138));
    CascadeMux I__7554 (
            .O(N__33145),
            .I(N__33129));
    InMux I__7553 (
            .O(N__33144),
            .I(N__33125));
    InMux I__7552 (
            .O(N__33143),
            .I(N__33119));
    InMux I__7551 (
            .O(N__33142),
            .I(N__33116));
    InMux I__7550 (
            .O(N__33141),
            .I(N__33112));
    InMux I__7549 (
            .O(N__33138),
            .I(N__33109));
    InMux I__7548 (
            .O(N__33137),
            .I(N__33101));
    InMux I__7547 (
            .O(N__33136),
            .I(N__33101));
    InMux I__7546 (
            .O(N__33135),
            .I(N__33098));
    InMux I__7545 (
            .O(N__33134),
            .I(N__33095));
    InMux I__7544 (
            .O(N__33133),
            .I(N__33090));
    InMux I__7543 (
            .O(N__33132),
            .I(N__33090));
    InMux I__7542 (
            .O(N__33129),
            .I(N__33082));
    InMux I__7541 (
            .O(N__33128),
            .I(N__33082));
    LocalMux I__7540 (
            .O(N__33125),
            .I(N__33079));
    InMux I__7539 (
            .O(N__33124),
            .I(N__33076));
    InMux I__7538 (
            .O(N__33123),
            .I(N__33073));
    InMux I__7537 (
            .O(N__33122),
            .I(N__33070));
    LocalMux I__7536 (
            .O(N__33119),
            .I(N__33065));
    LocalMux I__7535 (
            .O(N__33116),
            .I(N__33065));
    InMux I__7534 (
            .O(N__33115),
            .I(N__33062));
    LocalMux I__7533 (
            .O(N__33112),
            .I(N__33057));
    LocalMux I__7532 (
            .O(N__33109),
            .I(N__33057));
    InMux I__7531 (
            .O(N__33108),
            .I(N__33053));
    InMux I__7530 (
            .O(N__33107),
            .I(N__33048));
    InMux I__7529 (
            .O(N__33106),
            .I(N__33045));
    LocalMux I__7528 (
            .O(N__33101),
            .I(N__33042));
    LocalMux I__7527 (
            .O(N__33098),
            .I(N__33035));
    LocalMux I__7526 (
            .O(N__33095),
            .I(N__33035));
    LocalMux I__7525 (
            .O(N__33090),
            .I(N__33035));
    InMux I__7524 (
            .O(N__33089),
            .I(N__33028));
    InMux I__7523 (
            .O(N__33088),
            .I(N__33028));
    InMux I__7522 (
            .O(N__33087),
            .I(N__33028));
    LocalMux I__7521 (
            .O(N__33082),
            .I(N__33019));
    Span4Mux_h I__7520 (
            .O(N__33079),
            .I(N__33019));
    LocalMux I__7519 (
            .O(N__33076),
            .I(N__33019));
    LocalMux I__7518 (
            .O(N__33073),
            .I(N__33019));
    LocalMux I__7517 (
            .O(N__33070),
            .I(N__33016));
    Span4Mux_v I__7516 (
            .O(N__33065),
            .I(N__33013));
    LocalMux I__7515 (
            .O(N__33062),
            .I(N__33008));
    Span4Mux_v I__7514 (
            .O(N__33057),
            .I(N__33008));
    CascadeMux I__7513 (
            .O(N__33056),
            .I(N__33005));
    LocalMux I__7512 (
            .O(N__33053),
            .I(N__33002));
    InMux I__7511 (
            .O(N__33052),
            .I(N__32997));
    InMux I__7510 (
            .O(N__33051),
            .I(N__32997));
    LocalMux I__7509 (
            .O(N__33048),
            .I(N__32994));
    LocalMux I__7508 (
            .O(N__33045),
            .I(N__32985));
    Span4Mux_v I__7507 (
            .O(N__33042),
            .I(N__32985));
    Span4Mux_v I__7506 (
            .O(N__33035),
            .I(N__32985));
    LocalMux I__7505 (
            .O(N__33028),
            .I(N__32985));
    Span4Mux_v I__7504 (
            .O(N__33019),
            .I(N__32976));
    Span4Mux_v I__7503 (
            .O(N__33016),
            .I(N__32976));
    Span4Mux_s0_h I__7502 (
            .O(N__33013),
            .I(N__32976));
    Span4Mux_v I__7501 (
            .O(N__33008),
            .I(N__32976));
    InMux I__7500 (
            .O(N__33005),
            .I(N__32973));
    Odrv4 I__7499 (
            .O(N__33002),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__7498 (
            .O(N__32997),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv12 I__7497 (
            .O(N__32994),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__7496 (
            .O(N__32985),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__7495 (
            .O(N__32976),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__7494 (
            .O(N__32973),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__7493 (
            .O(N__32960),
            .I(N__32954));
    InMux I__7492 (
            .O(N__32959),
            .I(N__32950));
    CascadeMux I__7491 (
            .O(N__32958),
            .I(N__32947));
    CascadeMux I__7490 (
            .O(N__32957),
            .I(N__32943));
    LocalMux I__7489 (
            .O(N__32954),
            .I(N__32937));
    InMux I__7488 (
            .O(N__32953),
            .I(N__32934));
    LocalMux I__7487 (
            .O(N__32950),
            .I(N__32931));
    InMux I__7486 (
            .O(N__32947),
            .I(N__32926));
    InMux I__7485 (
            .O(N__32946),
            .I(N__32926));
    InMux I__7484 (
            .O(N__32943),
            .I(N__32921));
    InMux I__7483 (
            .O(N__32942),
            .I(N__32921));
    InMux I__7482 (
            .O(N__32941),
            .I(N__32916));
    InMux I__7481 (
            .O(N__32940),
            .I(N__32916));
    Span12Mux_s5_v I__7480 (
            .O(N__32937),
            .I(N__32911));
    LocalMux I__7479 (
            .O(N__32934),
            .I(N__32911));
    Odrv4 I__7478 (
            .O(N__32931),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    LocalMux I__7477 (
            .O(N__32926),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    LocalMux I__7476 (
            .O(N__32921),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    LocalMux I__7475 (
            .O(N__32916),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    Odrv12 I__7474 (
            .O(N__32911),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    InMux I__7473 (
            .O(N__32900),
            .I(N__32897));
    LocalMux I__7472 (
            .O(N__32897),
            .I(\POWERLED.g0_i_0_0_0 ));
    InMux I__7471 (
            .O(N__32894),
            .I(N__32891));
    LocalMux I__7470 (
            .O(N__32891),
            .I(N__32888));
    Span4Mux_v I__7469 (
            .O(N__32888),
            .I(N__32885));
    Span4Mux_v I__7468 (
            .O(N__32885),
            .I(N__32882));
    Span4Mux_h I__7467 (
            .O(N__32882),
            .I(N__32877));
    InMux I__7466 (
            .O(N__32881),
            .I(N__32872));
    InMux I__7465 (
            .O(N__32880),
            .I(N__32872));
    Odrv4 I__7464 (
            .O(N__32877),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    LocalMux I__7463 (
            .O(N__32872),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    IoInMux I__7462 (
            .O(N__32867),
            .I(N__32864));
    LocalMux I__7461 (
            .O(N__32864),
            .I(N__32861));
    Span4Mux_s0_h I__7460 (
            .O(N__32861),
            .I(N__32858));
    Odrv4 I__7459 (
            .O(N__32858),
            .I(vpp_en));
    CascadeMux I__7458 (
            .O(N__32855),
            .I(N__32841));
    CascadeMux I__7457 (
            .O(N__32854),
            .I(N__32838));
    CascadeMux I__7456 (
            .O(N__32853),
            .I(N__32833));
    InMux I__7455 (
            .O(N__32852),
            .I(N__32823));
    InMux I__7454 (
            .O(N__32851),
            .I(N__32823));
    InMux I__7453 (
            .O(N__32850),
            .I(N__32823));
    InMux I__7452 (
            .O(N__32849),
            .I(N__32818));
    InMux I__7451 (
            .O(N__32848),
            .I(N__32815));
    InMux I__7450 (
            .O(N__32847),
            .I(N__32807));
    InMux I__7449 (
            .O(N__32846),
            .I(N__32807));
    InMux I__7448 (
            .O(N__32845),
            .I(N__32802));
    InMux I__7447 (
            .O(N__32844),
            .I(N__32802));
    InMux I__7446 (
            .O(N__32841),
            .I(N__32797));
    InMux I__7445 (
            .O(N__32838),
            .I(N__32797));
    InMux I__7444 (
            .O(N__32837),
            .I(N__32790));
    InMux I__7443 (
            .O(N__32836),
            .I(N__32790));
    InMux I__7442 (
            .O(N__32833),
            .I(N__32790));
    InMux I__7441 (
            .O(N__32832),
            .I(N__32783));
    InMux I__7440 (
            .O(N__32831),
            .I(N__32783));
    InMux I__7439 (
            .O(N__32830),
            .I(N__32783));
    LocalMux I__7438 (
            .O(N__32823),
            .I(N__32780));
    CascadeMux I__7437 (
            .O(N__32822),
            .I(N__32777));
    CascadeMux I__7436 (
            .O(N__32821),
            .I(N__32774));
    LocalMux I__7435 (
            .O(N__32818),
            .I(N__32766));
    LocalMux I__7434 (
            .O(N__32815),
            .I(N__32763));
    InMux I__7433 (
            .O(N__32814),
            .I(N__32760));
    InMux I__7432 (
            .O(N__32813),
            .I(N__32757));
    InMux I__7431 (
            .O(N__32812),
            .I(N__32754));
    LocalMux I__7430 (
            .O(N__32807),
            .I(N__32751));
    LocalMux I__7429 (
            .O(N__32802),
            .I(N__32742));
    LocalMux I__7428 (
            .O(N__32797),
            .I(N__32742));
    LocalMux I__7427 (
            .O(N__32790),
            .I(N__32742));
    LocalMux I__7426 (
            .O(N__32783),
            .I(N__32742));
    Span4Mux_h I__7425 (
            .O(N__32780),
            .I(N__32739));
    InMux I__7424 (
            .O(N__32777),
            .I(N__32736));
    InMux I__7423 (
            .O(N__32774),
            .I(N__32731));
    InMux I__7422 (
            .O(N__32773),
            .I(N__32731));
    InMux I__7421 (
            .O(N__32772),
            .I(N__32728));
    InMux I__7420 (
            .O(N__32771),
            .I(N__32721));
    InMux I__7419 (
            .O(N__32770),
            .I(N__32721));
    InMux I__7418 (
            .O(N__32769),
            .I(N__32721));
    Span4Mux_h I__7417 (
            .O(N__32766),
            .I(N__32710));
    Span4Mux_h I__7416 (
            .O(N__32763),
            .I(N__32710));
    LocalMux I__7415 (
            .O(N__32760),
            .I(N__32710));
    LocalMux I__7414 (
            .O(N__32757),
            .I(N__32710));
    LocalMux I__7413 (
            .O(N__32754),
            .I(N__32710));
    Span4Mux_h I__7412 (
            .O(N__32751),
            .I(N__32701));
    Span4Mux_v I__7411 (
            .O(N__32742),
            .I(N__32701));
    Span4Mux_v I__7410 (
            .O(N__32739),
            .I(N__32701));
    LocalMux I__7409 (
            .O(N__32736),
            .I(N__32701));
    LocalMux I__7408 (
            .O(N__32731),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__7407 (
            .O(N__32728),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__7406 (
            .O(N__32721),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__7405 (
            .O(N__32710),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__7404 (
            .O(N__32701),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    InMux I__7403 (
            .O(N__32690),
            .I(N__32687));
    LocalMux I__7402 (
            .O(N__32687),
            .I(N__32684));
    Odrv12 I__7401 (
            .O(N__32684),
            .I(\POWERLED.G_7_i_o5_0 ));
    CascadeMux I__7400 (
            .O(N__32681),
            .I(N__32677));
    CascadeMux I__7399 (
            .O(N__32680),
            .I(N__32671));
    InMux I__7398 (
            .O(N__32677),
            .I(N__32659));
    InMux I__7397 (
            .O(N__32676),
            .I(N__32659));
    InMux I__7396 (
            .O(N__32675),
            .I(N__32659));
    InMux I__7395 (
            .O(N__32674),
            .I(N__32659));
    InMux I__7394 (
            .O(N__32671),
            .I(N__32638));
    InMux I__7393 (
            .O(N__32670),
            .I(N__32638));
    InMux I__7392 (
            .O(N__32669),
            .I(N__32638));
    InMux I__7391 (
            .O(N__32668),
            .I(N__32635));
    LocalMux I__7390 (
            .O(N__32659),
            .I(N__32630));
    InMux I__7389 (
            .O(N__32658),
            .I(N__32625));
    InMux I__7388 (
            .O(N__32657),
            .I(N__32625));
    InMux I__7387 (
            .O(N__32656),
            .I(N__32622));
    InMux I__7386 (
            .O(N__32655),
            .I(N__32615));
    InMux I__7385 (
            .O(N__32654),
            .I(N__32615));
    InMux I__7384 (
            .O(N__32653),
            .I(N__32615));
    InMux I__7383 (
            .O(N__32652),
            .I(N__32612));
    InMux I__7382 (
            .O(N__32651),
            .I(N__32609));
    InMux I__7381 (
            .O(N__32650),
            .I(N__32602));
    InMux I__7380 (
            .O(N__32649),
            .I(N__32602));
    InMux I__7379 (
            .O(N__32648),
            .I(N__32602));
    CascadeMux I__7378 (
            .O(N__32647),
            .I(N__32599));
    CascadeMux I__7377 (
            .O(N__32646),
            .I(N__32595));
    InMux I__7376 (
            .O(N__32645),
            .I(N__32592));
    LocalMux I__7375 (
            .O(N__32638),
            .I(N__32585));
    LocalMux I__7374 (
            .O(N__32635),
            .I(N__32585));
    InMux I__7373 (
            .O(N__32634),
            .I(N__32580));
    InMux I__7372 (
            .O(N__32633),
            .I(N__32580));
    Span4Mux_s2_v I__7371 (
            .O(N__32630),
            .I(N__32573));
    LocalMux I__7370 (
            .O(N__32625),
            .I(N__32573));
    LocalMux I__7369 (
            .O(N__32622),
            .I(N__32570));
    LocalMux I__7368 (
            .O(N__32615),
            .I(N__32567));
    LocalMux I__7367 (
            .O(N__32612),
            .I(N__32560));
    LocalMux I__7366 (
            .O(N__32609),
            .I(N__32560));
    LocalMux I__7365 (
            .O(N__32602),
            .I(N__32560));
    InMux I__7364 (
            .O(N__32599),
            .I(N__32557));
    InMux I__7363 (
            .O(N__32598),
            .I(N__32554));
    InMux I__7362 (
            .O(N__32595),
            .I(N__32551));
    LocalMux I__7361 (
            .O(N__32592),
            .I(N__32548));
    InMux I__7360 (
            .O(N__32591),
            .I(N__32545));
    CascadeMux I__7359 (
            .O(N__32590),
            .I(N__32542));
    Span4Mux_v I__7358 (
            .O(N__32585),
            .I(N__32535));
    LocalMux I__7357 (
            .O(N__32580),
            .I(N__32535));
    InMux I__7356 (
            .O(N__32579),
            .I(N__32530));
    InMux I__7355 (
            .O(N__32578),
            .I(N__32530));
    Span4Mux_v I__7354 (
            .O(N__32573),
            .I(N__32525));
    Span4Mux_v I__7353 (
            .O(N__32570),
            .I(N__32518));
    Span4Mux_h I__7352 (
            .O(N__32567),
            .I(N__32518));
    Span4Mux_v I__7351 (
            .O(N__32560),
            .I(N__32513));
    LocalMux I__7350 (
            .O(N__32557),
            .I(N__32513));
    LocalMux I__7349 (
            .O(N__32554),
            .I(N__32510));
    LocalMux I__7348 (
            .O(N__32551),
            .I(N__32503));
    Span4Mux_v I__7347 (
            .O(N__32548),
            .I(N__32503));
    LocalMux I__7346 (
            .O(N__32545),
            .I(N__32503));
    InMux I__7345 (
            .O(N__32542),
            .I(N__32500));
    InMux I__7344 (
            .O(N__32541),
            .I(N__32497));
    InMux I__7343 (
            .O(N__32540),
            .I(N__32494));
    Span4Mux_h I__7342 (
            .O(N__32535),
            .I(N__32491));
    LocalMux I__7341 (
            .O(N__32530),
            .I(N__32488));
    InMux I__7340 (
            .O(N__32529),
            .I(N__32485));
    InMux I__7339 (
            .O(N__32528),
            .I(N__32480));
    Span4Mux_v I__7338 (
            .O(N__32525),
            .I(N__32477));
    InMux I__7337 (
            .O(N__32524),
            .I(N__32472));
    InMux I__7336 (
            .O(N__32523),
            .I(N__32472));
    Span4Mux_v I__7335 (
            .O(N__32518),
            .I(N__32457));
    Span4Mux_h I__7334 (
            .O(N__32513),
            .I(N__32457));
    Span4Mux_v I__7333 (
            .O(N__32510),
            .I(N__32457));
    Span4Mux_h I__7332 (
            .O(N__32503),
            .I(N__32457));
    LocalMux I__7331 (
            .O(N__32500),
            .I(N__32457));
    LocalMux I__7330 (
            .O(N__32497),
            .I(N__32457));
    LocalMux I__7329 (
            .O(N__32494),
            .I(N__32457));
    Span4Mux_v I__7328 (
            .O(N__32491),
            .I(N__32450));
    Span4Mux_h I__7327 (
            .O(N__32488),
            .I(N__32450));
    LocalMux I__7326 (
            .O(N__32485),
            .I(N__32450));
    InMux I__7325 (
            .O(N__32484),
            .I(N__32445));
    InMux I__7324 (
            .O(N__32483),
            .I(N__32445));
    LocalMux I__7323 (
            .O(N__32480),
            .I(N__32442));
    Sp12to4 I__7322 (
            .O(N__32477),
            .I(N__32437));
    LocalMux I__7321 (
            .O(N__32472),
            .I(N__32437));
    Span4Mux_h I__7320 (
            .O(N__32457),
            .I(N__32434));
    Span4Mux_h I__7319 (
            .O(N__32450),
            .I(N__32431));
    LocalMux I__7318 (
            .O(N__32445),
            .I(N__32428));
    Span12Mux_s8_h I__7317 (
            .O(N__32442),
            .I(N__32425));
    Span12Mux_s8_h I__7316 (
            .O(N__32437),
            .I(N__32420));
    Sp12to4 I__7315 (
            .O(N__32434),
            .I(N__32420));
    Span4Mux_v I__7314 (
            .O(N__32431),
            .I(N__32415));
    Span4Mux_h I__7313 (
            .O(N__32428),
            .I(N__32415));
    Odrv12 I__7312 (
            .O(N__32425),
            .I(slp_s4n));
    Odrv12 I__7311 (
            .O(N__32420),
            .I(slp_s4n));
    Odrv4 I__7310 (
            .O(N__32415),
            .I(slp_s4n));
    InMux I__7309 (
            .O(N__32408),
            .I(N__32403));
    CascadeMux I__7308 (
            .O(N__32407),
            .I(N__32399));
    CascadeMux I__7307 (
            .O(N__32406),
            .I(N__32396));
    LocalMux I__7306 (
            .O(N__32403),
            .I(N__32391));
    CascadeMux I__7305 (
            .O(N__32402),
            .I(N__32388));
    InMux I__7304 (
            .O(N__32399),
            .I(N__32381));
    InMux I__7303 (
            .O(N__32396),
            .I(N__32378));
    InMux I__7302 (
            .O(N__32395),
            .I(N__32372));
    InMux I__7301 (
            .O(N__32394),
            .I(N__32369));
    Span4Mux_v I__7300 (
            .O(N__32391),
            .I(N__32366));
    InMux I__7299 (
            .O(N__32388),
            .I(N__32361));
    InMux I__7298 (
            .O(N__32387),
            .I(N__32361));
    InMux I__7297 (
            .O(N__32386),
            .I(N__32356));
    InMux I__7296 (
            .O(N__32385),
            .I(N__32356));
    CascadeMux I__7295 (
            .O(N__32384),
            .I(N__32353));
    LocalMux I__7294 (
            .O(N__32381),
            .I(N__32347));
    LocalMux I__7293 (
            .O(N__32378),
            .I(N__32347));
    InMux I__7292 (
            .O(N__32377),
            .I(N__32344));
    InMux I__7291 (
            .O(N__32376),
            .I(N__32341));
    InMux I__7290 (
            .O(N__32375),
            .I(N__32338));
    LocalMux I__7289 (
            .O(N__32372),
            .I(N__32333));
    LocalMux I__7288 (
            .O(N__32369),
            .I(N__32333));
    Span4Mux_h I__7287 (
            .O(N__32366),
            .I(N__32328));
    LocalMux I__7286 (
            .O(N__32361),
            .I(N__32328));
    LocalMux I__7285 (
            .O(N__32356),
            .I(N__32325));
    InMux I__7284 (
            .O(N__32353),
            .I(N__32322));
    InMux I__7283 (
            .O(N__32352),
            .I(N__32319));
    Span4Mux_v I__7282 (
            .O(N__32347),
            .I(N__32312));
    LocalMux I__7281 (
            .O(N__32344),
            .I(N__32312));
    LocalMux I__7280 (
            .O(N__32341),
            .I(N__32312));
    LocalMux I__7279 (
            .O(N__32338),
            .I(N__32309));
    Span4Mux_s3_v I__7278 (
            .O(N__32333),
            .I(N__32302));
    Span4Mux_v I__7277 (
            .O(N__32328),
            .I(N__32302));
    Span12Mux_v I__7276 (
            .O(N__32325),
            .I(N__32295));
    LocalMux I__7275 (
            .O(N__32322),
            .I(N__32295));
    LocalMux I__7274 (
            .O(N__32319),
            .I(N__32295));
    Span4Mux_v I__7273 (
            .O(N__32312),
            .I(N__32290));
    Span4Mux_v I__7272 (
            .O(N__32309),
            .I(N__32290));
    InMux I__7271 (
            .O(N__32308),
            .I(N__32285));
    InMux I__7270 (
            .O(N__32307),
            .I(N__32285));
    Odrv4 I__7269 (
            .O(N__32302),
            .I(gpio_fpga_soc_4));
    Odrv12 I__7268 (
            .O(N__32295),
            .I(gpio_fpga_soc_4));
    Odrv4 I__7267 (
            .O(N__32290),
            .I(gpio_fpga_soc_4));
    LocalMux I__7266 (
            .O(N__32285),
            .I(gpio_fpga_soc_4));
    InMux I__7265 (
            .O(N__32276),
            .I(N__32267));
    InMux I__7264 (
            .O(N__32275),
            .I(N__32262));
    InMux I__7263 (
            .O(N__32274),
            .I(N__32262));
    InMux I__7262 (
            .O(N__32273),
            .I(N__32259));
    InMux I__7261 (
            .O(N__32272),
            .I(N__32254));
    CascadeMux I__7260 (
            .O(N__32271),
            .I(N__32251));
    InMux I__7259 (
            .O(N__32270),
            .I(N__32245));
    LocalMux I__7258 (
            .O(N__32267),
            .I(N__32241));
    LocalMux I__7257 (
            .O(N__32262),
            .I(N__32238));
    LocalMux I__7256 (
            .O(N__32259),
            .I(N__32234));
    InMux I__7255 (
            .O(N__32258),
            .I(N__32231));
    InMux I__7254 (
            .O(N__32257),
            .I(N__32225));
    LocalMux I__7253 (
            .O(N__32254),
            .I(N__32222));
    InMux I__7252 (
            .O(N__32251),
            .I(N__32219));
    InMux I__7251 (
            .O(N__32250),
            .I(N__32216));
    CascadeMux I__7250 (
            .O(N__32249),
            .I(N__32212));
    CascadeMux I__7249 (
            .O(N__32248),
            .I(N__32209));
    LocalMux I__7248 (
            .O(N__32245),
            .I(N__32205));
    InMux I__7247 (
            .O(N__32244),
            .I(N__32202));
    Span4Mux_v I__7246 (
            .O(N__32241),
            .I(N__32197));
    Span4Mux_v I__7245 (
            .O(N__32238),
            .I(N__32197));
    CascadeMux I__7244 (
            .O(N__32237),
            .I(N__32194));
    Span4Mux_v I__7243 (
            .O(N__32234),
            .I(N__32187));
    LocalMux I__7242 (
            .O(N__32231),
            .I(N__32187));
    InMux I__7241 (
            .O(N__32230),
            .I(N__32182));
    InMux I__7240 (
            .O(N__32229),
            .I(N__32182));
    InMux I__7239 (
            .O(N__32228),
            .I(N__32179));
    LocalMux I__7238 (
            .O(N__32225),
            .I(N__32172));
    Span4Mux_h I__7237 (
            .O(N__32222),
            .I(N__32172));
    LocalMux I__7236 (
            .O(N__32219),
            .I(N__32172));
    LocalMux I__7235 (
            .O(N__32216),
            .I(N__32169));
    InMux I__7234 (
            .O(N__32215),
            .I(N__32164));
    InMux I__7233 (
            .O(N__32212),
            .I(N__32164));
    InMux I__7232 (
            .O(N__32209),
            .I(N__32159));
    InMux I__7231 (
            .O(N__32208),
            .I(N__32159));
    Span4Mux_v I__7230 (
            .O(N__32205),
            .I(N__32156));
    LocalMux I__7229 (
            .O(N__32202),
            .I(N__32153));
    Span4Mux_h I__7228 (
            .O(N__32197),
            .I(N__32150));
    InMux I__7227 (
            .O(N__32194),
            .I(N__32147));
    InMux I__7226 (
            .O(N__32193),
            .I(N__32144));
    InMux I__7225 (
            .O(N__32192),
            .I(N__32141));
    Span4Mux_h I__7224 (
            .O(N__32187),
            .I(N__32132));
    LocalMux I__7223 (
            .O(N__32182),
            .I(N__32132));
    LocalMux I__7222 (
            .O(N__32179),
            .I(N__32132));
    Span4Mux_h I__7221 (
            .O(N__32172),
            .I(N__32132));
    Span4Mux_v I__7220 (
            .O(N__32169),
            .I(N__32129));
    LocalMux I__7219 (
            .O(N__32164),
            .I(N__32120));
    LocalMux I__7218 (
            .O(N__32159),
            .I(N__32120));
    Span4Mux_h I__7217 (
            .O(N__32156),
            .I(N__32120));
    Span4Mux_s0_h I__7216 (
            .O(N__32153),
            .I(N__32120));
    Odrv4 I__7215 (
            .O(N__32150),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__7214 (
            .O(N__32147),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__7213 (
            .O(N__32144),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__7212 (
            .O(N__32141),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__7211 (
            .O(N__32132),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__7210 (
            .O(N__32129),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__7209 (
            .O(N__32120),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    InMux I__7208 (
            .O(N__32105),
            .I(N__32102));
    LocalMux I__7207 (
            .O(N__32102),
            .I(N__32099));
    Sp12to4 I__7206 (
            .O(N__32099),
            .I(N__32096));
    Odrv12 I__7205 (
            .O(N__32096),
            .I(\POWERLED.dutycycle_e_N_3L4_1 ));
    CascadeMux I__7204 (
            .O(N__32093),
            .I(N__32089));
    CascadeMux I__7203 (
            .O(N__32092),
            .I(N__32086));
    InMux I__7202 (
            .O(N__32089),
            .I(N__32076));
    InMux I__7201 (
            .O(N__32086),
            .I(N__32076));
    InMux I__7200 (
            .O(N__32085),
            .I(N__32071));
    InMux I__7199 (
            .O(N__32084),
            .I(N__32071));
    InMux I__7198 (
            .O(N__32083),
            .I(N__32068));
    InMux I__7197 (
            .O(N__32082),
            .I(N__32065));
    InMux I__7196 (
            .O(N__32081),
            .I(N__32059));
    LocalMux I__7195 (
            .O(N__32076),
            .I(N__32052));
    LocalMux I__7194 (
            .O(N__32071),
            .I(N__32052));
    LocalMux I__7193 (
            .O(N__32068),
            .I(N__32052));
    LocalMux I__7192 (
            .O(N__32065),
            .I(N__32049));
    InMux I__7191 (
            .O(N__32064),
            .I(N__32046));
    InMux I__7190 (
            .O(N__32063),
            .I(N__32041));
    InMux I__7189 (
            .O(N__32062),
            .I(N__32041));
    LocalMux I__7188 (
            .O(N__32059),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    Odrv4 I__7187 (
            .O(N__32052),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    Odrv4 I__7186 (
            .O(N__32049),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    LocalMux I__7185 (
            .O(N__32046),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    LocalMux I__7184 (
            .O(N__32041),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    InMux I__7183 (
            .O(N__32030),
            .I(N__32027));
    LocalMux I__7182 (
            .O(N__32027),
            .I(N__32022));
    CascadeMux I__7181 (
            .O(N__32026),
            .I(N__32018));
    CascadeMux I__7180 (
            .O(N__32025),
            .I(N__32015));
    Span4Mux_s1_v I__7179 (
            .O(N__32022),
            .I(N__32009));
    InMux I__7178 (
            .O(N__32021),
            .I(N__32004));
    InMux I__7177 (
            .O(N__32018),
            .I(N__31998));
    InMux I__7176 (
            .O(N__32015),
            .I(N__31998));
    InMux I__7175 (
            .O(N__32014),
            .I(N__31991));
    InMux I__7174 (
            .O(N__32013),
            .I(N__31991));
    InMux I__7173 (
            .O(N__32012),
            .I(N__31988));
    Span4Mux_v I__7172 (
            .O(N__32009),
            .I(N__31984));
    InMux I__7171 (
            .O(N__32008),
            .I(N__31979));
    InMux I__7170 (
            .O(N__32007),
            .I(N__31979));
    LocalMux I__7169 (
            .O(N__32004),
            .I(N__31976));
    InMux I__7168 (
            .O(N__32003),
            .I(N__31973));
    LocalMux I__7167 (
            .O(N__31998),
            .I(N__31970));
    InMux I__7166 (
            .O(N__31997),
            .I(N__31967));
    InMux I__7165 (
            .O(N__31996),
            .I(N__31964));
    LocalMux I__7164 (
            .O(N__31991),
            .I(N__31959));
    LocalMux I__7163 (
            .O(N__31988),
            .I(N__31959));
    InMux I__7162 (
            .O(N__31987),
            .I(N__31956));
    Sp12to4 I__7161 (
            .O(N__31984),
            .I(N__31950));
    LocalMux I__7160 (
            .O(N__31979),
            .I(N__31947));
    Span4Mux_v I__7159 (
            .O(N__31976),
            .I(N__31944));
    LocalMux I__7158 (
            .O(N__31973),
            .I(N__31941));
    Span4Mux_v I__7157 (
            .O(N__31970),
            .I(N__31932));
    LocalMux I__7156 (
            .O(N__31967),
            .I(N__31932));
    LocalMux I__7155 (
            .O(N__31964),
            .I(N__31932));
    Span4Mux_v I__7154 (
            .O(N__31959),
            .I(N__31932));
    LocalMux I__7153 (
            .O(N__31956),
            .I(N__31929));
    InMux I__7152 (
            .O(N__31955),
            .I(N__31924));
    InMux I__7151 (
            .O(N__31954),
            .I(N__31924));
    InMux I__7150 (
            .O(N__31953),
            .I(N__31921));
    Span12Mux_s8_h I__7149 (
            .O(N__31950),
            .I(N__31916));
    Span12Mux_s3_h I__7148 (
            .O(N__31947),
            .I(N__31916));
    Span4Mux_h I__7147 (
            .O(N__31944),
            .I(N__31913));
    Span4Mux_s1_v I__7146 (
            .O(N__31941),
            .I(N__31910));
    Span4Mux_v I__7145 (
            .O(N__31932),
            .I(N__31903));
    Span4Mux_s0_h I__7144 (
            .O(N__31929),
            .I(N__31903));
    LocalMux I__7143 (
            .O(N__31924),
            .I(N__31903));
    LocalMux I__7142 (
            .O(N__31921),
            .I(VCCST_EN_i_1));
    Odrv12 I__7141 (
            .O(N__31916),
            .I(VCCST_EN_i_1));
    Odrv4 I__7140 (
            .O(N__31913),
            .I(VCCST_EN_i_1));
    Odrv4 I__7139 (
            .O(N__31910),
            .I(VCCST_EN_i_1));
    Odrv4 I__7138 (
            .O(N__31903),
            .I(VCCST_EN_i_1));
    InMux I__7137 (
            .O(N__31892),
            .I(N__31888));
    InMux I__7136 (
            .O(N__31891),
            .I(N__31881));
    LocalMux I__7135 (
            .O(N__31888),
            .I(N__31878));
    InMux I__7134 (
            .O(N__31887),
            .I(N__31875));
    InMux I__7133 (
            .O(N__31886),
            .I(N__31870));
    InMux I__7132 (
            .O(N__31885),
            .I(N__31870));
    CascadeMux I__7131 (
            .O(N__31884),
            .I(N__31865));
    LocalMux I__7130 (
            .O(N__31881),
            .I(N__31861));
    Span4Mux_v I__7129 (
            .O(N__31878),
            .I(N__31856));
    LocalMux I__7128 (
            .O(N__31875),
            .I(N__31856));
    LocalMux I__7127 (
            .O(N__31870),
            .I(N__31853));
    InMux I__7126 (
            .O(N__31869),
            .I(N__31848));
    InMux I__7125 (
            .O(N__31868),
            .I(N__31848));
    InMux I__7124 (
            .O(N__31865),
            .I(N__31845));
    InMux I__7123 (
            .O(N__31864),
            .I(N__31842));
    Span4Mux_s1_h I__7122 (
            .O(N__31861),
            .I(N__31837));
    Span4Mux_h I__7121 (
            .O(N__31856),
            .I(N__31837));
    Odrv4 I__7120 (
            .O(N__31853),
            .I(\POWERLED.N_203 ));
    LocalMux I__7119 (
            .O(N__31848),
            .I(\POWERLED.N_203 ));
    LocalMux I__7118 (
            .O(N__31845),
            .I(\POWERLED.N_203 ));
    LocalMux I__7117 (
            .O(N__31842),
            .I(\POWERLED.N_203 ));
    Odrv4 I__7116 (
            .O(N__31837),
            .I(\POWERLED.N_203 ));
    CascadeMux I__7115 (
            .O(N__31826),
            .I(N__31817));
    CascadeMux I__7114 (
            .O(N__31825),
            .I(N__31814));
    InMux I__7113 (
            .O(N__31824),
            .I(N__31804));
    InMux I__7112 (
            .O(N__31823),
            .I(N__31799));
    InMux I__7111 (
            .O(N__31822),
            .I(N__31799));
    InMux I__7110 (
            .O(N__31821),
            .I(N__31789));
    InMux I__7109 (
            .O(N__31820),
            .I(N__31789));
    InMux I__7108 (
            .O(N__31817),
            .I(N__31789));
    InMux I__7107 (
            .O(N__31814),
            .I(N__31786));
    InMux I__7106 (
            .O(N__31813),
            .I(N__31781));
    InMux I__7105 (
            .O(N__31812),
            .I(N__31781));
    InMux I__7104 (
            .O(N__31811),
            .I(N__31778));
    CascadeMux I__7103 (
            .O(N__31810),
            .I(N__31775));
    CascadeMux I__7102 (
            .O(N__31809),
            .I(N__31770));
    InMux I__7101 (
            .O(N__31808),
            .I(N__31766));
    CascadeMux I__7100 (
            .O(N__31807),
            .I(N__31763));
    LocalMux I__7099 (
            .O(N__31804),
            .I(N__31760));
    LocalMux I__7098 (
            .O(N__31799),
            .I(N__31757));
    CascadeMux I__7097 (
            .O(N__31798),
            .I(N__31753));
    CascadeMux I__7096 (
            .O(N__31797),
            .I(N__31747));
    CascadeMux I__7095 (
            .O(N__31796),
            .I(N__31743));
    LocalMux I__7094 (
            .O(N__31789),
            .I(N__31739));
    LocalMux I__7093 (
            .O(N__31786),
            .I(N__31736));
    LocalMux I__7092 (
            .O(N__31781),
            .I(N__31733));
    LocalMux I__7091 (
            .O(N__31778),
            .I(N__31730));
    InMux I__7090 (
            .O(N__31775),
            .I(N__31723));
    InMux I__7089 (
            .O(N__31774),
            .I(N__31723));
    InMux I__7088 (
            .O(N__31773),
            .I(N__31723));
    InMux I__7087 (
            .O(N__31770),
            .I(N__31718));
    InMux I__7086 (
            .O(N__31769),
            .I(N__31718));
    LocalMux I__7085 (
            .O(N__31766),
            .I(N__31715));
    InMux I__7084 (
            .O(N__31763),
            .I(N__31712));
    Span4Mux_s2_h I__7083 (
            .O(N__31760),
            .I(N__31709));
    Span12Mux_s5_v I__7082 (
            .O(N__31757),
            .I(N__31706));
    InMux I__7081 (
            .O(N__31756),
            .I(N__31701));
    InMux I__7080 (
            .O(N__31753),
            .I(N__31701));
    InMux I__7079 (
            .O(N__31752),
            .I(N__31692));
    InMux I__7078 (
            .O(N__31751),
            .I(N__31692));
    InMux I__7077 (
            .O(N__31750),
            .I(N__31692));
    InMux I__7076 (
            .O(N__31747),
            .I(N__31692));
    InMux I__7075 (
            .O(N__31746),
            .I(N__31685));
    InMux I__7074 (
            .O(N__31743),
            .I(N__31685));
    InMux I__7073 (
            .O(N__31742),
            .I(N__31685));
    Span4Mux_v I__7072 (
            .O(N__31739),
            .I(N__31682));
    Span4Mux_s2_h I__7071 (
            .O(N__31736),
            .I(N__31679));
    Span12Mux_v I__7070 (
            .O(N__31733),
            .I(N__31676));
    Span4Mux_v I__7069 (
            .O(N__31730),
            .I(N__31665));
    LocalMux I__7068 (
            .O(N__31723),
            .I(N__31665));
    LocalMux I__7067 (
            .O(N__31718),
            .I(N__31665));
    Span4Mux_s3_h I__7066 (
            .O(N__31715),
            .I(N__31665));
    LocalMux I__7065 (
            .O(N__31712),
            .I(N__31665));
    Odrv4 I__7064 (
            .O(N__31709),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv12 I__7063 (
            .O(N__31706),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__7062 (
            .O(N__31701),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__7061 (
            .O(N__31692),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__7060 (
            .O(N__31685),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__7059 (
            .O(N__31682),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__7058 (
            .O(N__31679),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv12 I__7057 (
            .O(N__31676),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__7056 (
            .O(N__31665),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    CascadeMux I__7055 (
            .O(N__31646),
            .I(N__31643));
    InMux I__7054 (
            .O(N__31643),
            .I(N__31640));
    LocalMux I__7053 (
            .O(N__31640),
            .I(N__31637));
    Span4Mux_v I__7052 (
            .O(N__31637),
            .I(N__31634));
    Odrv4 I__7051 (
            .O(N__31634),
            .I(\POWERLED.N_505 ));
    CascadeMux I__7050 (
            .O(N__31631),
            .I(\POWERLED.dutycycleZ0Z_8_cascade_ ));
    InMux I__7049 (
            .O(N__31628),
            .I(N__31622));
    InMux I__7048 (
            .O(N__31627),
            .I(N__31622));
    LocalMux I__7047 (
            .O(N__31622),
            .I(\POWERLED.dutycycle_RNIHDMC5Z0Z_3 ));
    InMux I__7046 (
            .O(N__31619),
            .I(N__31615));
    InMux I__7045 (
            .O(N__31618),
            .I(N__31612));
    LocalMux I__7044 (
            .O(N__31615),
            .I(N__31607));
    LocalMux I__7043 (
            .O(N__31612),
            .I(N__31607));
    Span4Mux_s2_h I__7042 (
            .O(N__31607),
            .I(N__31604));
    Odrv4 I__7041 (
            .O(N__31604),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    CascadeMux I__7040 (
            .O(N__31601),
            .I(N__31597));
    InMux I__7039 (
            .O(N__31600),
            .I(N__31592));
    InMux I__7038 (
            .O(N__31597),
            .I(N__31592));
    LocalMux I__7037 (
            .O(N__31592),
            .I(\POWERLED.dutycycleZ1Z_3 ));
    SRMux I__7036 (
            .O(N__31589),
            .I(N__31586));
    LocalMux I__7035 (
            .O(N__31586),
            .I(N__31582));
    SRMux I__7034 (
            .O(N__31585),
            .I(N__31577));
    Span4Mux_h I__7033 (
            .O(N__31582),
            .I(N__31574));
    SRMux I__7032 (
            .O(N__31581),
            .I(N__31571));
    SRMux I__7031 (
            .O(N__31580),
            .I(N__31564));
    LocalMux I__7030 (
            .O(N__31577),
            .I(N__31560));
    IoSpan4Mux I__7029 (
            .O(N__31574),
            .I(N__31557));
    LocalMux I__7028 (
            .O(N__31571),
            .I(N__31553));
    SRMux I__7027 (
            .O(N__31570),
            .I(N__31550));
    SRMux I__7026 (
            .O(N__31569),
            .I(N__31547));
    SRMux I__7025 (
            .O(N__31568),
            .I(N__31544));
    SRMux I__7024 (
            .O(N__31567),
            .I(N__31540));
    LocalMux I__7023 (
            .O(N__31564),
            .I(N__31535));
    SRMux I__7022 (
            .O(N__31563),
            .I(N__31532));
    Span4Mux_h I__7021 (
            .O(N__31560),
            .I(N__31529));
    IoSpan4Mux I__7020 (
            .O(N__31557),
            .I(N__31526));
    SRMux I__7019 (
            .O(N__31556),
            .I(N__31523));
    Span4Mux_s3_h I__7018 (
            .O(N__31553),
            .I(N__31514));
    LocalMux I__7017 (
            .O(N__31550),
            .I(N__31514));
    LocalMux I__7016 (
            .O(N__31547),
            .I(N__31514));
    LocalMux I__7015 (
            .O(N__31544),
            .I(N__31514));
    SRMux I__7014 (
            .O(N__31543),
            .I(N__31511));
    LocalMux I__7013 (
            .O(N__31540),
            .I(N__31508));
    SRMux I__7012 (
            .O(N__31539),
            .I(N__31505));
    SRMux I__7011 (
            .O(N__31538),
            .I(N__31502));
    Span4Mux_v I__7010 (
            .O(N__31535),
            .I(N__31499));
    LocalMux I__7009 (
            .O(N__31532),
            .I(N__31494));
    Span4Mux_v I__7008 (
            .O(N__31529),
            .I(N__31494));
    Span4Mux_s3_h I__7007 (
            .O(N__31526),
            .I(N__31491));
    LocalMux I__7006 (
            .O(N__31523),
            .I(N__31486));
    Span4Mux_v I__7005 (
            .O(N__31514),
            .I(N__31486));
    LocalMux I__7004 (
            .O(N__31511),
            .I(N__31483));
    Span4Mux_v I__7003 (
            .O(N__31508),
            .I(N__31480));
    LocalMux I__7002 (
            .O(N__31505),
            .I(N__31477));
    LocalMux I__7001 (
            .O(N__31502),
            .I(N__31474));
    Span4Mux_v I__7000 (
            .O(N__31499),
            .I(N__31471));
    Span4Mux_v I__6999 (
            .O(N__31494),
            .I(N__31468));
    Sp12to4 I__6998 (
            .O(N__31491),
            .I(N__31465));
    Span4Mux_v I__6997 (
            .O(N__31486),
            .I(N__31462));
    Span4Mux_v I__6996 (
            .O(N__31483),
            .I(N__31455));
    Span4Mux_v I__6995 (
            .O(N__31480),
            .I(N__31455));
    Span4Mux_h I__6994 (
            .O(N__31477),
            .I(N__31455));
    Span4Mux_h I__6993 (
            .O(N__31474),
            .I(N__31452));
    Odrv4 I__6992 (
            .O(N__31471),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv4 I__6991 (
            .O(N__31468),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv12 I__6990 (
            .O(N__31465),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv4 I__6989 (
            .O(N__31462),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv4 I__6988 (
            .O(N__31455),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv4 I__6987 (
            .O(N__31452),
            .I(\POWERLED.N_430_iZ0 ));
    CascadeMux I__6986 (
            .O(N__31439),
            .I(\POWERLED.N_5_0_cascade_ ));
    InMux I__6985 (
            .O(N__31436),
            .I(N__31433));
    LocalMux I__6984 (
            .O(N__31433),
            .I(\POWERLED.N_12_2 ));
    CascadeMux I__6983 (
            .O(N__31430),
            .I(\POWERLED.g0_7_1_cascade_ ));
    InMux I__6982 (
            .O(N__31427),
            .I(N__31424));
    LocalMux I__6981 (
            .O(N__31424),
            .I(N__31421));
    Span4Mux_h I__6980 (
            .O(N__31421),
            .I(N__31418));
    Odrv4 I__6979 (
            .O(N__31418),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_4 ));
    InMux I__6978 (
            .O(N__31415),
            .I(N__31395));
    InMux I__6977 (
            .O(N__31414),
            .I(N__31395));
    InMux I__6976 (
            .O(N__31413),
            .I(N__31388));
    InMux I__6975 (
            .O(N__31412),
            .I(N__31388));
    InMux I__6974 (
            .O(N__31411),
            .I(N__31388));
    InMux I__6973 (
            .O(N__31410),
            .I(N__31383));
    InMux I__6972 (
            .O(N__31409),
            .I(N__31380));
    InMux I__6971 (
            .O(N__31408),
            .I(N__31373));
    InMux I__6970 (
            .O(N__31407),
            .I(N__31373));
    InMux I__6969 (
            .O(N__31406),
            .I(N__31373));
    CascadeMux I__6968 (
            .O(N__31405),
            .I(N__31370));
    InMux I__6967 (
            .O(N__31404),
            .I(N__31367));
    InMux I__6966 (
            .O(N__31403),
            .I(N__31364));
    InMux I__6965 (
            .O(N__31402),
            .I(N__31359));
    InMux I__6964 (
            .O(N__31401),
            .I(N__31359));
    InMux I__6963 (
            .O(N__31400),
            .I(N__31356));
    LocalMux I__6962 (
            .O(N__31395),
            .I(N__31353));
    LocalMux I__6961 (
            .O(N__31388),
            .I(N__31349));
    InMux I__6960 (
            .O(N__31387),
            .I(N__31342));
    InMux I__6959 (
            .O(N__31386),
            .I(N__31337));
    LocalMux I__6958 (
            .O(N__31383),
            .I(N__31334));
    LocalMux I__6957 (
            .O(N__31380),
            .I(N__31329));
    LocalMux I__6956 (
            .O(N__31373),
            .I(N__31329));
    InMux I__6955 (
            .O(N__31370),
            .I(N__31326));
    LocalMux I__6954 (
            .O(N__31367),
            .I(N__31319));
    LocalMux I__6953 (
            .O(N__31364),
            .I(N__31319));
    LocalMux I__6952 (
            .O(N__31359),
            .I(N__31319));
    LocalMux I__6951 (
            .O(N__31356),
            .I(N__31314));
    Span4Mux_v I__6950 (
            .O(N__31353),
            .I(N__31314));
    InMux I__6949 (
            .O(N__31352),
            .I(N__31311));
    Span4Mux_s0_h I__6948 (
            .O(N__31349),
            .I(N__31308));
    InMux I__6947 (
            .O(N__31348),
            .I(N__31303));
    InMux I__6946 (
            .O(N__31347),
            .I(N__31303));
    InMux I__6945 (
            .O(N__31346),
            .I(N__31298));
    InMux I__6944 (
            .O(N__31345),
            .I(N__31298));
    LocalMux I__6943 (
            .O(N__31342),
            .I(N__31295));
    InMux I__6942 (
            .O(N__31341),
            .I(N__31290));
    InMux I__6941 (
            .O(N__31340),
            .I(N__31290));
    LocalMux I__6940 (
            .O(N__31337),
            .I(N__31283));
    Span12Mux_s7_v I__6939 (
            .O(N__31334),
            .I(N__31283));
    Span12Mux_s8_v I__6938 (
            .O(N__31329),
            .I(N__31283));
    LocalMux I__6937 (
            .O(N__31326),
            .I(N__31276));
    Span4Mux_v I__6936 (
            .O(N__31319),
            .I(N__31276));
    Span4Mux_h I__6935 (
            .O(N__31314),
            .I(N__31276));
    LocalMux I__6934 (
            .O(N__31311),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6933 (
            .O(N__31308),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6932 (
            .O(N__31303),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6931 (
            .O(N__31298),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv12 I__6930 (
            .O(N__31295),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6929 (
            .O(N__31290),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv12 I__6928 (
            .O(N__31283),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6927 (
            .O(N__31276),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    InMux I__6926 (
            .O(N__31259),
            .I(N__31249));
    CascadeMux I__6925 (
            .O(N__31258),
            .I(N__31246));
    InMux I__6924 (
            .O(N__31257),
            .I(N__31235));
    InMux I__6923 (
            .O(N__31256),
            .I(N__31235));
    InMux I__6922 (
            .O(N__31255),
            .I(N__31235));
    CascadeMux I__6921 (
            .O(N__31254),
            .I(N__31231));
    CascadeMux I__6920 (
            .O(N__31253),
            .I(N__31227));
    CascadeMux I__6919 (
            .O(N__31252),
            .I(N__31221));
    LocalMux I__6918 (
            .O(N__31249),
            .I(N__31212));
    InMux I__6917 (
            .O(N__31246),
            .I(N__31207));
    InMux I__6916 (
            .O(N__31245),
            .I(N__31207));
    InMux I__6915 (
            .O(N__31244),
            .I(N__31204));
    InMux I__6914 (
            .O(N__31243),
            .I(N__31199));
    InMux I__6913 (
            .O(N__31242),
            .I(N__31199));
    LocalMux I__6912 (
            .O(N__31235),
            .I(N__31196));
    CascadeMux I__6911 (
            .O(N__31234),
            .I(N__31193));
    InMux I__6910 (
            .O(N__31231),
            .I(N__31188));
    InMux I__6909 (
            .O(N__31230),
            .I(N__31188));
    InMux I__6908 (
            .O(N__31227),
            .I(N__31183));
    InMux I__6907 (
            .O(N__31226),
            .I(N__31183));
    InMux I__6906 (
            .O(N__31225),
            .I(N__31176));
    InMux I__6905 (
            .O(N__31224),
            .I(N__31176));
    InMux I__6904 (
            .O(N__31221),
            .I(N__31176));
    InMux I__6903 (
            .O(N__31220),
            .I(N__31173));
    InMux I__6902 (
            .O(N__31219),
            .I(N__31166));
    InMux I__6901 (
            .O(N__31218),
            .I(N__31166));
    InMux I__6900 (
            .O(N__31217),
            .I(N__31166));
    InMux I__6899 (
            .O(N__31216),
            .I(N__31163));
    InMux I__6898 (
            .O(N__31215),
            .I(N__31160));
    Span4Mux_s3_h I__6897 (
            .O(N__31212),
            .I(N__31157));
    LocalMux I__6896 (
            .O(N__31207),
            .I(N__31154));
    LocalMux I__6895 (
            .O(N__31204),
            .I(N__31147));
    LocalMux I__6894 (
            .O(N__31199),
            .I(N__31147));
    Span4Mux_s3_h I__6893 (
            .O(N__31196),
            .I(N__31147));
    InMux I__6892 (
            .O(N__31193),
            .I(N__31144));
    LocalMux I__6891 (
            .O(N__31188),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6890 (
            .O(N__31183),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6889 (
            .O(N__31176),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6888 (
            .O(N__31173),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6887 (
            .O(N__31166),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6886 (
            .O(N__31163),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6885 (
            .O(N__31160),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__6884 (
            .O(N__31157),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__6883 (
            .O(N__31154),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__6882 (
            .O(N__31147),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__6881 (
            .O(N__31144),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    InMux I__6880 (
            .O(N__31121),
            .I(N__31118));
    LocalMux I__6879 (
            .O(N__31118),
            .I(N__31115));
    Span4Mux_v I__6878 (
            .O(N__31115),
            .I(N__31112));
    Odrv4 I__6877 (
            .O(N__31112),
            .I(\POWERLED.i2_mux ));
    InMux I__6876 (
            .O(N__31109),
            .I(N__31101));
    InMux I__6875 (
            .O(N__31108),
            .I(N__31098));
    InMux I__6874 (
            .O(N__31107),
            .I(N__31095));
    InMux I__6873 (
            .O(N__31106),
            .I(N__31090));
    InMux I__6872 (
            .O(N__31105),
            .I(N__31090));
    InMux I__6871 (
            .O(N__31104),
            .I(N__31087));
    LocalMux I__6870 (
            .O(N__31101),
            .I(N__31078));
    LocalMux I__6869 (
            .O(N__31098),
            .I(N__31078));
    LocalMux I__6868 (
            .O(N__31095),
            .I(N__31078));
    LocalMux I__6867 (
            .O(N__31090),
            .I(N__31075));
    LocalMux I__6866 (
            .O(N__31087),
            .I(N__31072));
    InMux I__6865 (
            .O(N__31086),
            .I(N__31069));
    InMux I__6864 (
            .O(N__31085),
            .I(N__31066));
    Span4Mux_v I__6863 (
            .O(N__31078),
            .I(N__31061));
    Span4Mux_s0_h I__6862 (
            .O(N__31075),
            .I(N__31061));
    Odrv4 I__6861 (
            .O(N__31072),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__6860 (
            .O(N__31069),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__6859 (
            .O(N__31066),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    Odrv4 I__6858 (
            .O(N__31061),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    InMux I__6857 (
            .O(N__31052),
            .I(N__31049));
    LocalMux I__6856 (
            .O(N__31049),
            .I(\POWERLED.g1_1cf0 ));
    InMux I__6855 (
            .O(N__31046),
            .I(N__31041));
    InMux I__6854 (
            .O(N__31045),
            .I(N__31036));
    InMux I__6853 (
            .O(N__31044),
            .I(N__31036));
    LocalMux I__6852 (
            .O(N__31041),
            .I(N__31032));
    LocalMux I__6851 (
            .O(N__31036),
            .I(N__31029));
    InMux I__6850 (
            .O(N__31035),
            .I(N__31021));
    Span4Mux_v I__6849 (
            .O(N__31032),
            .I(N__31011));
    Span4Mux_s0_h I__6848 (
            .O(N__31029),
            .I(N__31011));
    InMux I__6847 (
            .O(N__31028),
            .I(N__31008));
    InMux I__6846 (
            .O(N__31027),
            .I(N__31005));
    InMux I__6845 (
            .O(N__31026),
            .I(N__30998));
    InMux I__6844 (
            .O(N__31025),
            .I(N__30998));
    InMux I__6843 (
            .O(N__31024),
            .I(N__30998));
    LocalMux I__6842 (
            .O(N__31021),
            .I(N__30993));
    InMux I__6841 (
            .O(N__31020),
            .I(N__30988));
    InMux I__6840 (
            .O(N__31019),
            .I(N__30988));
    InMux I__6839 (
            .O(N__31018),
            .I(N__30985));
    InMux I__6838 (
            .O(N__31017),
            .I(N__30979));
    InMux I__6837 (
            .O(N__31016),
            .I(N__30979));
    Span4Mux_h I__6836 (
            .O(N__31011),
            .I(N__30972));
    LocalMux I__6835 (
            .O(N__31008),
            .I(N__30972));
    LocalMux I__6834 (
            .O(N__31005),
            .I(N__30972));
    LocalMux I__6833 (
            .O(N__30998),
            .I(N__30969));
    InMux I__6832 (
            .O(N__30997),
            .I(N__30966));
    CascadeMux I__6831 (
            .O(N__30996),
            .I(N__30963));
    Span4Mux_v I__6830 (
            .O(N__30993),
            .I(N__30960));
    LocalMux I__6829 (
            .O(N__30988),
            .I(N__30955));
    LocalMux I__6828 (
            .O(N__30985),
            .I(N__30955));
    InMux I__6827 (
            .O(N__30984),
            .I(N__30952));
    LocalMux I__6826 (
            .O(N__30979),
            .I(N__30943));
    Span4Mux_v I__6825 (
            .O(N__30972),
            .I(N__30943));
    Span4Mux_v I__6824 (
            .O(N__30969),
            .I(N__30943));
    LocalMux I__6823 (
            .O(N__30966),
            .I(N__30943));
    InMux I__6822 (
            .O(N__30963),
            .I(N__30940));
    Odrv4 I__6821 (
            .O(N__30960),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv12 I__6820 (
            .O(N__30955),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__6819 (
            .O(N__30952),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__6818 (
            .O(N__30943),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__6817 (
            .O(N__30940),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    CascadeMux I__6816 (
            .O(N__30929),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_3_cascade_ ));
    CascadeMux I__6815 (
            .O(N__30926),
            .I(N__30923));
    InMux I__6814 (
            .O(N__30923),
            .I(N__30920));
    LocalMux I__6813 (
            .O(N__30920),
            .I(N__30917));
    Span4Mux_v I__6812 (
            .O(N__30917),
            .I(N__30914));
    Span4Mux_h I__6811 (
            .O(N__30914),
            .I(N__30911));
    Odrv4 I__6810 (
            .O(N__30911),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5 ));
    CascadeMux I__6809 (
            .O(N__30908),
            .I(\POWERLED.un1_clk_100khz_32_and_i_0cf0_cascade_ ));
    CascadeMux I__6808 (
            .O(N__30905),
            .I(N__30902));
    InMux I__6807 (
            .O(N__30902),
            .I(N__30895));
    InMux I__6806 (
            .O(N__30901),
            .I(N__30892));
    InMux I__6805 (
            .O(N__30900),
            .I(N__30889));
    InMux I__6804 (
            .O(N__30899),
            .I(N__30886));
    InMux I__6803 (
            .O(N__30898),
            .I(N__30883));
    LocalMux I__6802 (
            .O(N__30895),
            .I(N__30879));
    LocalMux I__6801 (
            .O(N__30892),
            .I(N__30874));
    LocalMux I__6800 (
            .O(N__30889),
            .I(N__30874));
    LocalMux I__6799 (
            .O(N__30886),
            .I(N__30869));
    LocalMux I__6798 (
            .O(N__30883),
            .I(N__30869));
    InMux I__6797 (
            .O(N__30882),
            .I(N__30866));
    Span4Mux_s0_h I__6796 (
            .O(N__30879),
            .I(N__30863));
    Span4Mux_v I__6795 (
            .O(N__30874),
            .I(N__30858));
    Span4Mux_v I__6794 (
            .O(N__30869),
            .I(N__30858));
    LocalMux I__6793 (
            .O(N__30866),
            .I(N__30855));
    Span4Mux_h I__6792 (
            .O(N__30863),
            .I(N__30846));
    Span4Mux_h I__6791 (
            .O(N__30858),
            .I(N__30846));
    Span4Mux_v I__6790 (
            .O(N__30855),
            .I(N__30846));
    InMux I__6789 (
            .O(N__30854),
            .I(N__30843));
    InMux I__6788 (
            .O(N__30853),
            .I(N__30840));
    Odrv4 I__6787 (
            .O(N__30846),
            .I(RSMRSTn_fast));
    LocalMux I__6786 (
            .O(N__30843),
            .I(RSMRSTn_fast));
    LocalMux I__6785 (
            .O(N__30840),
            .I(RSMRSTn_fast));
    CascadeMux I__6784 (
            .O(N__30833),
            .I(N__30829));
    InMux I__6783 (
            .O(N__30832),
            .I(N__30824));
    InMux I__6782 (
            .O(N__30829),
            .I(N__30824));
    LocalMux I__6781 (
            .O(N__30824),
            .I(N__30821));
    Odrv12 I__6780 (
            .O(N__30821),
            .I(\POWERLED.un1_clk_100khz_32_and_i_0 ));
    IoInMux I__6779 (
            .O(N__30818),
            .I(N__30814));
    IoInMux I__6778 (
            .O(N__30817),
            .I(N__30811));
    LocalMux I__6777 (
            .O(N__30814),
            .I(N__30804));
    LocalMux I__6776 (
            .O(N__30811),
            .I(N__30804));
    CascadeMux I__6775 (
            .O(N__30810),
            .I(N__30801));
    InMux I__6774 (
            .O(N__30809),
            .I(N__30791));
    IoSpan4Mux I__6773 (
            .O(N__30804),
            .I(N__30787));
    InMux I__6772 (
            .O(N__30801),
            .I(N__30782));
    InMux I__6771 (
            .O(N__30800),
            .I(N__30782));
    InMux I__6770 (
            .O(N__30799),
            .I(N__30779));
    CascadeMux I__6769 (
            .O(N__30798),
            .I(N__30776));
    CascadeMux I__6768 (
            .O(N__30797),
            .I(N__30773));
    InMux I__6767 (
            .O(N__30796),
            .I(N__30770));
    InMux I__6766 (
            .O(N__30795),
            .I(N__30767));
    InMux I__6765 (
            .O(N__30794),
            .I(N__30764));
    LocalMux I__6764 (
            .O(N__30791),
            .I(N__30761));
    InMux I__6763 (
            .O(N__30790),
            .I(N__30758));
    IoSpan4Mux I__6762 (
            .O(N__30787),
            .I(N__30755));
    LocalMux I__6761 (
            .O(N__30782),
            .I(N__30752));
    LocalMux I__6760 (
            .O(N__30779),
            .I(N__30749));
    InMux I__6759 (
            .O(N__30776),
            .I(N__30746));
    InMux I__6758 (
            .O(N__30773),
            .I(N__30743));
    LocalMux I__6757 (
            .O(N__30770),
            .I(N__30739));
    LocalMux I__6756 (
            .O(N__30767),
            .I(N__30730));
    LocalMux I__6755 (
            .O(N__30764),
            .I(N__30730));
    Span4Mux_v I__6754 (
            .O(N__30761),
            .I(N__30730));
    LocalMux I__6753 (
            .O(N__30758),
            .I(N__30730));
    Span4Mux_s2_h I__6752 (
            .O(N__30755),
            .I(N__30724));
    Span4Mux_v I__6751 (
            .O(N__30752),
            .I(N__30724));
    Span4Mux_h I__6750 (
            .O(N__30749),
            .I(N__30721));
    LocalMux I__6749 (
            .O(N__30746),
            .I(N__30716));
    LocalMux I__6748 (
            .O(N__30743),
            .I(N__30716));
    InMux I__6747 (
            .O(N__30742),
            .I(N__30713));
    Span4Mux_v I__6746 (
            .O(N__30739),
            .I(N__30704));
    Span4Mux_v I__6745 (
            .O(N__30730),
            .I(N__30704));
    InMux I__6744 (
            .O(N__30729),
            .I(N__30701));
    Span4Mux_h I__6743 (
            .O(N__30724),
            .I(N__30698));
    Span4Mux_h I__6742 (
            .O(N__30721),
            .I(N__30691));
    Span4Mux_s3_h I__6741 (
            .O(N__30716),
            .I(N__30691));
    LocalMux I__6740 (
            .O(N__30713),
            .I(N__30691));
    InMux I__6739 (
            .O(N__30712),
            .I(N__30688));
    InMux I__6738 (
            .O(N__30711),
            .I(N__30681));
    InMux I__6737 (
            .O(N__30710),
            .I(N__30681));
    InMux I__6736 (
            .O(N__30709),
            .I(N__30681));
    Span4Mux_h I__6735 (
            .O(N__30704),
            .I(N__30676));
    LocalMux I__6734 (
            .O(N__30701),
            .I(N__30676));
    Odrv4 I__6733 (
            .O(N__30698),
            .I(v5s_enn));
    Odrv4 I__6732 (
            .O(N__30691),
            .I(v5s_enn));
    LocalMux I__6731 (
            .O(N__30688),
            .I(v5s_enn));
    LocalMux I__6730 (
            .O(N__30681),
            .I(v5s_enn));
    Odrv4 I__6729 (
            .O(N__30676),
            .I(v5s_enn));
    CascadeMux I__6728 (
            .O(N__30665),
            .I(N__30654));
    CascadeMux I__6727 (
            .O(N__30664),
            .I(N__30651));
    InMux I__6726 (
            .O(N__30663),
            .I(N__30648));
    InMux I__6725 (
            .O(N__30662),
            .I(N__30645));
    InMux I__6724 (
            .O(N__30661),
            .I(N__30641));
    CascadeMux I__6723 (
            .O(N__30660),
            .I(N__30636));
    CascadeMux I__6722 (
            .O(N__30659),
            .I(N__30633));
    CascadeMux I__6721 (
            .O(N__30658),
            .I(N__30626));
    InMux I__6720 (
            .O(N__30657),
            .I(N__30622));
    InMux I__6719 (
            .O(N__30654),
            .I(N__30617));
    InMux I__6718 (
            .O(N__30651),
            .I(N__30617));
    LocalMux I__6717 (
            .O(N__30648),
            .I(N__30611));
    LocalMux I__6716 (
            .O(N__30645),
            .I(N__30611));
    CascadeMux I__6715 (
            .O(N__30644),
            .I(N__30608));
    LocalMux I__6714 (
            .O(N__30641),
            .I(N__30605));
    InMux I__6713 (
            .O(N__30640),
            .I(N__30602));
    InMux I__6712 (
            .O(N__30639),
            .I(N__30591));
    InMux I__6711 (
            .O(N__30636),
            .I(N__30591));
    InMux I__6710 (
            .O(N__30633),
            .I(N__30591));
    InMux I__6709 (
            .O(N__30632),
            .I(N__30591));
    InMux I__6708 (
            .O(N__30631),
            .I(N__30591));
    InMux I__6707 (
            .O(N__30630),
            .I(N__30586));
    InMux I__6706 (
            .O(N__30629),
            .I(N__30586));
    InMux I__6705 (
            .O(N__30626),
            .I(N__30581));
    InMux I__6704 (
            .O(N__30625),
            .I(N__30581));
    LocalMux I__6703 (
            .O(N__30622),
            .I(N__30578));
    LocalMux I__6702 (
            .O(N__30617),
            .I(N__30571));
    InMux I__6701 (
            .O(N__30616),
            .I(N__30568));
    Span4Mux_v I__6700 (
            .O(N__30611),
            .I(N__30565));
    InMux I__6699 (
            .O(N__30608),
            .I(N__30562));
    Span4Mux_v I__6698 (
            .O(N__30605),
            .I(N__30552));
    LocalMux I__6697 (
            .O(N__30602),
            .I(N__30552));
    LocalMux I__6696 (
            .O(N__30591),
            .I(N__30552));
    LocalMux I__6695 (
            .O(N__30586),
            .I(N__30547));
    LocalMux I__6694 (
            .O(N__30581),
            .I(N__30547));
    Span4Mux_s2_h I__6693 (
            .O(N__30578),
            .I(N__30544));
    CascadeMux I__6692 (
            .O(N__30577),
            .I(N__30541));
    InMux I__6691 (
            .O(N__30576),
            .I(N__30532));
    InMux I__6690 (
            .O(N__30575),
            .I(N__30532));
    InMux I__6689 (
            .O(N__30574),
            .I(N__30532));
    Span4Mux_s2_h I__6688 (
            .O(N__30571),
            .I(N__30529));
    LocalMux I__6687 (
            .O(N__30568),
            .I(N__30526));
    Span4Mux_v I__6686 (
            .O(N__30565),
            .I(N__30523));
    LocalMux I__6685 (
            .O(N__30562),
            .I(N__30520));
    InMux I__6684 (
            .O(N__30561),
            .I(N__30517));
    InMux I__6683 (
            .O(N__30560),
            .I(N__30514));
    InMux I__6682 (
            .O(N__30559),
            .I(N__30511));
    Span4Mux_v I__6681 (
            .O(N__30552),
            .I(N__30508));
    Span4Mux_h I__6680 (
            .O(N__30547),
            .I(N__30503));
    Span4Mux_v I__6679 (
            .O(N__30544),
            .I(N__30503));
    InMux I__6678 (
            .O(N__30541),
            .I(N__30500));
    InMux I__6677 (
            .O(N__30540),
            .I(N__30495));
    InMux I__6676 (
            .O(N__30539),
            .I(N__30495));
    LocalMux I__6675 (
            .O(N__30532),
            .I(N__30488));
    Span4Mux_v I__6674 (
            .O(N__30529),
            .I(N__30488));
    Span4Mux_s2_h I__6673 (
            .O(N__30526),
            .I(N__30488));
    Odrv4 I__6672 (
            .O(N__30523),
            .I(\POWERLED.N_2291_i ));
    Odrv12 I__6671 (
            .O(N__30520),
            .I(\POWERLED.N_2291_i ));
    LocalMux I__6670 (
            .O(N__30517),
            .I(\POWERLED.N_2291_i ));
    LocalMux I__6669 (
            .O(N__30514),
            .I(\POWERLED.N_2291_i ));
    LocalMux I__6668 (
            .O(N__30511),
            .I(\POWERLED.N_2291_i ));
    Odrv4 I__6667 (
            .O(N__30508),
            .I(\POWERLED.N_2291_i ));
    Odrv4 I__6666 (
            .O(N__30503),
            .I(\POWERLED.N_2291_i ));
    LocalMux I__6665 (
            .O(N__30500),
            .I(\POWERLED.N_2291_i ));
    LocalMux I__6664 (
            .O(N__30495),
            .I(\POWERLED.N_2291_i ));
    Odrv4 I__6663 (
            .O(N__30488),
            .I(\POWERLED.N_2291_i ));
    InMux I__6662 (
            .O(N__30467),
            .I(N__30458));
    InMux I__6661 (
            .O(N__30466),
            .I(N__30458));
    InMux I__6660 (
            .O(N__30465),
            .I(N__30458));
    LocalMux I__6659 (
            .O(N__30458),
            .I(N__30455));
    Span4Mux_s3_h I__6658 (
            .O(N__30455),
            .I(N__30452));
    Odrv4 I__6657 (
            .O(N__30452),
            .I(\POWERLED.N_676 ));
    InMux I__6656 (
            .O(N__30449),
            .I(N__30446));
    LocalMux I__6655 (
            .O(N__30446),
            .I(\POWERLED.dutycycle_RNI6SKJ1Z0Z_3 ));
    CascadeMux I__6654 (
            .O(N__30443),
            .I(\POWERLED.func_state_RNILP0FZ0Z_1_cascade_ ));
    InMux I__6653 (
            .O(N__30440),
            .I(N__30437));
    LocalMux I__6652 (
            .O(N__30437),
            .I(\POWERLED.N_523 ));
    CascadeMux I__6651 (
            .O(N__30434),
            .I(N__30431));
    InMux I__6650 (
            .O(N__30431),
            .I(N__30428));
    LocalMux I__6649 (
            .O(N__30428),
            .I(\POWERLED.G_11_i_o10_1_0 ));
    InMux I__6648 (
            .O(N__30425),
            .I(N__30421));
    CascadeMux I__6647 (
            .O(N__30424),
            .I(N__30412));
    LocalMux I__6646 (
            .O(N__30421),
            .I(N__30409));
    InMux I__6645 (
            .O(N__30420),
            .I(N__30406));
    InMux I__6644 (
            .O(N__30419),
            .I(N__30401));
    InMux I__6643 (
            .O(N__30418),
            .I(N__30401));
    InMux I__6642 (
            .O(N__30417),
            .I(N__30397));
    CascadeMux I__6641 (
            .O(N__30416),
            .I(N__30391));
    InMux I__6640 (
            .O(N__30415),
            .I(N__30387));
    InMux I__6639 (
            .O(N__30412),
            .I(N__30384));
    Span4Mux_v I__6638 (
            .O(N__30409),
            .I(N__30381));
    LocalMux I__6637 (
            .O(N__30406),
            .I(N__30378));
    LocalMux I__6636 (
            .O(N__30401),
            .I(N__30375));
    CascadeMux I__6635 (
            .O(N__30400),
            .I(N__30372));
    LocalMux I__6634 (
            .O(N__30397),
            .I(N__30369));
    InMux I__6633 (
            .O(N__30396),
            .I(N__30364));
    InMux I__6632 (
            .O(N__30395),
            .I(N__30364));
    InMux I__6631 (
            .O(N__30394),
            .I(N__30359));
    InMux I__6630 (
            .O(N__30391),
            .I(N__30359));
    InMux I__6629 (
            .O(N__30390),
            .I(N__30355));
    LocalMux I__6628 (
            .O(N__30387),
            .I(N__30350));
    LocalMux I__6627 (
            .O(N__30384),
            .I(N__30350));
    Span4Mux_h I__6626 (
            .O(N__30381),
            .I(N__30345));
    Span4Mux_v I__6625 (
            .O(N__30378),
            .I(N__30345));
    Span4Mux_v I__6624 (
            .O(N__30375),
            .I(N__30342));
    InMux I__6623 (
            .O(N__30372),
            .I(N__30339));
    Sp12to4 I__6622 (
            .O(N__30369),
            .I(N__30332));
    LocalMux I__6621 (
            .O(N__30364),
            .I(N__30332));
    LocalMux I__6620 (
            .O(N__30359),
            .I(N__30332));
    InMux I__6619 (
            .O(N__30358),
            .I(N__30329));
    LocalMux I__6618 (
            .O(N__30355),
            .I(N__30324));
    Span4Mux_v I__6617 (
            .O(N__30350),
            .I(N__30324));
    Odrv4 I__6616 (
            .O(N__30345),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__6615 (
            .O(N__30342),
            .I(\POWERLED.dutycycle ));
    LocalMux I__6614 (
            .O(N__30339),
            .I(\POWERLED.dutycycle ));
    Odrv12 I__6613 (
            .O(N__30332),
            .I(\POWERLED.dutycycle ));
    LocalMux I__6612 (
            .O(N__30329),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__6611 (
            .O(N__30324),
            .I(\POWERLED.dutycycle ));
    InMux I__6610 (
            .O(N__30311),
            .I(N__30307));
    InMux I__6609 (
            .O(N__30310),
            .I(N__30304));
    LocalMux I__6608 (
            .O(N__30307),
            .I(N__30299));
    LocalMux I__6607 (
            .O(N__30304),
            .I(N__30299));
    Odrv4 I__6606 (
            .O(N__30299),
            .I(N_9_0));
    CascadeMux I__6605 (
            .O(N__30296),
            .I(N__30292));
    InMux I__6604 (
            .O(N__30295),
            .I(N__30284));
    InMux I__6603 (
            .O(N__30292),
            .I(N__30284));
    InMux I__6602 (
            .O(N__30291),
            .I(N__30278));
    InMux I__6601 (
            .O(N__30290),
            .I(N__30278));
    InMux I__6600 (
            .O(N__30289),
            .I(N__30272));
    LocalMux I__6599 (
            .O(N__30284),
            .I(N__30268));
    InMux I__6598 (
            .O(N__30283),
            .I(N__30265));
    LocalMux I__6597 (
            .O(N__30278),
            .I(N__30261));
    InMux I__6596 (
            .O(N__30277),
            .I(N__30257));
    InMux I__6595 (
            .O(N__30276),
            .I(N__30252));
    InMux I__6594 (
            .O(N__30275),
            .I(N__30252));
    LocalMux I__6593 (
            .O(N__30272),
            .I(N__30249));
    InMux I__6592 (
            .O(N__30271),
            .I(N__30246));
    Span4Mux_v I__6591 (
            .O(N__30268),
            .I(N__30241));
    LocalMux I__6590 (
            .O(N__30265),
            .I(N__30241));
    InMux I__6589 (
            .O(N__30264),
            .I(N__30238));
    Span12Mux_v I__6588 (
            .O(N__30261),
            .I(N__30235));
    InMux I__6587 (
            .O(N__30260),
            .I(N__30232));
    LocalMux I__6586 (
            .O(N__30257),
            .I(N__30229));
    LocalMux I__6585 (
            .O(N__30252),
            .I(N__30224));
    Span4Mux_s3_h I__6584 (
            .O(N__30249),
            .I(N__30224));
    LocalMux I__6583 (
            .O(N__30246),
            .I(N__30219));
    Span4Mux_v I__6582 (
            .O(N__30241),
            .I(N__30219));
    LocalMux I__6581 (
            .O(N__30238),
            .I(RSMRSTn_rep2));
    Odrv12 I__6580 (
            .O(N__30235),
            .I(RSMRSTn_rep2));
    LocalMux I__6579 (
            .O(N__30232),
            .I(RSMRSTn_rep2));
    Odrv4 I__6578 (
            .O(N__30229),
            .I(RSMRSTn_rep2));
    Odrv4 I__6577 (
            .O(N__30224),
            .I(RSMRSTn_rep2));
    Odrv4 I__6576 (
            .O(N__30219),
            .I(RSMRSTn_rep2));
    CascadeMux I__6575 (
            .O(N__30206),
            .I(N__30201));
    CascadeMux I__6574 (
            .O(N__30205),
            .I(N__30198));
    CascadeMux I__6573 (
            .O(N__30204),
            .I(N__30191));
    InMux I__6572 (
            .O(N__30201),
            .I(N__30188));
    InMux I__6571 (
            .O(N__30198),
            .I(N__30185));
    InMux I__6570 (
            .O(N__30197),
            .I(N__30182));
    InMux I__6569 (
            .O(N__30196),
            .I(N__30179));
    CascadeMux I__6568 (
            .O(N__30195),
            .I(N__30176));
    InMux I__6567 (
            .O(N__30194),
            .I(N__30172));
    InMux I__6566 (
            .O(N__30191),
            .I(N__30169));
    LocalMux I__6565 (
            .O(N__30188),
            .I(N__30166));
    LocalMux I__6564 (
            .O(N__30185),
            .I(N__30163));
    LocalMux I__6563 (
            .O(N__30182),
            .I(N__30160));
    LocalMux I__6562 (
            .O(N__30179),
            .I(N__30157));
    InMux I__6561 (
            .O(N__30176),
            .I(N__30154));
    CascadeMux I__6560 (
            .O(N__30175),
            .I(N__30151));
    LocalMux I__6559 (
            .O(N__30172),
            .I(N__30141));
    LocalMux I__6558 (
            .O(N__30169),
            .I(N__30141));
    Span4Mux_v I__6557 (
            .O(N__30166),
            .I(N__30141));
    Span4Mux_h I__6556 (
            .O(N__30163),
            .I(N__30141));
    Span4Mux_v I__6555 (
            .O(N__30160),
            .I(N__30135));
    Span4Mux_v I__6554 (
            .O(N__30157),
            .I(N__30135));
    LocalMux I__6553 (
            .O(N__30154),
            .I(N__30132));
    InMux I__6552 (
            .O(N__30151),
            .I(N__30127));
    InMux I__6551 (
            .O(N__30150),
            .I(N__30127));
    Span4Mux_v I__6550 (
            .O(N__30141),
            .I(N__30124));
    InMux I__6549 (
            .O(N__30140),
            .I(N__30121));
    Span4Mux_h I__6548 (
            .O(N__30135),
            .I(N__30118));
    Odrv12 I__6547 (
            .O(N__30132),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__6546 (
            .O(N__30127),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__6545 (
            .O(N__30124),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__6544 (
            .O(N__30121),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__6543 (
            .O(N__30118),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__6542 (
            .O(N__30107),
            .I(N__30104));
    LocalMux I__6541 (
            .O(N__30104),
            .I(\POWERLED.N_488 ));
    InMux I__6540 (
            .O(N__30101),
            .I(N__30098));
    LocalMux I__6539 (
            .O(N__30098),
            .I(N__30095));
    Sp12to4 I__6538 (
            .O(N__30095),
            .I(N__30092));
    Odrv12 I__6537 (
            .O(N__30092),
            .I(\POWERLED.N_540_1 ));
    InMux I__6536 (
            .O(N__30089),
            .I(N__30086));
    LocalMux I__6535 (
            .O(N__30086),
            .I(N__30083));
    Span4Mux_h I__6534 (
            .O(N__30083),
            .I(N__30079));
    InMux I__6533 (
            .O(N__30082),
            .I(N__30076));
    Odrv4 I__6532 (
            .O(N__30079),
            .I(POWERLED_un1_dutycycle_172_m0_0));
    LocalMux I__6531 (
            .O(N__30076),
            .I(POWERLED_un1_dutycycle_172_m0_0));
    InMux I__6530 (
            .O(N__30071),
            .I(N__30065));
    InMux I__6529 (
            .O(N__30070),
            .I(N__30062));
    InMux I__6528 (
            .O(N__30069),
            .I(N__30059));
    InMux I__6527 (
            .O(N__30068),
            .I(N__30056));
    LocalMux I__6526 (
            .O(N__30065),
            .I(N__30047));
    LocalMux I__6525 (
            .O(N__30062),
            .I(N__30047));
    LocalMux I__6524 (
            .O(N__30059),
            .I(N__30044));
    LocalMux I__6523 (
            .O(N__30056),
            .I(N__30041));
    InMux I__6522 (
            .O(N__30055),
            .I(N__30034));
    InMux I__6521 (
            .O(N__30054),
            .I(N__30034));
    InMux I__6520 (
            .O(N__30053),
            .I(N__30034));
    InMux I__6519 (
            .O(N__30052),
            .I(N__30030));
    Span4Mux_v I__6518 (
            .O(N__30047),
            .I(N__30027));
    Span4Mux_s2_h I__6517 (
            .O(N__30044),
            .I(N__30024));
    Span4Mux_v I__6516 (
            .O(N__30041),
            .I(N__30019));
    LocalMux I__6515 (
            .O(N__30034),
            .I(N__30019));
    InMux I__6514 (
            .O(N__30033),
            .I(N__30016));
    LocalMux I__6513 (
            .O(N__30030),
            .I(N__30013));
    Odrv4 I__6512 (
            .O(N__30027),
            .I(\POWERLED.N_435 ));
    Odrv4 I__6511 (
            .O(N__30024),
            .I(\POWERLED.N_435 ));
    Odrv4 I__6510 (
            .O(N__30019),
            .I(\POWERLED.N_435 ));
    LocalMux I__6509 (
            .O(N__30016),
            .I(\POWERLED.N_435 ));
    Odrv12 I__6508 (
            .O(N__30013),
            .I(\POWERLED.N_435 ));
    InMux I__6507 (
            .O(N__30002),
            .I(N__29999));
    LocalMux I__6506 (
            .O(N__29999),
            .I(N__29996));
    Span4Mux_v I__6505 (
            .O(N__29996),
            .I(N__29992));
    InMux I__6504 (
            .O(N__29995),
            .I(N__29989));
    Odrv4 I__6503 (
            .O(N__29992),
            .I(\POWERLED.func_state_RNI_4Z0Z_1 ));
    LocalMux I__6502 (
            .O(N__29989),
            .I(\POWERLED.func_state_RNI_4Z0Z_1 ));
    InMux I__6501 (
            .O(N__29984),
            .I(N__29981));
    LocalMux I__6500 (
            .O(N__29981),
            .I(\POWERLED.un1_dutycycle_172_m0_ns_1_0 ));
    CascadeMux I__6499 (
            .O(N__29978),
            .I(\POWERLED.func_state_RNI_4Z0Z_1_cascade_ ));
    InMux I__6498 (
            .O(N__29975),
            .I(N__29972));
    LocalMux I__6497 (
            .O(N__29972),
            .I(\POWERLED.dutycycle_RNI5DLRZ0Z_5 ));
    InMux I__6496 (
            .O(N__29969),
            .I(N__29965));
    InMux I__6495 (
            .O(N__29968),
            .I(N__29962));
    LocalMux I__6494 (
            .O(N__29965),
            .I(N__29955));
    LocalMux I__6493 (
            .O(N__29962),
            .I(N__29952));
    InMux I__6492 (
            .O(N__29961),
            .I(N__29949));
    InMux I__6491 (
            .O(N__29960),
            .I(N__29946));
    InMux I__6490 (
            .O(N__29959),
            .I(N__29940));
    InMux I__6489 (
            .O(N__29958),
            .I(N__29940));
    Span4Mux_v I__6488 (
            .O(N__29955),
            .I(N__29934));
    Span4Mux_s1_h I__6487 (
            .O(N__29952),
            .I(N__29934));
    LocalMux I__6486 (
            .O(N__29949),
            .I(N__29929));
    LocalMux I__6485 (
            .O(N__29946),
            .I(N__29929));
    CascadeMux I__6484 (
            .O(N__29945),
            .I(N__29925));
    LocalMux I__6483 (
            .O(N__29940),
            .I(N__29922));
    InMux I__6482 (
            .O(N__29939),
            .I(N__29919));
    Span4Mux_h I__6481 (
            .O(N__29934),
            .I(N__29916));
    Span12Mux_s7_v I__6480 (
            .O(N__29929),
            .I(N__29913));
    InMux I__6479 (
            .O(N__29928),
            .I(N__29908));
    InMux I__6478 (
            .O(N__29925),
            .I(N__29908));
    Odrv12 I__6477 (
            .O(N__29922),
            .I(SUSWARN_N_rep1));
    LocalMux I__6476 (
            .O(N__29919),
            .I(SUSWARN_N_rep1));
    Odrv4 I__6475 (
            .O(N__29916),
            .I(SUSWARN_N_rep1));
    Odrv12 I__6474 (
            .O(N__29913),
            .I(SUSWARN_N_rep1));
    LocalMux I__6473 (
            .O(N__29908),
            .I(SUSWARN_N_rep1));
    CascadeMux I__6472 (
            .O(N__29897),
            .I(\POWERLED.dutycycle_RNI7ABC3Z0Z_5_cascade_ ));
    CascadeMux I__6471 (
            .O(N__29894),
            .I(N__29890));
    InMux I__6470 (
            .O(N__29893),
            .I(N__29880));
    InMux I__6469 (
            .O(N__29890),
            .I(N__29880));
    InMux I__6468 (
            .O(N__29889),
            .I(N__29877));
    CascadeMux I__6467 (
            .O(N__29888),
            .I(N__29874));
    InMux I__6466 (
            .O(N__29887),
            .I(N__29867));
    InMux I__6465 (
            .O(N__29886),
            .I(N__29867));
    InMux I__6464 (
            .O(N__29885),
            .I(N__29864));
    LocalMux I__6463 (
            .O(N__29880),
            .I(N__29861));
    LocalMux I__6462 (
            .O(N__29877),
            .I(N__29858));
    InMux I__6461 (
            .O(N__29874),
            .I(N__29853));
    InMux I__6460 (
            .O(N__29873),
            .I(N__29853));
    CascadeMux I__6459 (
            .O(N__29872),
            .I(N__29850));
    LocalMux I__6458 (
            .O(N__29867),
            .I(N__29838));
    LocalMux I__6457 (
            .O(N__29864),
            .I(N__29835));
    Span4Mux_v I__6456 (
            .O(N__29861),
            .I(N__29832));
    Span4Mux_h I__6455 (
            .O(N__29858),
            .I(N__29827));
    LocalMux I__6454 (
            .O(N__29853),
            .I(N__29827));
    InMux I__6453 (
            .O(N__29850),
            .I(N__29820));
    InMux I__6452 (
            .O(N__29849),
            .I(N__29820));
    InMux I__6451 (
            .O(N__29848),
            .I(N__29820));
    InMux I__6450 (
            .O(N__29847),
            .I(N__29817));
    InMux I__6449 (
            .O(N__29846),
            .I(N__29812));
    InMux I__6448 (
            .O(N__29845),
            .I(N__29812));
    InMux I__6447 (
            .O(N__29844),
            .I(N__29803));
    InMux I__6446 (
            .O(N__29843),
            .I(N__29803));
    InMux I__6445 (
            .O(N__29842),
            .I(N__29803));
    InMux I__6444 (
            .O(N__29841),
            .I(N__29803));
    Span4Mux_v I__6443 (
            .O(N__29838),
            .I(N__29798));
    Span4Mux_h I__6442 (
            .O(N__29835),
            .I(N__29798));
    Span4Mux_h I__6441 (
            .O(N__29832),
            .I(N__29793));
    Span4Mux_v I__6440 (
            .O(N__29827),
            .I(N__29793));
    LocalMux I__6439 (
            .O(N__29820),
            .I(N__29790));
    LocalMux I__6438 (
            .O(N__29817),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__6437 (
            .O(N__29812),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__6436 (
            .O(N__29803),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__6435 (
            .O(N__29798),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__6434 (
            .O(N__29793),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__6433 (
            .O(N__29790),
            .I(COUNTER_un4_counter_7_THRU_CO));
    InMux I__6432 (
            .O(N__29777),
            .I(N__29774));
    LocalMux I__6431 (
            .O(N__29774),
            .I(N__29771));
    Span4Mux_v I__6430 (
            .O(N__29771),
            .I(N__29768));
    Odrv4 I__6429 (
            .O(N__29768),
            .I(\POWERLED.g2_1_1 ));
    InMux I__6428 (
            .O(N__29765),
            .I(N__29762));
    LocalMux I__6427 (
            .O(N__29762),
            .I(v5s_ok));
    InMux I__6426 (
            .O(N__29759),
            .I(N__29756));
    LocalMux I__6425 (
            .O(N__29756),
            .I(N__29753));
    Span4Mux_v I__6424 (
            .O(N__29753),
            .I(N__29750));
    Odrv4 I__6423 (
            .O(N__29750),
            .I(vccst_cpu_ok));
    CascadeMux I__6422 (
            .O(N__29747),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_1_cascade_ ));
    InMux I__6421 (
            .O(N__29744),
            .I(N__29741));
    LocalMux I__6420 (
            .O(N__29741),
            .I(N__29738));
    Span12Mux_v I__6419 (
            .O(N__29738),
            .I(N__29735));
    Odrv12 I__6418 (
            .O(N__29735),
            .I(v33s_ok));
    IoInMux I__6417 (
            .O(N__29732),
            .I(N__29729));
    LocalMux I__6416 (
            .O(N__29729),
            .I(N__29726));
    Span4Mux_s2_v I__6415 (
            .O(N__29726),
            .I(N__29723));
    Span4Mux_v I__6414 (
            .O(N__29723),
            .I(N__29720));
    Span4Mux_v I__6413 (
            .O(N__29720),
            .I(N__29717));
    Odrv4 I__6412 (
            .O(N__29717),
            .I(vccin_en));
    InMux I__6411 (
            .O(N__29714),
            .I(N__29711));
    LocalMux I__6410 (
            .O(N__29711),
            .I(N__29707));
    InMux I__6409 (
            .O(N__29710),
            .I(N__29704));
    Span4Mux_v I__6408 (
            .O(N__29707),
            .I(N__29698));
    LocalMux I__6407 (
            .O(N__29704),
            .I(N__29698));
    InMux I__6406 (
            .O(N__29703),
            .I(N__29694));
    Span4Mux_h I__6405 (
            .O(N__29698),
            .I(N__29691));
    InMux I__6404 (
            .O(N__29697),
            .I(N__29688));
    LocalMux I__6403 (
            .O(N__29694),
            .I(\POWERLED.N_253 ));
    Odrv4 I__6402 (
            .O(N__29691),
            .I(\POWERLED.N_253 ));
    LocalMux I__6401 (
            .O(N__29688),
            .I(\POWERLED.N_253 ));
    CascadeMux I__6400 (
            .O(N__29681),
            .I(N__29676));
    CascadeMux I__6399 (
            .O(N__29680),
            .I(N__29673));
    InMux I__6398 (
            .O(N__29679),
            .I(N__29669));
    InMux I__6397 (
            .O(N__29676),
            .I(N__29664));
    InMux I__6396 (
            .O(N__29673),
            .I(N__29664));
    InMux I__6395 (
            .O(N__29672),
            .I(N__29661));
    LocalMux I__6394 (
            .O(N__29669),
            .I(N__29658));
    LocalMux I__6393 (
            .O(N__29664),
            .I(N__29653));
    LocalMux I__6392 (
            .O(N__29661),
            .I(N__29653));
    Span4Mux_h I__6391 (
            .O(N__29658),
            .I(N__29650));
    Odrv12 I__6390 (
            .O(N__29653),
            .I(\POWERLED.func_state_RNI_6Z0Z_1 ));
    Odrv4 I__6389 (
            .O(N__29650),
            .I(\POWERLED.func_state_RNI_6Z0Z_1 ));
    InMux I__6388 (
            .O(N__29645),
            .I(N__29642));
    LocalMux I__6387 (
            .O(N__29642),
            .I(N__29638));
    InMux I__6386 (
            .O(N__29641),
            .I(N__29635));
    Odrv12 I__6385 (
            .O(N__29638),
            .I(\POWERLED.g1_1 ));
    LocalMux I__6384 (
            .O(N__29635),
            .I(\POWERLED.g1_1 ));
    CascadeMux I__6383 (
            .O(N__29630),
            .I(\POWERLED.func_state_RNI_6Z0Z_1_cascade_ ));
    CascadeMux I__6382 (
            .O(N__29627),
            .I(\POWERLED.N_2361_0_cascade_ ));
    InMux I__6381 (
            .O(N__29624),
            .I(N__29618));
    InMux I__6380 (
            .O(N__29623),
            .I(N__29618));
    LocalMux I__6379 (
            .O(N__29618),
            .I(N__29615));
    Odrv4 I__6378 (
            .O(N__29615),
            .I(N_6_0));
    InMux I__6377 (
            .O(N__29612),
            .I(N__29609));
    LocalMux I__6376 (
            .O(N__29609),
            .I(\POWERLED.dutycycle_e_N_6L11_1 ));
    CascadeMux I__6375 (
            .O(N__29606),
            .I(\POWERLED.dutycycle_RNI2MQDZ0Z_4_cascade_ ));
    CascadeMux I__6374 (
            .O(N__29603),
            .I(N__29600));
    InMux I__6373 (
            .O(N__29600),
            .I(N__29597));
    LocalMux I__6372 (
            .O(N__29597),
            .I(\POWERLED.dutycycle_RNIOGRSZ0Z_4 ));
    CascadeMux I__6371 (
            .O(N__29594),
            .I(\POWERLED.un1_func_state25_6_0_0_a6_1_0_cascade_ ));
    InMux I__6370 (
            .O(N__29591),
            .I(N__29588));
    LocalMux I__6369 (
            .O(N__29588),
            .I(N__29585));
    Odrv12 I__6368 (
            .O(N__29585),
            .I(\POWERLED.un1_func_state25_6_0_o_N_4 ));
    InMux I__6367 (
            .O(N__29582),
            .I(N__29579));
    LocalMux I__6366 (
            .O(N__29579),
            .I(\POWERLED.un1_func_state25_6_0_0_0_2_1 ));
    CascadeMux I__6365 (
            .O(N__29576),
            .I(\POWERLED.un1_func_state25_6_0_o_N_5_cascade_ ));
    InMux I__6364 (
            .O(N__29573),
            .I(N__29563));
    CascadeMux I__6363 (
            .O(N__29572),
            .I(N__29560));
    CascadeMux I__6362 (
            .O(N__29571),
            .I(N__29556));
    InMux I__6361 (
            .O(N__29570),
            .I(N__29552));
    InMux I__6360 (
            .O(N__29569),
            .I(N__29547));
    InMux I__6359 (
            .O(N__29568),
            .I(N__29547));
    InMux I__6358 (
            .O(N__29567),
            .I(N__29542));
    InMux I__6357 (
            .O(N__29566),
            .I(N__29542));
    LocalMux I__6356 (
            .O(N__29563),
            .I(N__29539));
    InMux I__6355 (
            .O(N__29560),
            .I(N__29535));
    InMux I__6354 (
            .O(N__29559),
            .I(N__29532));
    InMux I__6353 (
            .O(N__29556),
            .I(N__29525));
    InMux I__6352 (
            .O(N__29555),
            .I(N__29525));
    LocalMux I__6351 (
            .O(N__29552),
            .I(N__29522));
    LocalMux I__6350 (
            .O(N__29547),
            .I(N__29517));
    LocalMux I__6349 (
            .O(N__29542),
            .I(N__29517));
    Span4Mux_v I__6348 (
            .O(N__29539),
            .I(N__29514));
    CascadeMux I__6347 (
            .O(N__29538),
            .I(N__29511));
    LocalMux I__6346 (
            .O(N__29535),
            .I(N__29503));
    LocalMux I__6345 (
            .O(N__29532),
            .I(N__29503));
    InMux I__6344 (
            .O(N__29531),
            .I(N__29498));
    InMux I__6343 (
            .O(N__29530),
            .I(N__29498));
    LocalMux I__6342 (
            .O(N__29525),
            .I(N__29495));
    Span4Mux_h I__6341 (
            .O(N__29522),
            .I(N__29492));
    Span4Mux_h I__6340 (
            .O(N__29517),
            .I(N__29487));
    Span4Mux_h I__6339 (
            .O(N__29514),
            .I(N__29487));
    InMux I__6338 (
            .O(N__29511),
            .I(N__29478));
    InMux I__6337 (
            .O(N__29510),
            .I(N__29478));
    InMux I__6336 (
            .O(N__29509),
            .I(N__29478));
    InMux I__6335 (
            .O(N__29508),
            .I(N__29478));
    Odrv12 I__6334 (
            .O(N__29503),
            .I(\POWERLED.N_421 ));
    LocalMux I__6333 (
            .O(N__29498),
            .I(\POWERLED.N_421 ));
    Odrv4 I__6332 (
            .O(N__29495),
            .I(\POWERLED.N_421 ));
    Odrv4 I__6331 (
            .O(N__29492),
            .I(\POWERLED.N_421 ));
    Odrv4 I__6330 (
            .O(N__29487),
            .I(\POWERLED.N_421 ));
    LocalMux I__6329 (
            .O(N__29478),
            .I(\POWERLED.N_421 ));
    CascadeMux I__6328 (
            .O(N__29465),
            .I(\POWERLED.un1_func_state25_6_0_0_0_2_cascade_ ));
    InMux I__6327 (
            .O(N__29462),
            .I(N__29453));
    InMux I__6326 (
            .O(N__29461),
            .I(N__29453));
    CascadeMux I__6325 (
            .O(N__29460),
            .I(N__29449));
    CEMux I__6324 (
            .O(N__29459),
            .I(N__29443));
    InMux I__6323 (
            .O(N__29458),
            .I(N__29440));
    LocalMux I__6322 (
            .O(N__29453),
            .I(N__29437));
    CEMux I__6321 (
            .O(N__29452),
            .I(N__29432));
    InMux I__6320 (
            .O(N__29449),
            .I(N__29423));
    InMux I__6319 (
            .O(N__29448),
            .I(N__29423));
    InMux I__6318 (
            .O(N__29447),
            .I(N__29423));
    InMux I__6317 (
            .O(N__29446),
            .I(N__29423));
    LocalMux I__6316 (
            .O(N__29443),
            .I(N__29420));
    LocalMux I__6315 (
            .O(N__29440),
            .I(N__29417));
    Span4Mux_v I__6314 (
            .O(N__29437),
            .I(N__29414));
    CascadeMux I__6313 (
            .O(N__29436),
            .I(N__29408));
    CascadeMux I__6312 (
            .O(N__29435),
            .I(N__29403));
    LocalMux I__6311 (
            .O(N__29432),
            .I(N__29397));
    LocalMux I__6310 (
            .O(N__29423),
            .I(N__29397));
    Span4Mux_v I__6309 (
            .O(N__29420),
            .I(N__29390));
    Span4Mux_v I__6308 (
            .O(N__29417),
            .I(N__29390));
    Span4Mux_h I__6307 (
            .O(N__29414),
            .I(N__29390));
    CascadeMux I__6306 (
            .O(N__29413),
            .I(N__29386));
    CEMux I__6305 (
            .O(N__29412),
            .I(N__29382));
    CEMux I__6304 (
            .O(N__29411),
            .I(N__29379));
    InMux I__6303 (
            .O(N__29408),
            .I(N__29370));
    InMux I__6302 (
            .O(N__29407),
            .I(N__29370));
    InMux I__6301 (
            .O(N__29406),
            .I(N__29370));
    InMux I__6300 (
            .O(N__29403),
            .I(N__29370));
    InMux I__6299 (
            .O(N__29402),
            .I(N__29364));
    Span4Mux_s3_v I__6298 (
            .O(N__29397),
            .I(N__29359));
    Span4Mux_v I__6297 (
            .O(N__29390),
            .I(N__29359));
    CEMux I__6296 (
            .O(N__29389),
            .I(N__29352));
    InMux I__6295 (
            .O(N__29386),
            .I(N__29352));
    InMux I__6294 (
            .O(N__29385),
            .I(N__29352));
    LocalMux I__6293 (
            .O(N__29382),
            .I(N__29345));
    LocalMux I__6292 (
            .O(N__29379),
            .I(N__29345));
    LocalMux I__6291 (
            .O(N__29370),
            .I(N__29345));
    CEMux I__6290 (
            .O(N__29369),
            .I(N__29338));
    InMux I__6289 (
            .O(N__29368),
            .I(N__29338));
    InMux I__6288 (
            .O(N__29367),
            .I(N__29338));
    LocalMux I__6287 (
            .O(N__29364),
            .I(\POWERLED.func_state_RNI31IBHZ0Z_0 ));
    Odrv4 I__6286 (
            .O(N__29359),
            .I(\POWERLED.func_state_RNI31IBHZ0Z_0 ));
    LocalMux I__6285 (
            .O(N__29352),
            .I(\POWERLED.func_state_RNI31IBHZ0Z_0 ));
    Odrv4 I__6284 (
            .O(N__29345),
            .I(\POWERLED.func_state_RNI31IBHZ0Z_0 ));
    LocalMux I__6283 (
            .O(N__29338),
            .I(\POWERLED.func_state_RNI31IBHZ0Z_0 ));
    InMux I__6282 (
            .O(N__29327),
            .I(N__29324));
    LocalMux I__6281 (
            .O(N__29324),
            .I(N__29321));
    Odrv4 I__6280 (
            .O(N__29321),
            .I(\POWERLED.N_6_2 ));
    InMux I__6279 (
            .O(N__29318),
            .I(N__29315));
    LocalMux I__6278 (
            .O(N__29315),
            .I(N__29311));
    InMux I__6277 (
            .O(N__29314),
            .I(N__29306));
    Span4Mux_v I__6276 (
            .O(N__29311),
            .I(N__29303));
    InMux I__6275 (
            .O(N__29310),
            .I(N__29298));
    InMux I__6274 (
            .O(N__29309),
            .I(N__29298));
    LocalMux I__6273 (
            .O(N__29306),
            .I(N__29295));
    IoSpan4Mux I__6272 (
            .O(N__29303),
            .I(N__29289));
    LocalMux I__6271 (
            .O(N__29298),
            .I(N__29289));
    Span12Mux_v I__6270 (
            .O(N__29295),
            .I(N__29286));
    InMux I__6269 (
            .O(N__29294),
            .I(N__29283));
    Span4Mux_s2_h I__6268 (
            .O(N__29289),
            .I(N__29280));
    Odrv12 I__6267 (
            .O(N__29286),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    LocalMux I__6266 (
            .O(N__29283),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    Odrv4 I__6265 (
            .O(N__29280),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    CascadeMux I__6264 (
            .O(N__29273),
            .I(N__29270));
    InMux I__6263 (
            .O(N__29270),
            .I(N__29267));
    LocalMux I__6262 (
            .O(N__29267),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0 ));
    InMux I__6261 (
            .O(N__29264),
            .I(N__29257));
    InMux I__6260 (
            .O(N__29263),
            .I(N__29254));
    InMux I__6259 (
            .O(N__29262),
            .I(N__29251));
    InMux I__6258 (
            .O(N__29261),
            .I(N__29248));
    CascadeMux I__6257 (
            .O(N__29260),
            .I(N__29242));
    LocalMux I__6256 (
            .O(N__29257),
            .I(N__29235));
    LocalMux I__6255 (
            .O(N__29254),
            .I(N__29235));
    LocalMux I__6254 (
            .O(N__29251),
            .I(N__29232));
    LocalMux I__6253 (
            .O(N__29248),
            .I(N__29229));
    InMux I__6252 (
            .O(N__29247),
            .I(N__29226));
    InMux I__6251 (
            .O(N__29246),
            .I(N__29221));
    InMux I__6250 (
            .O(N__29245),
            .I(N__29221));
    InMux I__6249 (
            .O(N__29242),
            .I(N__29216));
    InMux I__6248 (
            .O(N__29241),
            .I(N__29216));
    InMux I__6247 (
            .O(N__29240),
            .I(N__29213));
    Span4Mux_v I__6246 (
            .O(N__29235),
            .I(N__29208));
    Span4Mux_h I__6245 (
            .O(N__29232),
            .I(N__29208));
    Span4Mux_h I__6244 (
            .O(N__29229),
            .I(N__29205));
    LocalMux I__6243 (
            .O(N__29226),
            .I(N__29202));
    LocalMux I__6242 (
            .O(N__29221),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    LocalMux I__6241 (
            .O(N__29216),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    LocalMux I__6240 (
            .O(N__29213),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__6239 (
            .O(N__29208),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__6238 (
            .O(N__29205),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv12 I__6237 (
            .O(N__29202),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    InMux I__6236 (
            .O(N__29189),
            .I(N__29182));
    InMux I__6235 (
            .O(N__29188),
            .I(N__29177));
    InMux I__6234 (
            .O(N__29187),
            .I(N__29177));
    InMux I__6233 (
            .O(N__29186),
            .I(N__29174));
    InMux I__6232 (
            .O(N__29185),
            .I(N__29171));
    LocalMux I__6231 (
            .O(N__29182),
            .I(N__29168));
    LocalMux I__6230 (
            .O(N__29177),
            .I(N__29165));
    LocalMux I__6229 (
            .O(N__29174),
            .I(N__29160));
    LocalMux I__6228 (
            .O(N__29171),
            .I(N__29160));
    Span4Mux_v I__6227 (
            .O(N__29168),
            .I(N__29157));
    Span12Mux_s7_v I__6226 (
            .O(N__29165),
            .I(N__29154));
    Odrv12 I__6225 (
            .O(N__29160),
            .I(\POWERLED.func_state_RNI_3Z0Z_1 ));
    Odrv4 I__6224 (
            .O(N__29157),
            .I(\POWERLED.func_state_RNI_3Z0Z_1 ));
    Odrv12 I__6223 (
            .O(N__29154),
            .I(\POWERLED.func_state_RNI_3Z0Z_1 ));
    CascadeMux I__6222 (
            .O(N__29147),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0_cascade_ ));
    InMux I__6221 (
            .O(N__29144),
            .I(N__29141));
    LocalMux I__6220 (
            .O(N__29141),
            .I(\POWERLED.func_state_1_m0_1_1 ));
    InMux I__6219 (
            .O(N__29138),
            .I(N__29135));
    LocalMux I__6218 (
            .O(N__29135),
            .I(\POWERLED.un1_func_state25_6_0_o_N_7_2 ));
    InMux I__6217 (
            .O(N__29132),
            .I(N__29127));
    CascadeMux I__6216 (
            .O(N__29131),
            .I(N__29124));
    CascadeMux I__6215 (
            .O(N__29130),
            .I(N__29120));
    LocalMux I__6214 (
            .O(N__29127),
            .I(N__29112));
    InMux I__6213 (
            .O(N__29124),
            .I(N__29103));
    InMux I__6212 (
            .O(N__29123),
            .I(N__29103));
    InMux I__6211 (
            .O(N__29120),
            .I(N__29103));
    InMux I__6210 (
            .O(N__29119),
            .I(N__29103));
    InMux I__6209 (
            .O(N__29118),
            .I(N__29096));
    InMux I__6208 (
            .O(N__29117),
            .I(N__29096));
    InMux I__6207 (
            .O(N__29116),
            .I(N__29096));
    InMux I__6206 (
            .O(N__29115),
            .I(N__29093));
    Span4Mux_v I__6205 (
            .O(N__29112),
            .I(N__29090));
    LocalMux I__6204 (
            .O(N__29103),
            .I(N__29087));
    LocalMux I__6203 (
            .O(N__29096),
            .I(N__29082));
    LocalMux I__6202 (
            .O(N__29093),
            .I(N__29082));
    Span4Mux_h I__6201 (
            .O(N__29090),
            .I(N__29079));
    Span4Mux_h I__6200 (
            .O(N__29087),
            .I(N__29076));
    Span4Mux_h I__6199 (
            .O(N__29082),
            .I(N__29073));
    Odrv4 I__6198 (
            .O(N__29079),
            .I(rsmrst_pwrgd_signal));
    Odrv4 I__6197 (
            .O(N__29076),
            .I(rsmrst_pwrgd_signal));
    Odrv4 I__6196 (
            .O(N__29073),
            .I(rsmrst_pwrgd_signal));
    InMux I__6195 (
            .O(N__29066),
            .I(N__29063));
    LocalMux I__6194 (
            .O(N__29063),
            .I(N__29060));
    Odrv4 I__6193 (
            .O(N__29060),
            .I(\POWERLED.count_off_0_13 ));
    InMux I__6192 (
            .O(N__29057),
            .I(N__29054));
    LocalMux I__6191 (
            .O(N__29054),
            .I(N__29050));
    InMux I__6190 (
            .O(N__29053),
            .I(N__29047));
    Odrv4 I__6189 (
            .O(N__29050),
            .I(\POWERLED.count_off_1_13 ));
    LocalMux I__6188 (
            .O(N__29047),
            .I(\POWERLED.count_off_1_13 ));
    CascadeMux I__6187 (
            .O(N__29042),
            .I(N__29039));
    InMux I__6186 (
            .O(N__29039),
            .I(N__29036));
    LocalMux I__6185 (
            .O(N__29036),
            .I(\POWERLED.count_offZ0Z_13 ));
    CascadeMux I__6184 (
            .O(N__29033),
            .I(N__29029));
    InMux I__6183 (
            .O(N__29032),
            .I(N__29026));
    InMux I__6182 (
            .O(N__29029),
            .I(N__29023));
    LocalMux I__6181 (
            .O(N__29026),
            .I(N__29020));
    LocalMux I__6180 (
            .O(N__29023),
            .I(N__29017));
    Odrv4 I__6179 (
            .O(N__29020),
            .I(\POWERLED.count_offZ0Z_14 ));
    Odrv4 I__6178 (
            .O(N__29017),
            .I(\POWERLED.count_offZ0Z_14 ));
    CascadeMux I__6177 (
            .O(N__29012),
            .I(\POWERLED.count_offZ0Z_13_cascade_ ));
    InMux I__6176 (
            .O(N__29009),
            .I(N__29005));
    InMux I__6175 (
            .O(N__29008),
            .I(N__29002));
    LocalMux I__6174 (
            .O(N__29005),
            .I(N__28999));
    LocalMux I__6173 (
            .O(N__29002),
            .I(N__28996));
    Span4Mux_v I__6172 (
            .O(N__28999),
            .I(N__28993));
    Span4Mux_v I__6171 (
            .O(N__28996),
            .I(N__28990));
    Span4Mux_v I__6170 (
            .O(N__28993),
            .I(N__28985));
    Span4Mux_v I__6169 (
            .O(N__28990),
            .I(N__28985));
    Odrv4 I__6168 (
            .O(N__28985),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__6167 (
            .O(N__28982),
            .I(N__28979));
    LocalMux I__6166 (
            .O(N__28979),
            .I(N__28976));
    Odrv4 I__6165 (
            .O(N__28976),
            .I(\POWERLED.un34_clk_100khz_10 ));
    InMux I__6164 (
            .O(N__28973),
            .I(N__28970));
    LocalMux I__6163 (
            .O(N__28970),
            .I(\POWERLED.count_off_0_0 ));
    CascadeMux I__6162 (
            .O(N__28967),
            .I(\POWERLED.count_off_1_0_cascade_ ));
    CascadeMux I__6161 (
            .O(N__28964),
            .I(N__28958));
    InMux I__6160 (
            .O(N__28963),
            .I(N__28951));
    InMux I__6159 (
            .O(N__28962),
            .I(N__28951));
    InMux I__6158 (
            .O(N__28961),
            .I(N__28951));
    InMux I__6157 (
            .O(N__28958),
            .I(N__28948));
    LocalMux I__6156 (
            .O(N__28951),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__6155 (
            .O(N__28948),
            .I(\POWERLED.count_offZ0Z_0 ));
    CascadeMux I__6154 (
            .O(N__28943),
            .I(\POWERLED.count_offZ0Z_0_cascade_ ));
    InMux I__6153 (
            .O(N__28940),
            .I(N__28937));
    LocalMux I__6152 (
            .O(N__28937),
            .I(\POWERLED.count_off_RNIZ0Z_1 ));
    CascadeMux I__6151 (
            .O(N__28934),
            .I(N__28912));
    InMux I__6150 (
            .O(N__28933),
            .I(N__28905));
    InMux I__6149 (
            .O(N__28932),
            .I(N__28905));
    InMux I__6148 (
            .O(N__28931),
            .I(N__28905));
    InMux I__6147 (
            .O(N__28930),
            .I(N__28900));
    InMux I__6146 (
            .O(N__28929),
            .I(N__28900));
    InMux I__6145 (
            .O(N__28928),
            .I(N__28893));
    InMux I__6144 (
            .O(N__28927),
            .I(N__28893));
    InMux I__6143 (
            .O(N__28926),
            .I(N__28893));
    InMux I__6142 (
            .O(N__28925),
            .I(N__28884));
    InMux I__6141 (
            .O(N__28924),
            .I(N__28884));
    InMux I__6140 (
            .O(N__28923),
            .I(N__28884));
    InMux I__6139 (
            .O(N__28922),
            .I(N__28884));
    InMux I__6138 (
            .O(N__28921),
            .I(N__28875));
    InMux I__6137 (
            .O(N__28920),
            .I(N__28875));
    InMux I__6136 (
            .O(N__28919),
            .I(N__28875));
    InMux I__6135 (
            .O(N__28918),
            .I(N__28875));
    InMux I__6134 (
            .O(N__28917),
            .I(N__28866));
    InMux I__6133 (
            .O(N__28916),
            .I(N__28866));
    InMux I__6132 (
            .O(N__28915),
            .I(N__28866));
    InMux I__6131 (
            .O(N__28912),
            .I(N__28866));
    LocalMux I__6130 (
            .O(N__28905),
            .I(N__28859));
    LocalMux I__6129 (
            .O(N__28900),
            .I(N__28859));
    LocalMux I__6128 (
            .O(N__28893),
            .I(N__28859));
    LocalMux I__6127 (
            .O(N__28884),
            .I(N__28854));
    LocalMux I__6126 (
            .O(N__28875),
            .I(N__28854));
    LocalMux I__6125 (
            .O(N__28866),
            .I(\POWERLED.N_123 ));
    Odrv12 I__6124 (
            .O(N__28859),
            .I(\POWERLED.N_123 ));
    Odrv4 I__6123 (
            .O(N__28854),
            .I(\POWERLED.N_123 ));
    InMux I__6122 (
            .O(N__28847),
            .I(N__28844));
    LocalMux I__6121 (
            .O(N__28844),
            .I(\POWERLED.count_off_0_1 ));
    CascadeMux I__6120 (
            .O(N__28841),
            .I(\POWERLED.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__6119 (
            .O(N__28838),
            .I(N__28834));
    InMux I__6118 (
            .O(N__28837),
            .I(N__28830));
    LocalMux I__6117 (
            .O(N__28834),
            .I(N__28827));
    InMux I__6116 (
            .O(N__28833),
            .I(N__28824));
    LocalMux I__6115 (
            .O(N__28830),
            .I(\POWERLED.count_offZ0Z_1 ));
    Odrv4 I__6114 (
            .O(N__28827),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__6113 (
            .O(N__28824),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__6112 (
            .O(N__28817),
            .I(N__28811));
    InMux I__6111 (
            .O(N__28816),
            .I(N__28811));
    LocalMux I__6110 (
            .O(N__28811),
            .I(\POWERLED.count_off_1_2 ));
    InMux I__6109 (
            .O(N__28808),
            .I(N__28805));
    LocalMux I__6108 (
            .O(N__28805),
            .I(\POWERLED.count_off_0_2 ));
    InMux I__6107 (
            .O(N__28802),
            .I(N__28796));
    InMux I__6106 (
            .O(N__28801),
            .I(N__28796));
    LocalMux I__6105 (
            .O(N__28796),
            .I(\POWERLED.count_off_1_5 ));
    InMux I__6104 (
            .O(N__28793),
            .I(N__28790));
    LocalMux I__6103 (
            .O(N__28790),
            .I(\POWERLED.count_off_0_5 ));
    InMux I__6102 (
            .O(N__28787),
            .I(N__28784));
    LocalMux I__6101 (
            .O(N__28784),
            .I(\POWERLED.count_off_0_6 ));
    InMux I__6100 (
            .O(N__28781),
            .I(N__28775));
    InMux I__6099 (
            .O(N__28780),
            .I(N__28775));
    LocalMux I__6098 (
            .O(N__28775),
            .I(\POWERLED.count_off_1_6 ));
    CascadeMux I__6097 (
            .O(N__28772),
            .I(N__28769));
    InMux I__6096 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__6095 (
            .O(N__28766),
            .I(\POWERLED.count_offZ0Z_6 ));
    CascadeMux I__6094 (
            .O(N__28763),
            .I(N__28759));
    InMux I__6093 (
            .O(N__28762),
            .I(N__28756));
    InMux I__6092 (
            .O(N__28759),
            .I(N__28753));
    LocalMux I__6091 (
            .O(N__28756),
            .I(\POWERLED.count_offZ0Z_5 ));
    LocalMux I__6090 (
            .O(N__28753),
            .I(\POWERLED.count_offZ0Z_5 ));
    CascadeMux I__6089 (
            .O(N__28748),
            .I(N__28744));
    InMux I__6088 (
            .O(N__28747),
            .I(N__28741));
    InMux I__6087 (
            .O(N__28744),
            .I(N__28738));
    LocalMux I__6086 (
            .O(N__28741),
            .I(\POWERLED.count_offZ0Z_2 ));
    LocalMux I__6085 (
            .O(N__28738),
            .I(\POWERLED.count_offZ0Z_2 ));
    CascadeMux I__6084 (
            .O(N__28733),
            .I(\POWERLED.count_offZ0Z_6_cascade_ ));
    InMux I__6083 (
            .O(N__28730),
            .I(N__28727));
    LocalMux I__6082 (
            .O(N__28727),
            .I(N__28724));
    Odrv4 I__6081 (
            .O(N__28724),
            .I(\POWERLED.un34_clk_100khz_9 ));
    InMux I__6080 (
            .O(N__28721),
            .I(N__28718));
    LocalMux I__6079 (
            .O(N__28718),
            .I(\POWERLED.count_off_0_11 ));
    InMux I__6078 (
            .O(N__28715),
            .I(N__28712));
    LocalMux I__6077 (
            .O(N__28712),
            .I(N__28708));
    InMux I__6076 (
            .O(N__28711),
            .I(N__28705));
    Odrv4 I__6075 (
            .O(N__28708),
            .I(\POWERLED.count_off_1_11 ));
    LocalMux I__6074 (
            .O(N__28705),
            .I(\POWERLED.count_off_1_11 ));
    CascadeMux I__6073 (
            .O(N__28700),
            .I(N__28696));
    InMux I__6072 (
            .O(N__28699),
            .I(N__28693));
    InMux I__6071 (
            .O(N__28696),
            .I(N__28690));
    LocalMux I__6070 (
            .O(N__28693),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__6069 (
            .O(N__28690),
            .I(\POWERLED.count_offZ0Z_11 ));
    CascadeMux I__6068 (
            .O(N__28685),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ));
    CascadeMux I__6067 (
            .O(N__28682),
            .I(\POWERLED.count_clkZ0Z_0_cascade_ ));
    CascadeMux I__6066 (
            .O(N__28679),
            .I(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ));
    InMux I__6065 (
            .O(N__28676),
            .I(N__28671));
    InMux I__6064 (
            .O(N__28675),
            .I(N__28666));
    InMux I__6063 (
            .O(N__28674),
            .I(N__28666));
    LocalMux I__6062 (
            .O(N__28671),
            .I(N__28660));
    LocalMux I__6061 (
            .O(N__28666),
            .I(N__28660));
    InMux I__6060 (
            .O(N__28665),
            .I(N__28657));
    Span4Mux_h I__6059 (
            .O(N__28660),
            .I(N__28654));
    LocalMux I__6058 (
            .O(N__28657),
            .I(\POWERLED.count_clkZ0Z_1 ));
    Odrv4 I__6057 (
            .O(N__28654),
            .I(\POWERLED.count_clkZ0Z_1 ));
    CascadeMux I__6056 (
            .O(N__28649),
            .I(\POWERLED.count_clkZ0Z_1_cascade_ ));
    InMux I__6055 (
            .O(N__28646),
            .I(N__28643));
    LocalMux I__6054 (
            .O(N__28643),
            .I(\POWERLED.count_clk_0_1 ));
    InMux I__6053 (
            .O(N__28640),
            .I(N__28637));
    LocalMux I__6052 (
            .O(N__28637),
            .I(N__28633));
    InMux I__6051 (
            .O(N__28636),
            .I(N__28630));
    Span4Mux_s3_v I__6050 (
            .O(N__28633),
            .I(N__28627));
    LocalMux I__6049 (
            .O(N__28630),
            .I(N__28624));
    Odrv4 I__6048 (
            .O(N__28627),
            .I(\POWERLED.count_off_1_14 ));
    Odrv4 I__6047 (
            .O(N__28624),
            .I(\POWERLED.count_off_1_14 ));
    InMux I__6046 (
            .O(N__28619),
            .I(N__28616));
    LocalMux I__6045 (
            .O(N__28616),
            .I(\POWERLED.count_off_0_14 ));
    InMux I__6044 (
            .O(N__28613),
            .I(N__28610));
    LocalMux I__6043 (
            .O(N__28610),
            .I(N__28607));
    Span4Mux_h I__6042 (
            .O(N__28607),
            .I(N__28604));
    Span4Mux_v I__6041 (
            .O(N__28604),
            .I(N__28600));
    InMux I__6040 (
            .O(N__28603),
            .I(N__28597));
    Span4Mux_v I__6039 (
            .O(N__28600),
            .I(N__28594));
    LocalMux I__6038 (
            .O(N__28597),
            .I(\POWERLED.count_off_1_7 ));
    Odrv4 I__6037 (
            .O(N__28594),
            .I(\POWERLED.count_off_1_7 ));
    InMux I__6036 (
            .O(N__28589),
            .I(N__28586));
    LocalMux I__6035 (
            .O(N__28586),
            .I(N__28583));
    Span12Mux_s7_h I__6034 (
            .O(N__28583),
            .I(N__28580));
    Span12Mux_v I__6033 (
            .O(N__28580),
            .I(N__28577));
    Odrv12 I__6032 (
            .O(N__28577),
            .I(\POWERLED.count_off_0_7 ));
    InMux I__6031 (
            .O(N__28574),
            .I(N__28571));
    LocalMux I__6030 (
            .O(N__28571),
            .I(N__28568));
    Span4Mux_h I__6029 (
            .O(N__28568),
            .I(N__28565));
    Span4Mux_v I__6028 (
            .O(N__28565),
            .I(N__28561));
    InMux I__6027 (
            .O(N__28564),
            .I(N__28558));
    Span4Mux_v I__6026 (
            .O(N__28561),
            .I(N__28555));
    LocalMux I__6025 (
            .O(N__28558),
            .I(\POWERLED.count_off_1_8 ));
    Odrv4 I__6024 (
            .O(N__28555),
            .I(\POWERLED.count_off_1_8 ));
    CascadeMux I__6023 (
            .O(N__28550),
            .I(N__28547));
    InMux I__6022 (
            .O(N__28547),
            .I(N__28544));
    LocalMux I__6021 (
            .O(N__28544),
            .I(N__28541));
    Span12Mux_s8_h I__6020 (
            .O(N__28541),
            .I(N__28538));
    Span12Mux_v I__6019 (
            .O(N__28538),
            .I(N__28535));
    Odrv12 I__6018 (
            .O(N__28535),
            .I(\POWERLED.count_off_0_8 ));
    CascadeMux I__6017 (
            .O(N__28532),
            .I(\POWERLED.N_518_cascade_ ));
    InMux I__6016 (
            .O(N__28529),
            .I(N__28522));
    InMux I__6015 (
            .O(N__28528),
            .I(N__28515));
    InMux I__6014 (
            .O(N__28527),
            .I(N__28515));
    InMux I__6013 (
            .O(N__28526),
            .I(N__28515));
    CascadeMux I__6012 (
            .O(N__28525),
            .I(N__28512));
    LocalMux I__6011 (
            .O(N__28522),
            .I(N__28505));
    LocalMux I__6010 (
            .O(N__28515),
            .I(N__28502));
    InMux I__6009 (
            .O(N__28512),
            .I(N__28499));
    InMux I__6008 (
            .O(N__28511),
            .I(N__28496));
    CascadeMux I__6007 (
            .O(N__28510),
            .I(N__28492));
    CascadeMux I__6006 (
            .O(N__28509),
            .I(N__28487));
    InMux I__6005 (
            .O(N__28508),
            .I(N__28484));
    Span12Mux_s7_h I__6004 (
            .O(N__28505),
            .I(N__28481));
    Span4Mux_h I__6003 (
            .O(N__28502),
            .I(N__28476));
    LocalMux I__6002 (
            .O(N__28499),
            .I(N__28476));
    LocalMux I__6001 (
            .O(N__28496),
            .I(N__28473));
    InMux I__6000 (
            .O(N__28495),
            .I(N__28470));
    InMux I__5999 (
            .O(N__28492),
            .I(N__28463));
    InMux I__5998 (
            .O(N__28491),
            .I(N__28463));
    InMux I__5997 (
            .O(N__28490),
            .I(N__28463));
    InMux I__5996 (
            .O(N__28487),
            .I(N__28460));
    LocalMux I__5995 (
            .O(N__28484),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv12 I__5994 (
            .O(N__28481),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5993 (
            .O(N__28476),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5992 (
            .O(N__28473),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__5991 (
            .O(N__28470),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__5990 (
            .O(N__28463),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__5989 (
            .O(N__28460),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    InMux I__5988 (
            .O(N__28445),
            .I(N__28442));
    LocalMux I__5987 (
            .O(N__28442),
            .I(\POWERLED.dutycycle_RNIE3861_0Z0Z_12 ));
    CascadeMux I__5986 (
            .O(N__28439),
            .I(\POWERLED.N_520_cascade_ ));
    InMux I__5985 (
            .O(N__28436),
            .I(N__28430));
    InMux I__5984 (
            .O(N__28435),
            .I(N__28430));
    LocalMux I__5983 (
            .O(N__28430),
            .I(N__28427));
    Span4Mux_h I__5982 (
            .O(N__28427),
            .I(N__28424));
    Odrv4 I__5981 (
            .O(N__28424),
            .I(\POWERLED.dutycycle_RNIPK9V4Z0Z_12 ));
    InMux I__5980 (
            .O(N__28421),
            .I(N__28417));
    InMux I__5979 (
            .O(N__28420),
            .I(N__28414));
    LocalMux I__5978 (
            .O(N__28417),
            .I(N__28409));
    LocalMux I__5977 (
            .O(N__28414),
            .I(N__28409));
    Span12Mux_s6_v I__5976 (
            .O(N__28409),
            .I(N__28406));
    Odrv12 I__5975 (
            .O(N__28406),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIN405GZ0 ));
    InMux I__5974 (
            .O(N__28403),
            .I(N__28400));
    LocalMux I__5973 (
            .O(N__28400),
            .I(\POWERLED.count_off_0_15 ));
    CascadeMux I__5972 (
            .O(N__28397),
            .I(N__28394));
    InMux I__5971 (
            .O(N__28394),
            .I(N__28391));
    LocalMux I__5970 (
            .O(N__28391),
            .I(N__28388));
    Span4Mux_v I__5969 (
            .O(N__28388),
            .I(N__28385));
    Span4Mux_v I__5968 (
            .O(N__28385),
            .I(N__28381));
    InMux I__5967 (
            .O(N__28384),
            .I(N__28378));
    Odrv4 I__5966 (
            .O(N__28381),
            .I(\POWERLED.count_off_RNI8AQHZ0Z_10 ));
    LocalMux I__5965 (
            .O(N__28378),
            .I(\POWERLED.count_off_RNI8AQHZ0Z_10 ));
    InMux I__5964 (
            .O(N__28373),
            .I(N__28370));
    LocalMux I__5963 (
            .O(N__28370),
            .I(N__28367));
    Odrv12 I__5962 (
            .O(N__28367),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_5 ));
    InMux I__5961 (
            .O(N__28364),
            .I(N__28360));
    InMux I__5960 (
            .O(N__28363),
            .I(N__28357));
    LocalMux I__5959 (
            .O(N__28360),
            .I(N__28352));
    LocalMux I__5958 (
            .O(N__28357),
            .I(N__28352));
    Odrv12 I__5957 (
            .O(N__28352),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__5956 (
            .O(N__28349),
            .I(N__28343));
    InMux I__5955 (
            .O(N__28348),
            .I(N__28343));
    LocalMux I__5954 (
            .O(N__28343),
            .I(N__28340));
    Odrv12 I__5953 (
            .O(N__28340),
            .I(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ));
    CascadeMux I__5952 (
            .O(N__28337),
            .I(N__28334));
    InMux I__5951 (
            .O(N__28334),
            .I(N__28331));
    LocalMux I__5950 (
            .O(N__28331),
            .I(\POWERLED.count_clk_0_11 ));
    CascadeMux I__5949 (
            .O(N__28328),
            .I(\POWERLED.N_514_cascade_ ));
    InMux I__5948 (
            .O(N__28325),
            .I(N__28319));
    InMux I__5947 (
            .O(N__28324),
            .I(N__28319));
    LocalMux I__5946 (
            .O(N__28319),
            .I(N__28316));
    Span4Mux_h I__5945 (
            .O(N__28316),
            .I(N__28313));
    Odrv4 I__5944 (
            .O(N__28313),
            .I(\POWERLED.dutycycle_RNIHDMC5Z0Z_11 ));
    InMux I__5943 (
            .O(N__28310),
            .I(N__28305));
    InMux I__5942 (
            .O(N__28309),
            .I(N__28299));
    CascadeMux I__5941 (
            .O(N__28308),
            .I(N__28295));
    LocalMux I__5940 (
            .O(N__28305),
            .I(N__28292));
    InMux I__5939 (
            .O(N__28304),
            .I(N__28285));
    InMux I__5938 (
            .O(N__28303),
            .I(N__28285));
    InMux I__5937 (
            .O(N__28302),
            .I(N__28285));
    LocalMux I__5936 (
            .O(N__28299),
            .I(N__28281));
    CascadeMux I__5935 (
            .O(N__28298),
            .I(N__28275));
    InMux I__5934 (
            .O(N__28295),
            .I(N__28268));
    Span4Mux_v I__5933 (
            .O(N__28292),
            .I(N__28265));
    LocalMux I__5932 (
            .O(N__28285),
            .I(N__28262));
    InMux I__5931 (
            .O(N__28284),
            .I(N__28259));
    Span4Mux_h I__5930 (
            .O(N__28281),
            .I(N__28256));
    InMux I__5929 (
            .O(N__28280),
            .I(N__28251));
    InMux I__5928 (
            .O(N__28279),
            .I(N__28251));
    InMux I__5927 (
            .O(N__28278),
            .I(N__28246));
    InMux I__5926 (
            .O(N__28275),
            .I(N__28246));
    InMux I__5925 (
            .O(N__28274),
            .I(N__28241));
    InMux I__5924 (
            .O(N__28273),
            .I(N__28241));
    InMux I__5923 (
            .O(N__28272),
            .I(N__28236));
    InMux I__5922 (
            .O(N__28271),
            .I(N__28236));
    LocalMux I__5921 (
            .O(N__28268),
            .I(N__28233));
    Odrv4 I__5920 (
            .O(N__28265),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv12 I__5919 (
            .O(N__28262),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__5918 (
            .O(N__28259),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__5917 (
            .O(N__28256),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__5916 (
            .O(N__28251),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__5915 (
            .O(N__28246),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__5914 (
            .O(N__28241),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__5913 (
            .O(N__28236),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__5912 (
            .O(N__28233),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    InMux I__5911 (
            .O(N__28214),
            .I(N__28211));
    LocalMux I__5910 (
            .O(N__28211),
            .I(N__28208));
    Odrv12 I__5909 (
            .O(N__28208),
            .I(\POWERLED.N_508 ));
    CascadeMux I__5908 (
            .O(N__28205),
            .I(\POWERLED.N_512_cascade_ ));
    InMux I__5907 (
            .O(N__28202),
            .I(N__28195));
    InMux I__5906 (
            .O(N__28201),
            .I(N__28190));
    InMux I__5905 (
            .O(N__28200),
            .I(N__28190));
    InMux I__5904 (
            .O(N__28199),
            .I(N__28187));
    InMux I__5903 (
            .O(N__28198),
            .I(N__28184));
    LocalMux I__5902 (
            .O(N__28195),
            .I(N__28176));
    LocalMux I__5901 (
            .O(N__28190),
            .I(N__28171));
    LocalMux I__5900 (
            .O(N__28187),
            .I(N__28171));
    LocalMux I__5899 (
            .O(N__28184),
            .I(N__28168));
    CascadeMux I__5898 (
            .O(N__28183),
            .I(N__28159));
    CascadeMux I__5897 (
            .O(N__28182),
            .I(N__28156));
    InMux I__5896 (
            .O(N__28181),
            .I(N__28151));
    InMux I__5895 (
            .O(N__28180),
            .I(N__28151));
    CascadeMux I__5894 (
            .O(N__28179),
            .I(N__28148));
    Span4Mux_v I__5893 (
            .O(N__28176),
            .I(N__28141));
    Span4Mux_v I__5892 (
            .O(N__28171),
            .I(N__28141));
    Span4Mux_v I__5891 (
            .O(N__28168),
            .I(N__28141));
    InMux I__5890 (
            .O(N__28167),
            .I(N__28136));
    InMux I__5889 (
            .O(N__28166),
            .I(N__28136));
    InMux I__5888 (
            .O(N__28165),
            .I(N__28131));
    InMux I__5887 (
            .O(N__28164),
            .I(N__28131));
    InMux I__5886 (
            .O(N__28163),
            .I(N__28122));
    InMux I__5885 (
            .O(N__28162),
            .I(N__28122));
    InMux I__5884 (
            .O(N__28159),
            .I(N__28122));
    InMux I__5883 (
            .O(N__28156),
            .I(N__28122));
    LocalMux I__5882 (
            .O(N__28151),
            .I(N__28119));
    InMux I__5881 (
            .O(N__28148),
            .I(N__28116));
    Odrv4 I__5880 (
            .O(N__28141),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__5879 (
            .O(N__28136),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__5878 (
            .O(N__28131),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__5877 (
            .O(N__28122),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__5876 (
            .O(N__28119),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__5875 (
            .O(N__28116),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    InMux I__5874 (
            .O(N__28103),
            .I(N__28100));
    LocalMux I__5873 (
            .O(N__28100),
            .I(\POWERLED.dutycycle_RNI6SKJ1_0Z0Z_11 ));
    CascadeMux I__5872 (
            .O(N__28097),
            .I(\POWERLED.N_526_cascade_ ));
    InMux I__5871 (
            .O(N__28094),
            .I(N__28091));
    LocalMux I__5870 (
            .O(N__28091),
            .I(\POWERLED.un1_clk_100khz_47_and_i_1 ));
    CascadeMux I__5869 (
            .O(N__28088),
            .I(N__28084));
    InMux I__5868 (
            .O(N__28087),
            .I(N__28079));
    InMux I__5867 (
            .O(N__28084),
            .I(N__28079));
    LocalMux I__5866 (
            .O(N__28079),
            .I(N__28076));
    Odrv4 I__5865 (
            .O(N__28076),
            .I(\POWERLED.dutycycle_en_11 ));
    InMux I__5864 (
            .O(N__28073),
            .I(N__28070));
    LocalMux I__5863 (
            .O(N__28070),
            .I(\POWERLED.N_2075_tz_tz ));
    CascadeMux I__5862 (
            .O(N__28067),
            .I(N__28063));
    InMux I__5861 (
            .O(N__28066),
            .I(N__28060));
    InMux I__5860 (
            .O(N__28063),
            .I(N__28057));
    LocalMux I__5859 (
            .O(N__28060),
            .I(N__28052));
    LocalMux I__5858 (
            .O(N__28057),
            .I(N__28049));
    InMux I__5857 (
            .O(N__28056),
            .I(N__28046));
    InMux I__5856 (
            .O(N__28055),
            .I(N__28043));
    Span4Mux_s1_h I__5855 (
            .O(N__28052),
            .I(N__28040));
    Span4Mux_v I__5854 (
            .O(N__28049),
            .I(N__28033));
    LocalMux I__5853 (
            .O(N__28046),
            .I(N__28033));
    LocalMux I__5852 (
            .O(N__28043),
            .I(N__28033));
    Span4Mux_h I__5851 (
            .O(N__28040),
            .I(N__28030));
    Span4Mux_h I__5850 (
            .O(N__28033),
            .I(N__28027));
    Odrv4 I__5849 (
            .O(N__28030),
            .I(\POWERLED.N_600 ));
    Odrv4 I__5848 (
            .O(N__28027),
            .I(\POWERLED.N_600 ));
    InMux I__5847 (
            .O(N__28022),
            .I(N__28019));
    LocalMux I__5846 (
            .O(N__28019),
            .I(N__28016));
    Span4Mux_v I__5845 (
            .O(N__28016),
            .I(N__28013));
    Odrv4 I__5844 (
            .O(N__28013),
            .I(\POWERLED.count_clk_en_0 ));
    CascadeMux I__5843 (
            .O(N__28010),
            .I(N__28007));
    InMux I__5842 (
            .O(N__28007),
            .I(N__28004));
    LocalMux I__5841 (
            .O(N__28004),
            .I(N__28001));
    Odrv4 I__5840 (
            .O(N__28001),
            .I(\POWERLED.N_443 ));
    InMux I__5839 (
            .O(N__27998),
            .I(N__27995));
    LocalMux I__5838 (
            .O(N__27995),
            .I(N__27992));
    Odrv12 I__5837 (
            .O(N__27992),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_1 ));
    CascadeMux I__5836 (
            .O(N__27989),
            .I(\POWERLED.N_443_cascade_ ));
    InMux I__5835 (
            .O(N__27986),
            .I(N__27982));
    InMux I__5834 (
            .O(N__27985),
            .I(N__27978));
    LocalMux I__5833 (
            .O(N__27982),
            .I(N__27975));
    CascadeMux I__5832 (
            .O(N__27981),
            .I(N__27972));
    LocalMux I__5831 (
            .O(N__27978),
            .I(N__27969));
    Span4Mux_v I__5830 (
            .O(N__27975),
            .I(N__27966));
    InMux I__5829 (
            .O(N__27972),
            .I(N__27963));
    Span4Mux_v I__5828 (
            .O(N__27969),
            .I(N__27960));
    Span4Mux_h I__5827 (
            .O(N__27966),
            .I(N__27955));
    LocalMux I__5826 (
            .O(N__27963),
            .I(N__27955));
    Span4Mux_v I__5825 (
            .O(N__27960),
            .I(N__27952));
    Span4Mux_v I__5824 (
            .O(N__27955),
            .I(N__27949));
    Odrv4 I__5823 (
            .O(N__27952),
            .I(\POWERLED.count_clk_RNINSEUCZ0Z_7 ));
    Odrv4 I__5822 (
            .O(N__27949),
            .I(\POWERLED.count_clk_RNINSEUCZ0Z_7 ));
    InMux I__5821 (
            .O(N__27944),
            .I(N__27940));
    CascadeMux I__5820 (
            .O(N__27943),
            .I(N__27937));
    LocalMux I__5819 (
            .O(N__27940),
            .I(N__27934));
    InMux I__5818 (
            .O(N__27937),
            .I(N__27931));
    Span4Mux_v I__5817 (
            .O(N__27934),
            .I(N__27928));
    LocalMux I__5816 (
            .O(N__27931),
            .I(N__27924));
    Span4Mux_v I__5815 (
            .O(N__27928),
            .I(N__27921));
    InMux I__5814 (
            .O(N__27927),
            .I(N__27918));
    Span4Mux_s2_h I__5813 (
            .O(N__27924),
            .I(N__27915));
    IoSpan4Mux I__5812 (
            .O(N__27921),
            .I(N__27910));
    LocalMux I__5811 (
            .O(N__27918),
            .I(N__27910));
    Span4Mux_v I__5810 (
            .O(N__27915),
            .I(N__27905));
    Span4Mux_s2_h I__5809 (
            .O(N__27910),
            .I(N__27905));
    Odrv4 I__5808 (
            .O(N__27905),
            .I(\POWERLED.N_668 ));
    InMux I__5807 (
            .O(N__27902),
            .I(N__27899));
    LocalMux I__5806 (
            .O(N__27899),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_2 ));
    CascadeMux I__5805 (
            .O(N__27896),
            .I(N__27892));
    CascadeMux I__5804 (
            .O(N__27895),
            .I(N__27887));
    InMux I__5803 (
            .O(N__27892),
            .I(N__27883));
    InMux I__5802 (
            .O(N__27891),
            .I(N__27878));
    InMux I__5801 (
            .O(N__27890),
            .I(N__27878));
    InMux I__5800 (
            .O(N__27887),
            .I(N__27875));
    CascadeMux I__5799 (
            .O(N__27886),
            .I(N__27870));
    LocalMux I__5798 (
            .O(N__27883),
            .I(N__27865));
    LocalMux I__5797 (
            .O(N__27878),
            .I(N__27862));
    LocalMux I__5796 (
            .O(N__27875),
            .I(N__27859));
    InMux I__5795 (
            .O(N__27874),
            .I(N__27854));
    InMux I__5794 (
            .O(N__27873),
            .I(N__27854));
    InMux I__5793 (
            .O(N__27870),
            .I(N__27851));
    InMux I__5792 (
            .O(N__27869),
            .I(N__27846));
    InMux I__5791 (
            .O(N__27868),
            .I(N__27846));
    Span4Mux_v I__5790 (
            .O(N__27865),
            .I(N__27843));
    Span4Mux_v I__5789 (
            .O(N__27862),
            .I(N__27838));
    Span4Mux_h I__5788 (
            .O(N__27859),
            .I(N__27838));
    LocalMux I__5787 (
            .O(N__27854),
            .I(N__27833));
    LocalMux I__5786 (
            .O(N__27851),
            .I(N__27833));
    LocalMux I__5785 (
            .O(N__27846),
            .I(N__27830));
    Odrv4 I__5784 (
            .O(N__27843),
            .I(N_247));
    Odrv4 I__5783 (
            .O(N__27838),
            .I(N_247));
    Odrv12 I__5782 (
            .O(N__27833),
            .I(N_247));
    Odrv12 I__5781 (
            .O(N__27830),
            .I(N_247));
    InMux I__5780 (
            .O(N__27821),
            .I(N__27818));
    LocalMux I__5779 (
            .O(N__27818),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_0 ));
    InMux I__5778 (
            .O(N__27815),
            .I(N__27811));
    CascadeMux I__5777 (
            .O(N__27814),
            .I(N__27808));
    LocalMux I__5776 (
            .O(N__27811),
            .I(N__27803));
    InMux I__5775 (
            .O(N__27808),
            .I(N__27800));
    InMux I__5774 (
            .O(N__27807),
            .I(N__27792));
    InMux I__5773 (
            .O(N__27806),
            .I(N__27792));
    Span4Mux_h I__5772 (
            .O(N__27803),
            .I(N__27787));
    LocalMux I__5771 (
            .O(N__27800),
            .I(N__27787));
    CascadeMux I__5770 (
            .O(N__27799),
            .I(N__27784));
    CascadeMux I__5769 (
            .O(N__27798),
            .I(N__27781));
    InMux I__5768 (
            .O(N__27797),
            .I(N__27778));
    LocalMux I__5767 (
            .O(N__27792),
            .I(N__27775));
    Span4Mux_v I__5766 (
            .O(N__27787),
            .I(N__27772));
    InMux I__5765 (
            .O(N__27784),
            .I(N__27767));
    InMux I__5764 (
            .O(N__27781),
            .I(N__27767));
    LocalMux I__5763 (
            .O(N__27778),
            .I(RSMRSTn_rep1));
    Odrv4 I__5762 (
            .O(N__27775),
            .I(RSMRSTn_rep1));
    Odrv4 I__5761 (
            .O(N__27772),
            .I(RSMRSTn_rep1));
    LocalMux I__5760 (
            .O(N__27767),
            .I(RSMRSTn_rep1));
    CascadeMux I__5759 (
            .O(N__27758),
            .I(\POWERLED.N_506_cascade_ ));
    CascadeMux I__5758 (
            .O(N__27755),
            .I(N__27752));
    InMux I__5757 (
            .O(N__27752),
            .I(N__27749));
    LocalMux I__5756 (
            .O(N__27749),
            .I(N__27746));
    Span4Mux_h I__5755 (
            .O(N__27746),
            .I(N__27743));
    Odrv4 I__5754 (
            .O(N__27743),
            .I(\POWERLED.dutycycle_RNI6SKJ1_0Z0Z_10 ));
    InMux I__5753 (
            .O(N__27740),
            .I(N__27737));
    LocalMux I__5752 (
            .O(N__27737),
            .I(N__27734));
    Span4Mux_h I__5751 (
            .O(N__27734),
            .I(N__27731));
    Odrv4 I__5750 (
            .O(N__27731),
            .I(\POWERLED.g0_i_0_1 ));
    CascadeMux I__5749 (
            .O(N__27728),
            .I(\POWERLED.un1_dutycycle_53_25_0_tz_1_1_cascade_ ));
    InMux I__5748 (
            .O(N__27725),
            .I(N__27721));
    InMux I__5747 (
            .O(N__27724),
            .I(N__27718));
    LocalMux I__5746 (
            .O(N__27721),
            .I(N__27713));
    LocalMux I__5745 (
            .O(N__27718),
            .I(N__27713));
    Span4Mux_h I__5744 (
            .O(N__27713),
            .I(N__27710));
    Odrv4 I__5743 (
            .O(N__27710),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_4 ));
    CascadeMux I__5742 (
            .O(N__27707),
            .I(N__27704));
    InMux I__5741 (
            .O(N__27704),
            .I(N__27700));
    InMux I__5740 (
            .O(N__27703),
            .I(N__27697));
    LocalMux I__5739 (
            .O(N__27700),
            .I(N__27694));
    LocalMux I__5738 (
            .O(N__27697),
            .I(N__27689));
    Span4Mux_s2_h I__5737 (
            .O(N__27694),
            .I(N__27689));
    Span4Mux_v I__5736 (
            .O(N__27689),
            .I(N__27686));
    Odrv4 I__5735 (
            .O(N__27686),
            .I(\POWERLED.func_state_RNI_0Z0Z_1 ));
    InMux I__5734 (
            .O(N__27683),
            .I(N__27678));
    InMux I__5733 (
            .O(N__27682),
            .I(N__27673));
    CascadeMux I__5732 (
            .O(N__27681),
            .I(N__27670));
    LocalMux I__5731 (
            .O(N__27678),
            .I(N__27667));
    InMux I__5730 (
            .O(N__27677),
            .I(N__27662));
    InMux I__5729 (
            .O(N__27676),
            .I(N__27662));
    LocalMux I__5728 (
            .O(N__27673),
            .I(N__27657));
    InMux I__5727 (
            .O(N__27670),
            .I(N__27652));
    Span4Mux_v I__5726 (
            .O(N__27667),
            .I(N__27647));
    LocalMux I__5725 (
            .O(N__27662),
            .I(N__27647));
    InMux I__5724 (
            .O(N__27661),
            .I(N__27642));
    InMux I__5723 (
            .O(N__27660),
            .I(N__27642));
    Span4Mux_s1_h I__5722 (
            .O(N__27657),
            .I(N__27639));
    InMux I__5721 (
            .O(N__27656),
            .I(N__27634));
    InMux I__5720 (
            .O(N__27655),
            .I(N__27634));
    LocalMux I__5719 (
            .O(N__27652),
            .I(N__27629));
    Span4Mux_h I__5718 (
            .O(N__27647),
            .I(N__27629));
    LocalMux I__5717 (
            .O(N__27642),
            .I(N__27626));
    Odrv4 I__5716 (
            .O(N__27639),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    LocalMux I__5715 (
            .O(N__27634),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    Odrv4 I__5714 (
            .O(N__27629),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    Odrv12 I__5713 (
            .O(N__27626),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    CascadeMux I__5712 (
            .O(N__27617),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1_cascade_ ));
    CascadeMux I__5711 (
            .O(N__27614),
            .I(\POWERLED.func_state_RNI_8Z0Z_1_cascade_ ));
    InMux I__5710 (
            .O(N__27611),
            .I(N__27608));
    LocalMux I__5709 (
            .O(N__27608),
            .I(N__27605));
    Odrv4 I__5708 (
            .O(N__27605),
            .I(\POWERLED.func_state_RNIMQ0F_0Z0Z_1 ));
    InMux I__5707 (
            .O(N__27602),
            .I(N__27599));
    LocalMux I__5706 (
            .O(N__27599),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d ));
    CascadeMux I__5705 (
            .O(N__27596),
            .I(\POWERLED.func_state_RNIMQ0F_0Z0Z_1_cascade_ ));
    InMux I__5704 (
            .O(N__27593),
            .I(N__27590));
    LocalMux I__5703 (
            .O(N__27590),
            .I(\POWERLED.dutycycle_RNI2MQDZ0Z_7 ));
    CascadeMux I__5702 (
            .O(N__27587),
            .I(N__27584));
    InMux I__5701 (
            .O(N__27584),
            .I(N__27581));
    LocalMux I__5700 (
            .O(N__27581),
            .I(N__27578));
    Odrv12 I__5699 (
            .O(N__27578),
            .I(\POWERLED.dutycycle_RNIEBSB1Z0Z_7 ));
    InMux I__5698 (
            .O(N__27575),
            .I(N__27572));
    LocalMux I__5697 (
            .O(N__27572),
            .I(N__27569));
    Span12Mux_s3_h I__5696 (
            .O(N__27569),
            .I(N__27566));
    Odrv12 I__5695 (
            .O(N__27566),
            .I(\POWERLED.N_545 ));
    InMux I__5694 (
            .O(N__27563),
            .I(N__27560));
    LocalMux I__5693 (
            .O(N__27560),
            .I(N__27557));
    Span4Mux_s2_h I__5692 (
            .O(N__27557),
            .I(N__27554));
    Odrv4 I__5691 (
            .O(N__27554),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ));
    InMux I__5690 (
            .O(N__27551),
            .I(N__27545));
    InMux I__5689 (
            .O(N__27550),
            .I(N__27545));
    LocalMux I__5688 (
            .O(N__27545),
            .I(N__27542));
    Span4Mux_h I__5687 (
            .O(N__27542),
            .I(N__27539));
    Span4Mux_v I__5686 (
            .O(N__27539),
            .I(N__27536));
    Odrv4 I__5685 (
            .O(N__27536),
            .I(\POWERLED.N_71 ));
    InMux I__5684 (
            .O(N__27533),
            .I(N__27527));
    InMux I__5683 (
            .O(N__27532),
            .I(N__27527));
    LocalMux I__5682 (
            .O(N__27527),
            .I(N__27524));
    Span4Mux_s2_h I__5681 (
            .O(N__27524),
            .I(N__27521));
    Odrv4 I__5680 (
            .O(N__27521),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_a2_d ));
    InMux I__5679 (
            .O(N__27518),
            .I(N__27515));
    LocalMux I__5678 (
            .O(N__27515),
            .I(N__27512));
    Odrv12 I__5677 (
            .O(N__27512),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    InMux I__5676 (
            .O(N__27509),
            .I(N__27506));
    LocalMux I__5675 (
            .O(N__27506),
            .I(\POWERLED.dutycycle_e_1_4 ));
    CascadeMux I__5674 (
            .O(N__27503),
            .I(\POWERLED.dutycycle_e_1_4_cascade_ ));
    InMux I__5673 (
            .O(N__27500),
            .I(N__27494));
    InMux I__5672 (
            .O(N__27499),
            .I(N__27494));
    LocalMux I__5671 (
            .O(N__27494),
            .I(\POWERLED.func_state_RNIJ17U4Z0Z_1 ));
    InMux I__5670 (
            .O(N__27491),
            .I(N__27487));
    InMux I__5669 (
            .O(N__27490),
            .I(N__27484));
    LocalMux I__5668 (
            .O(N__27487),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    LocalMux I__5667 (
            .O(N__27484),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    InMux I__5666 (
            .O(N__27479),
            .I(N__27476));
    LocalMux I__5665 (
            .O(N__27476),
            .I(N__27473));
    Odrv4 I__5664 (
            .O(N__27473),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    InMux I__5663 (
            .O(N__27470),
            .I(N__27467));
    LocalMux I__5662 (
            .O(N__27467),
            .I(\POWERLED.dutycycle_e_1_7 ));
    InMux I__5661 (
            .O(N__27464),
            .I(N__27460));
    InMux I__5660 (
            .O(N__27463),
            .I(N__27457));
    LocalMux I__5659 (
            .O(N__27460),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    LocalMux I__5658 (
            .O(N__27457),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    CascadeMux I__5657 (
            .O(N__27452),
            .I(\POWERLED.dutycycle_e_1_7_cascade_ ));
    InMux I__5656 (
            .O(N__27449),
            .I(N__27443));
    InMux I__5655 (
            .O(N__27448),
            .I(N__27443));
    LocalMux I__5654 (
            .O(N__27443),
            .I(\POWERLED.func_state_RNI9S7D5Z0Z_1 ));
    CascadeMux I__5653 (
            .O(N__27440),
            .I(\POWERLED.dutycycleZ1Z_6_cascade_ ));
    InMux I__5652 (
            .O(N__27437),
            .I(N__27433));
    InMux I__5651 (
            .O(N__27436),
            .I(N__27430));
    LocalMux I__5650 (
            .O(N__27433),
            .I(N__27425));
    LocalMux I__5649 (
            .O(N__27430),
            .I(N__27425));
    Odrv4 I__5648 (
            .O(N__27425),
            .I(\POWERLED.N_133 ));
    CascadeMux I__5647 (
            .O(N__27422),
            .I(N__27417));
    CascadeMux I__5646 (
            .O(N__27421),
            .I(N__27412));
    InMux I__5645 (
            .O(N__27420),
            .I(N__27409));
    InMux I__5644 (
            .O(N__27417),
            .I(N__27406));
    InMux I__5643 (
            .O(N__27416),
            .I(N__27403));
    InMux I__5642 (
            .O(N__27415),
            .I(N__27400));
    InMux I__5641 (
            .O(N__27412),
            .I(N__27397));
    LocalMux I__5640 (
            .O(N__27409),
            .I(N__27393));
    LocalMux I__5639 (
            .O(N__27406),
            .I(N__27390));
    LocalMux I__5638 (
            .O(N__27403),
            .I(N__27386));
    LocalMux I__5637 (
            .O(N__27400),
            .I(N__27381));
    LocalMux I__5636 (
            .O(N__27397),
            .I(N__27381));
    InMux I__5635 (
            .O(N__27396),
            .I(N__27378));
    Span4Mux_v I__5634 (
            .O(N__27393),
            .I(N__27373));
    Span4Mux_v I__5633 (
            .O(N__27390),
            .I(N__27373));
    InMux I__5632 (
            .O(N__27389),
            .I(N__27370));
    Span4Mux_s2_h I__5631 (
            .O(N__27386),
            .I(N__27365));
    Span4Mux_h I__5630 (
            .O(N__27381),
            .I(N__27365));
    LocalMux I__5629 (
            .O(N__27378),
            .I(N__27362));
    Odrv4 I__5628 (
            .O(N__27373),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__5627 (
            .O(N__27370),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__5626 (
            .O(N__27365),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__5625 (
            .O(N__27362),
            .I(\POWERLED.func_stateZ0Z_0 ));
    CascadeMux I__5624 (
            .O(N__27353),
            .I(N__27349));
    InMux I__5623 (
            .O(N__27352),
            .I(N__27342));
    InMux I__5622 (
            .O(N__27349),
            .I(N__27342));
    InMux I__5621 (
            .O(N__27348),
            .I(N__27333));
    InMux I__5620 (
            .O(N__27347),
            .I(N__27333));
    LocalMux I__5619 (
            .O(N__27342),
            .I(N__27329));
    InMux I__5618 (
            .O(N__27341),
            .I(N__27326));
    InMux I__5617 (
            .O(N__27340),
            .I(N__27321));
    InMux I__5616 (
            .O(N__27339),
            .I(N__27321));
    InMux I__5615 (
            .O(N__27338),
            .I(N__27318));
    LocalMux I__5614 (
            .O(N__27333),
            .I(N__27313));
    InMux I__5613 (
            .O(N__27332),
            .I(N__27310));
    Span4Mux_v I__5612 (
            .O(N__27329),
            .I(N__27307));
    LocalMux I__5611 (
            .O(N__27326),
            .I(N__27300));
    LocalMux I__5610 (
            .O(N__27321),
            .I(N__27300));
    LocalMux I__5609 (
            .O(N__27318),
            .I(N__27300));
    InMux I__5608 (
            .O(N__27317),
            .I(N__27297));
    InMux I__5607 (
            .O(N__27316),
            .I(N__27294));
    Span4Mux_s3_h I__5606 (
            .O(N__27313),
            .I(N__27289));
    LocalMux I__5605 (
            .O(N__27310),
            .I(N__27289));
    Span4Mux_v I__5604 (
            .O(N__27307),
            .I(N__27284));
    Span4Mux_v I__5603 (
            .O(N__27300),
            .I(N__27284));
    LocalMux I__5602 (
            .O(N__27297),
            .I(\POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0 ));
    LocalMux I__5601 (
            .O(N__27294),
            .I(\POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0 ));
    Odrv4 I__5600 (
            .O(N__27289),
            .I(\POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0 ));
    Odrv4 I__5599 (
            .O(N__27284),
            .I(\POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0 ));
    InMux I__5598 (
            .O(N__27275),
            .I(N__27272));
    LocalMux I__5597 (
            .O(N__27272),
            .I(\POWERLED.N_490 ));
    InMux I__5596 (
            .O(N__27269),
            .I(N__27266));
    LocalMux I__5595 (
            .O(N__27266),
            .I(N__27263));
    Span4Mux_v I__5594 (
            .O(N__27263),
            .I(N__27260));
    Odrv4 I__5593 (
            .O(N__27260),
            .I(\POWERLED.g1_0_2 ));
    CascadeMux I__5592 (
            .O(N__27257),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_0_cascade_ ));
    InMux I__5591 (
            .O(N__27254),
            .I(N__27251));
    LocalMux I__5590 (
            .O(N__27251),
            .I(N__27248));
    Span4Mux_v I__5589 (
            .O(N__27248),
            .I(N__27245));
    Odrv4 I__5588 (
            .O(N__27245),
            .I(\POWERLED.dutycycle_eena_13_1_0 ));
    InMux I__5587 (
            .O(N__27242),
            .I(N__27239));
    LocalMux I__5586 (
            .O(N__27239),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6 ));
    CascadeMux I__5585 (
            .O(N__27236),
            .I(N__27232));
    InMux I__5584 (
            .O(N__27235),
            .I(N__27229));
    InMux I__5583 (
            .O(N__27232),
            .I(N__27226));
    LocalMux I__5582 (
            .O(N__27229),
            .I(N__27223));
    LocalMux I__5581 (
            .O(N__27226),
            .I(N__27220));
    Span4Mux_s1_h I__5580 (
            .O(N__27223),
            .I(N__27215));
    Span4Mux_v I__5579 (
            .O(N__27220),
            .I(N__27215));
    Span4Mux_h I__5578 (
            .O(N__27215),
            .I(N__27212));
    Span4Mux_v I__5577 (
            .O(N__27212),
            .I(N__27209));
    Odrv4 I__5576 (
            .O(N__27209),
            .I(\POWERLED.count_offZ0Z_7 ));
    CascadeMux I__5575 (
            .O(N__27206),
            .I(\POWERLED.count_offZ0Z_3_cascade_ ));
    CascadeMux I__5574 (
            .O(N__27203),
            .I(N__27199));
    InMux I__5573 (
            .O(N__27202),
            .I(N__27196));
    InMux I__5572 (
            .O(N__27199),
            .I(N__27193));
    LocalMux I__5571 (
            .O(N__27196),
            .I(N__27190));
    LocalMux I__5570 (
            .O(N__27193),
            .I(N__27187));
    Span12Mux_s5_h I__5569 (
            .O(N__27190),
            .I(N__27184));
    Span12Mux_v I__5568 (
            .O(N__27187),
            .I(N__27181));
    Odrv12 I__5567 (
            .O(N__27184),
            .I(\POWERLED.count_offZ0Z_8 ));
    Odrv12 I__5566 (
            .O(N__27181),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__5565 (
            .O(N__27176),
            .I(N__27173));
    LocalMux I__5564 (
            .O(N__27173),
            .I(N__27170));
    Span4Mux_v I__5563 (
            .O(N__27170),
            .I(N__27167));
    Odrv4 I__5562 (
            .O(N__27167),
            .I(\POWERLED.un34_clk_100khz_11 ));
    CascadeMux I__5561 (
            .O(N__27164),
            .I(\POWERLED.un34_clk_100khz_8_cascade_ ));
    CascadeMux I__5560 (
            .O(N__27161),
            .I(\POWERLED.count_off_RNI_0Z0Z_10_cascade_ ));
    CascadeMux I__5559 (
            .O(N__27158),
            .I(\POWERLED.count_off_RNI8AQHZ0Z_10_cascade_ ));
    InMux I__5558 (
            .O(N__27155),
            .I(N__27152));
    LocalMux I__5557 (
            .O(N__27152),
            .I(\POWERLED.func_state_1_m2_ns_1_1 ));
    InMux I__5556 (
            .O(N__27149),
            .I(N__27146));
    LocalMux I__5555 (
            .O(N__27146),
            .I(N__27143));
    Span4Mux_v I__5554 (
            .O(N__27143),
            .I(N__27140));
    Span4Mux_v I__5553 (
            .O(N__27140),
            .I(N__27137));
    Odrv4 I__5552 (
            .O(N__27137),
            .I(\POWERLED.N_494 ));
    CascadeMux I__5551 (
            .O(N__27134),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_ ));
    InMux I__5550 (
            .O(N__27131),
            .I(N__27128));
    LocalMux I__5549 (
            .O(N__27128),
            .I(N__27125));
    Span4Mux_s2_h I__5548 (
            .O(N__27125),
            .I(N__27122));
    Odrv4 I__5547 (
            .O(N__27122),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ));
    CascadeMux I__5546 (
            .O(N__27119),
            .I(\POWERLED.dutycycle_1_0_iv_i_i_m2_1_6_cascade_ ));
    InMux I__5545 (
            .O(N__27116),
            .I(N__27113));
    LocalMux I__5544 (
            .O(N__27113),
            .I(N__27110));
    Span4Mux_v I__5543 (
            .O(N__27110),
            .I(N__27107));
    Span4Mux_h I__5542 (
            .O(N__27107),
            .I(N__27104));
    Odrv4 I__5541 (
            .O(N__27104),
            .I(\POWERLED.N_453 ));
    InMux I__5540 (
            .O(N__27101),
            .I(N__27098));
    LocalMux I__5539 (
            .O(N__27098),
            .I(N__27095));
    Odrv4 I__5538 (
            .O(N__27095),
            .I(\POWERLED.N_426_i ));
    InMux I__5537 (
            .O(N__27092),
            .I(N__27089));
    LocalMux I__5536 (
            .O(N__27089),
            .I(\POWERLED.N_562 ));
    CascadeMux I__5535 (
            .O(N__27086),
            .I(N__27083));
    InMux I__5534 (
            .O(N__27083),
            .I(N__27079));
    InMux I__5533 (
            .O(N__27082),
            .I(N__27076));
    LocalMux I__5532 (
            .O(N__27079),
            .I(N__27071));
    LocalMux I__5531 (
            .O(N__27076),
            .I(N__27071));
    Odrv12 I__5530 (
            .O(N__27071),
            .I(\POWERLED.func_state_enZ0 ));
    InMux I__5529 (
            .O(N__27068),
            .I(N__27065));
    LocalMux I__5528 (
            .O(N__27065),
            .I(\POWERLED.func_state_1_m2_1 ));
    InMux I__5527 (
            .O(N__27062),
            .I(N__27056));
    InMux I__5526 (
            .O(N__27061),
            .I(N__27056));
    LocalMux I__5525 (
            .O(N__27056),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__5524 (
            .O(N__27053),
            .I(N__27050));
    LocalMux I__5523 (
            .O(N__27050),
            .I(\POWERLED.count_off_0_4 ));
    CascadeMux I__5522 (
            .O(N__27047),
            .I(N__27044));
    InMux I__5521 (
            .O(N__27044),
            .I(N__27038));
    InMux I__5520 (
            .O(N__27043),
            .I(N__27038));
    LocalMux I__5519 (
            .O(N__27038),
            .I(N__27035));
    Odrv4 I__5518 (
            .O(N__27035),
            .I(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ));
    InMux I__5517 (
            .O(N__27032),
            .I(N__27029));
    LocalMux I__5516 (
            .O(N__27029),
            .I(\POWERLED.count_off_0_3 ));
    InMux I__5515 (
            .O(N__27026),
            .I(N__27020));
    InMux I__5514 (
            .O(N__27025),
            .I(N__27020));
    LocalMux I__5513 (
            .O(N__27020),
            .I(N__27017));
    Odrv4 I__5512 (
            .O(N__27017),
            .I(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ));
    InMux I__5511 (
            .O(N__27014),
            .I(N__27011));
    LocalMux I__5510 (
            .O(N__27011),
            .I(N__27008));
    Odrv4 I__5509 (
            .O(N__27008),
            .I(\POWERLED.count_offZ0Z_3 ));
    CascadeMux I__5508 (
            .O(N__27005),
            .I(N__27002));
    InMux I__5507 (
            .O(N__27002),
            .I(N__26998));
    InMux I__5506 (
            .O(N__27001),
            .I(N__26995));
    LocalMux I__5505 (
            .O(N__26998),
            .I(N__26992));
    LocalMux I__5504 (
            .O(N__26995),
            .I(\POWERLED.count_offZ0Z_4 ));
    Odrv4 I__5503 (
            .O(N__26992),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__5502 (
            .O(N__26987),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    CascadeMux I__5501 (
            .O(N__26984),
            .I(N__26981));
    InMux I__5500 (
            .O(N__26981),
            .I(N__26977));
    InMux I__5499 (
            .O(N__26980),
            .I(N__26974));
    LocalMux I__5498 (
            .O(N__26977),
            .I(N__26971));
    LocalMux I__5497 (
            .O(N__26974),
            .I(\POWERLED.count_offZ0Z_12 ));
    Odrv4 I__5496 (
            .O(N__26971),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__5495 (
            .O(N__26966),
            .I(N__26960));
    InMux I__5494 (
            .O(N__26965),
            .I(N__26960));
    LocalMux I__5493 (
            .O(N__26960),
            .I(N__26957));
    Odrv4 I__5492 (
            .O(N__26957),
            .I(\POWERLED.count_off_1_12 ));
    InMux I__5491 (
            .O(N__26954),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__5490 (
            .O(N__26951),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__5489 (
            .O(N__26948),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__5488 (
            .O(N__26945),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__5487 (
            .O(N__26942),
            .I(N__26939));
    LocalMux I__5486 (
            .O(N__26939),
            .I(N__26936));
    Span4Mux_v I__5485 (
            .O(N__26936),
            .I(N__26933));
    Odrv4 I__5484 (
            .O(N__26933),
            .I(\POWERLED.N_627 ));
    CascadeMux I__5483 (
            .O(N__26930),
            .I(N__26927));
    InMux I__5482 (
            .O(N__26927),
            .I(N__26924));
    LocalMux I__5481 (
            .O(N__26924),
            .I(N__26921));
    Odrv12 I__5480 (
            .O(N__26921),
            .I(\POWERLED.N_688 ));
    InMux I__5479 (
            .O(N__26918),
            .I(N__26914));
    InMux I__5478 (
            .O(N__26917),
            .I(N__26911));
    LocalMux I__5477 (
            .O(N__26914),
            .I(N__26908));
    LocalMux I__5476 (
            .O(N__26911),
            .I(N__26904));
    Span4Mux_h I__5475 (
            .O(N__26908),
            .I(N__26901));
    CascadeMux I__5474 (
            .O(N__26907),
            .I(N__26898));
    Span4Mux_s3_h I__5473 (
            .O(N__26904),
            .I(N__26893));
    Span4Mux_v I__5472 (
            .O(N__26901),
            .I(N__26893));
    InMux I__5471 (
            .O(N__26898),
            .I(N__26890));
    Odrv4 I__5470 (
            .O(N__26893),
            .I(\POWERLED.N_74 ));
    LocalMux I__5469 (
            .O(N__26890),
            .I(\POWERLED.N_74 ));
    CascadeMux I__5468 (
            .O(N__26885),
            .I(\POWERLED.N_6_1_cascade_ ));
    CascadeMux I__5467 (
            .O(N__26882),
            .I(\POWERLED.func_state_1_m2_1_cascade_ ));
    CascadeMux I__5466 (
            .O(N__26879),
            .I(\POWERLED.func_state_cascade_ ));
    InMux I__5465 (
            .O(N__26876),
            .I(\POWERLED.un3_count_off_1_cry_1 ));
    InMux I__5464 (
            .O(N__26873),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    InMux I__5463 (
            .O(N__26870),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    InMux I__5462 (
            .O(N__26867),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    InMux I__5461 (
            .O(N__26864),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    InMux I__5460 (
            .O(N__26861),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__5459 (
            .O(N__26858),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__5458 (
            .O(N__26855),
            .I(N__26852));
    LocalMux I__5457 (
            .O(N__26852),
            .I(N__26849));
    Odrv4 I__5456 (
            .O(N__26849),
            .I(\POWERLED.count_offZ0Z_9 ));
    InMux I__5455 (
            .O(N__26846),
            .I(N__26840));
    InMux I__5454 (
            .O(N__26845),
            .I(N__26840));
    LocalMux I__5453 (
            .O(N__26840),
            .I(N__26837));
    Odrv4 I__5452 (
            .O(N__26837),
            .I(\POWERLED.count_off_1_9 ));
    InMux I__5451 (
            .O(N__26834),
            .I(bfn_11_4_0_));
    CascadeMux I__5450 (
            .O(N__26831),
            .I(N__26828));
    InMux I__5449 (
            .O(N__26828),
            .I(N__26824));
    InMux I__5448 (
            .O(N__26827),
            .I(N__26821));
    LocalMux I__5447 (
            .O(N__26824),
            .I(N__26818));
    LocalMux I__5446 (
            .O(N__26821),
            .I(\POWERLED.count_offZ0Z_10 ));
    Odrv4 I__5445 (
            .O(N__26818),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__5444 (
            .O(N__26813),
            .I(N__26807));
    InMux I__5443 (
            .O(N__26812),
            .I(N__26807));
    LocalMux I__5442 (
            .O(N__26807),
            .I(N__26804));
    Odrv4 I__5441 (
            .O(N__26804),
            .I(\POWERLED.count_off_1_10 ));
    InMux I__5440 (
            .O(N__26801),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    InMux I__5439 (
            .O(N__26798),
            .I(N__26794));
    InMux I__5438 (
            .O(N__26797),
            .I(N__26791));
    LocalMux I__5437 (
            .O(N__26794),
            .I(\POWERLED.count_clkZ0Z_14 ));
    LocalMux I__5436 (
            .O(N__26791),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__5435 (
            .O(N__26786),
            .I(N__26783));
    LocalMux I__5434 (
            .O(N__26783),
            .I(\POWERLED.count_off_0_9 ));
    CascadeMux I__5433 (
            .O(N__26780),
            .I(\POWERLED.count_offZ0Z_9_cascade_ ));
    InMux I__5432 (
            .O(N__26777),
            .I(N__26774));
    LocalMux I__5431 (
            .O(N__26774),
            .I(\POWERLED.count_off_0_10 ));
    InMux I__5430 (
            .O(N__26771),
            .I(N__26768));
    LocalMux I__5429 (
            .O(N__26768),
            .I(\POWERLED.count_off_0_12 ));
    InMux I__5428 (
            .O(N__26765),
            .I(N__26758));
    InMux I__5427 (
            .O(N__26764),
            .I(N__26758));
    InMux I__5426 (
            .O(N__26763),
            .I(N__26755));
    LocalMux I__5425 (
            .O(N__26758),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__5424 (
            .O(N__26755),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__5423 (
            .O(N__26750),
            .I(N__26746));
    InMux I__5422 (
            .O(N__26749),
            .I(N__26743));
    LocalMux I__5421 (
            .O(N__26746),
            .I(\POWERLED.count_clkZ0Z_9 ));
    LocalMux I__5420 (
            .O(N__26743),
            .I(\POWERLED.count_clkZ0Z_9 ));
    CascadeMux I__5419 (
            .O(N__26738),
            .I(\POWERLED.count_clkZ0Z_7_cascade_ ));
    InMux I__5418 (
            .O(N__26735),
            .I(N__26732));
    LocalMux I__5417 (
            .O(N__26732),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3 ));
    InMux I__5416 (
            .O(N__26729),
            .I(N__26723));
    InMux I__5415 (
            .O(N__26728),
            .I(N__26723));
    LocalMux I__5414 (
            .O(N__26723),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    InMux I__5413 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__5412 (
            .O(N__26717),
            .I(\POWERLED.count_clk_0_7 ));
    InMux I__5411 (
            .O(N__26714),
            .I(N__26711));
    LocalMux I__5410 (
            .O(N__26711),
            .I(N__26707));
    InMux I__5409 (
            .O(N__26710),
            .I(N__26704));
    Span4Mux_h I__5408 (
            .O(N__26707),
            .I(N__26699));
    LocalMux I__5407 (
            .O(N__26704),
            .I(N__26699));
    Odrv4 I__5406 (
            .O(N__26699),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__5405 (
            .O(N__26696),
            .I(N__26693));
    LocalMux I__5404 (
            .O(N__26693),
            .I(N__26688));
    InMux I__5403 (
            .O(N__26692),
            .I(N__26685));
    InMux I__5402 (
            .O(N__26691),
            .I(N__26682));
    Span4Mux_h I__5401 (
            .O(N__26688),
            .I(N__26679));
    LocalMux I__5400 (
            .O(N__26685),
            .I(\POWERLED.count_clk_1_10 ));
    LocalMux I__5399 (
            .O(N__26682),
            .I(\POWERLED.count_clk_1_10 ));
    Odrv4 I__5398 (
            .O(N__26679),
            .I(\POWERLED.count_clk_1_10 ));
    InMux I__5397 (
            .O(N__26672),
            .I(N__26669));
    LocalMux I__5396 (
            .O(N__26669),
            .I(N__26665));
    InMux I__5395 (
            .O(N__26668),
            .I(N__26662));
    Span4Mux_s2_v I__5394 (
            .O(N__26665),
            .I(N__26659));
    LocalMux I__5393 (
            .O(N__26662),
            .I(N__26656));
    Odrv4 I__5392 (
            .O(N__26659),
            .I(\POWERLED.count_clkZ0Z_15 ));
    Odrv4 I__5391 (
            .O(N__26656),
            .I(\POWERLED.count_clkZ0Z_15 ));
    CascadeMux I__5390 (
            .O(N__26651),
            .I(N__26647));
    InMux I__5389 (
            .O(N__26650),
            .I(N__26644));
    InMux I__5388 (
            .O(N__26647),
            .I(N__26641));
    LocalMux I__5387 (
            .O(N__26644),
            .I(N__26638));
    LocalMux I__5386 (
            .O(N__26641),
            .I(N__26635));
    Odrv4 I__5385 (
            .O(N__26638),
            .I(\POWERLED.count_clkZ0Z_10 ));
    Odrv4 I__5384 (
            .O(N__26635),
            .I(\POWERLED.count_clkZ0Z_10 ));
    InMux I__5383 (
            .O(N__26630),
            .I(N__26627));
    LocalMux I__5382 (
            .O(N__26627),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_0 ));
    CascadeMux I__5381 (
            .O(N__26624),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_2_cascade_ ));
    InMux I__5380 (
            .O(N__26621),
            .I(N__26618));
    LocalMux I__5379 (
            .O(N__26618),
            .I(N__26614));
    InMux I__5378 (
            .O(N__26617),
            .I(N__26611));
    Odrv4 I__5377 (
            .O(N__26614),
            .I(\POWERLED.count_clk_RNINSEUCZ0Z_10 ));
    LocalMux I__5376 (
            .O(N__26611),
            .I(\POWERLED.count_clk_RNINSEUCZ0Z_10 ));
    InMux I__5375 (
            .O(N__26606),
            .I(N__26603));
    LocalMux I__5374 (
            .O(N__26603),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_1 ));
    InMux I__5373 (
            .O(N__26600),
            .I(N__26594));
    InMux I__5372 (
            .O(N__26599),
            .I(N__26594));
    LocalMux I__5371 (
            .O(N__26594),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__5370 (
            .O(N__26591),
            .I(N__26582));
    InMux I__5369 (
            .O(N__26590),
            .I(N__26582));
    InMux I__5368 (
            .O(N__26589),
            .I(N__26582));
    LocalMux I__5367 (
            .O(N__26582),
            .I(\POWERLED.count_clk_1_12 ));
    InMux I__5366 (
            .O(N__26579),
            .I(N__26576));
    LocalMux I__5365 (
            .O(N__26576),
            .I(\POWERLED.un1_count_clk_2_axb_12 ));
    InMux I__5364 (
            .O(N__26573),
            .I(N__26566));
    InMux I__5363 (
            .O(N__26572),
            .I(N__26566));
    InMux I__5362 (
            .O(N__26571),
            .I(N__26563));
    LocalMux I__5361 (
            .O(N__26566),
            .I(\POWERLED.count_clk_1_14 ));
    LocalMux I__5360 (
            .O(N__26563),
            .I(\POWERLED.count_clk_1_14 ));
    InMux I__5359 (
            .O(N__26558),
            .I(N__26552));
    InMux I__5358 (
            .O(N__26557),
            .I(N__26552));
    LocalMux I__5357 (
            .O(N__26552),
            .I(\POWERLED.count_clk_0_3 ));
    InMux I__5356 (
            .O(N__26549),
            .I(N__26543));
    InMux I__5355 (
            .O(N__26548),
            .I(N__26543));
    LocalMux I__5354 (
            .O(N__26543),
            .I(N__26539));
    InMux I__5353 (
            .O(N__26542),
            .I(N__26536));
    Odrv4 I__5352 (
            .O(N__26539),
            .I(\POWERLED.count_clkZ0Z_8 ));
    LocalMux I__5351 (
            .O(N__26536),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__5350 (
            .O(N__26531),
            .I(N__26524));
    InMux I__5349 (
            .O(N__26530),
            .I(N__26524));
    InMux I__5348 (
            .O(N__26529),
            .I(N__26521));
    LocalMux I__5347 (
            .O(N__26524),
            .I(N__26518));
    LocalMux I__5346 (
            .O(N__26521),
            .I(N__26515));
    Span4Mux_s3_h I__5345 (
            .O(N__26518),
            .I(N__26510));
    Span4Mux_s2_v I__5344 (
            .O(N__26515),
            .I(N__26510));
    Odrv4 I__5343 (
            .O(N__26510),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__5342 (
            .O(N__26507),
            .I(N__26502));
    InMux I__5341 (
            .O(N__26506),
            .I(N__26499));
    InMux I__5340 (
            .O(N__26505),
            .I(N__26496));
    LocalMux I__5339 (
            .O(N__26502),
            .I(N__26493));
    LocalMux I__5338 (
            .O(N__26499),
            .I(N__26488));
    LocalMux I__5337 (
            .O(N__26496),
            .I(N__26488));
    Span4Mux_s2_v I__5336 (
            .O(N__26493),
            .I(N__26485));
    Odrv4 I__5335 (
            .O(N__26488),
            .I(\POWERLED.count_clkZ0Z_4 ));
    Odrv4 I__5334 (
            .O(N__26485),
            .I(\POWERLED.count_clkZ0Z_4 ));
    CascadeMux I__5333 (
            .O(N__26480),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_ ));
    InMux I__5332 (
            .O(N__26477),
            .I(N__26472));
    InMux I__5331 (
            .O(N__26476),
            .I(N__26467));
    InMux I__5330 (
            .O(N__26475),
            .I(N__26467));
    LocalMux I__5329 (
            .O(N__26472),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__5328 (
            .O(N__26467),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__5327 (
            .O(N__26462),
            .I(N__26459));
    LocalMux I__5326 (
            .O(N__26459),
            .I(\POWERLED.N_625 ));
    CascadeMux I__5325 (
            .O(N__26456),
            .I(\POWERLED.N_625_cascade_ ));
    CascadeMux I__5324 (
            .O(N__26453),
            .I(\POWERLED.count_clkZ0Z_9_cascade_ ));
    InMux I__5323 (
            .O(N__26450),
            .I(N__26444));
    InMux I__5322 (
            .O(N__26449),
            .I(N__26444));
    LocalMux I__5321 (
            .O(N__26444),
            .I(\POWERLED.count_clk_RNINSEUC_0Z0Z_10 ));
    InMux I__5320 (
            .O(N__26441),
            .I(N__26435));
    InMux I__5319 (
            .O(N__26440),
            .I(N__26435));
    LocalMux I__5318 (
            .O(N__26435),
            .I(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ));
    InMux I__5317 (
            .O(N__26432),
            .I(N__26429));
    LocalMux I__5316 (
            .O(N__26429),
            .I(\POWERLED.count_clk_0_9 ));
    InMux I__5315 (
            .O(N__26426),
            .I(N__26423));
    LocalMux I__5314 (
            .O(N__26423),
            .I(N__26420));
    Odrv4 I__5313 (
            .O(N__26420),
            .I(\POWERLED.count_clk_0_5 ));
    InMux I__5312 (
            .O(N__26417),
            .I(N__26411));
    InMux I__5311 (
            .O(N__26416),
            .I(N__26411));
    LocalMux I__5310 (
            .O(N__26411),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    InMux I__5309 (
            .O(N__26408),
            .I(N__26401));
    InMux I__5308 (
            .O(N__26407),
            .I(N__26401));
    InMux I__5307 (
            .O(N__26406),
            .I(N__26398));
    LocalMux I__5306 (
            .O(N__26401),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__5305 (
            .O(N__26398),
            .I(\POWERLED.count_clkZ0Z_7 ));
    InMux I__5304 (
            .O(N__26393),
            .I(N__26387));
    InMux I__5303 (
            .O(N__26392),
            .I(N__26387));
    LocalMux I__5302 (
            .O(N__26387),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__5301 (
            .O(N__26384),
            .I(N__26380));
    InMux I__5300 (
            .O(N__26383),
            .I(N__26375));
    InMux I__5299 (
            .O(N__26380),
            .I(N__26375));
    LocalMux I__5298 (
            .O(N__26375),
            .I(N__26372));
    Odrv12 I__5297 (
            .O(N__26372),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ));
    InMux I__5296 (
            .O(N__26369),
            .I(N__26366));
    LocalMux I__5295 (
            .O(N__26366),
            .I(\POWERLED.dutycycle_RNIHDMC5Z0Z_9 ));
    CascadeMux I__5294 (
            .O(N__26363),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    CascadeMux I__5293 (
            .O(N__26360),
            .I(\POWERLED.N_17_cascade_ ));
    InMux I__5292 (
            .O(N__26357),
            .I(N__26354));
    LocalMux I__5291 (
            .O(N__26354),
            .I(N__26351));
    Odrv4 I__5290 (
            .O(N__26351),
            .I(\POWERLED.N_8_2 ));
    InMux I__5289 (
            .O(N__26348),
            .I(N__26345));
    LocalMux I__5288 (
            .O(N__26345),
            .I(\POWERLED.G_7_i_0 ));
    InMux I__5287 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__5286 (
            .O(N__26339),
            .I(\POWERLED.count_clkZ0Z_3 ));
    CascadeMux I__5285 (
            .O(N__26336),
            .I(\POWERLED.count_clkZ0Z_3_cascade_ ));
    CascadeMux I__5284 (
            .O(N__26333),
            .I(\POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_ ));
    InMux I__5283 (
            .O(N__26330),
            .I(N__26321));
    InMux I__5282 (
            .O(N__26329),
            .I(N__26321));
    InMux I__5281 (
            .O(N__26328),
            .I(N__26321));
    LocalMux I__5280 (
            .O(N__26321),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    CascadeMux I__5279 (
            .O(N__26318),
            .I(\POWERLED.dutycycleZ0Z_2_cascade_ ));
    InMux I__5278 (
            .O(N__26315),
            .I(N__26312));
    LocalMux I__5277 (
            .O(N__26312),
            .I(\POWERLED.g0_9_1 ));
    InMux I__5276 (
            .O(N__26309),
            .I(N__26306));
    LocalMux I__5275 (
            .O(N__26306),
            .I(\POWERLED.g0_9_1_1_0 ));
    InMux I__5274 (
            .O(N__26303),
            .I(N__26299));
    CascadeMux I__5273 (
            .O(N__26302),
            .I(N__26296));
    LocalMux I__5272 (
            .O(N__26299),
            .I(N__26293));
    InMux I__5271 (
            .O(N__26296),
            .I(N__26290));
    Odrv4 I__5270 (
            .O(N__26293),
            .I(\POWERLED.dutycycle_RNIHDMC5Z0Z_10 ));
    LocalMux I__5269 (
            .O(N__26290),
            .I(\POWERLED.dutycycle_RNIHDMC5Z0Z_10 ));
    InMux I__5268 (
            .O(N__26285),
            .I(N__26279));
    InMux I__5267 (
            .O(N__26284),
            .I(N__26279));
    LocalMux I__5266 (
            .O(N__26279),
            .I(N__26276));
    Odrv4 I__5265 (
            .O(N__26276),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ));
    CascadeMux I__5264 (
            .O(N__26273),
            .I(N__26270));
    InMux I__5263 (
            .O(N__26270),
            .I(N__26264));
    InMux I__5262 (
            .O(N__26269),
            .I(N__26264));
    LocalMux I__5261 (
            .O(N__26264),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    InMux I__5260 (
            .O(N__26261),
            .I(N__26258));
    LocalMux I__5259 (
            .O(N__26258),
            .I(N__26255));
    Span4Mux_v I__5258 (
            .O(N__26255),
            .I(N__26252));
    Span4Mux_v I__5257 (
            .O(N__26252),
            .I(N__26249));
    Odrv4 I__5256 (
            .O(N__26249),
            .I(\POWERLED.dutycycle_RNI6SKJ1Z0Z_9 ));
    CascadeMux I__5255 (
            .O(N__26246),
            .I(\POWERLED.dutycycle_RNIHDMC5Z0Z_9_cascade_ ));
    InMux I__5254 (
            .O(N__26243),
            .I(N__26239));
    InMux I__5253 (
            .O(N__26242),
            .I(N__26234));
    LocalMux I__5252 (
            .O(N__26239),
            .I(N__26229));
    CascadeMux I__5251 (
            .O(N__26238),
            .I(N__26224));
    InMux I__5250 (
            .O(N__26237),
            .I(N__26221));
    LocalMux I__5249 (
            .O(N__26234),
            .I(N__26218));
    InMux I__5248 (
            .O(N__26233),
            .I(N__26213));
    InMux I__5247 (
            .O(N__26232),
            .I(N__26213));
    Span4Mux_v I__5246 (
            .O(N__26229),
            .I(N__26210));
    InMux I__5245 (
            .O(N__26228),
            .I(N__26207));
    InMux I__5244 (
            .O(N__26227),
            .I(N__26204));
    InMux I__5243 (
            .O(N__26224),
            .I(N__26201));
    LocalMux I__5242 (
            .O(N__26221),
            .I(N__26196));
    Span4Mux_h I__5241 (
            .O(N__26218),
            .I(N__26196));
    LocalMux I__5240 (
            .O(N__26213),
            .I(N__26193));
    Odrv4 I__5239 (
            .O(N__26210),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__5238 (
            .O(N__26207),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__5237 (
            .O(N__26204),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__5236 (
            .O(N__26201),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__5235 (
            .O(N__26196),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv12 I__5234 (
            .O(N__26193),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    InMux I__5233 (
            .O(N__26180),
            .I(N__26177));
    LocalMux I__5232 (
            .O(N__26177),
            .I(\POWERLED.un1_dutycycle_53_7_0 ));
    CascadeMux I__5231 (
            .O(N__26174),
            .I(\POWERLED.un1_dutycycle_53_41_0_cascade_ ));
    CascadeMux I__5230 (
            .O(N__26171),
            .I(N__26168));
    InMux I__5229 (
            .O(N__26168),
            .I(N__26165));
    LocalMux I__5228 (
            .O(N__26165),
            .I(N__26162));
    Span4Mux_h I__5227 (
            .O(N__26162),
            .I(N__26159));
    Odrv4 I__5226 (
            .O(N__26159),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_13 ));
    InMux I__5225 (
            .O(N__26156),
            .I(N__26153));
    LocalMux I__5224 (
            .O(N__26153),
            .I(\POWERLED.un1_dutycycle_53_59_a0_0 ));
    CascadeMux I__5223 (
            .O(N__26150),
            .I(N__26147));
    InMux I__5222 (
            .O(N__26147),
            .I(N__26141));
    InMux I__5221 (
            .O(N__26146),
            .I(N__26141));
    LocalMux I__5220 (
            .O(N__26141),
            .I(\POWERLED.dutycycleZ1Z_11 ));
    CascadeMux I__5219 (
            .O(N__26138),
            .I(N__26134));
    InMux I__5218 (
            .O(N__26137),
            .I(N__26129));
    InMux I__5217 (
            .O(N__26134),
            .I(N__26129));
    LocalMux I__5216 (
            .O(N__26129),
            .I(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ));
    CascadeMux I__5215 (
            .O(N__26126),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    CascadeMux I__5214 (
            .O(N__26123),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_12_cascade_ ));
    InMux I__5213 (
            .O(N__26120),
            .I(N__26116));
    InMux I__5212 (
            .O(N__26119),
            .I(N__26113));
    LocalMux I__5211 (
            .O(N__26116),
            .I(\POWERLED.un1_dutycycle_53_56_a1_2 ));
    LocalMux I__5210 (
            .O(N__26113),
            .I(\POWERLED.un1_dutycycle_53_56_a1_2 ));
    CascadeMux I__5209 (
            .O(N__26108),
            .I(N__26105));
    InMux I__5208 (
            .O(N__26105),
            .I(N__26102));
    LocalMux I__5207 (
            .O(N__26102),
            .I(N__26099));
    Span4Mux_h I__5206 (
            .O(N__26099),
            .I(N__26096));
    Odrv4 I__5205 (
            .O(N__26096),
            .I(\POWERLED.un1_dutycycle_53_8_2 ));
    InMux I__5204 (
            .O(N__26093),
            .I(N__26090));
    LocalMux I__5203 (
            .O(N__26090),
            .I(\POWERLED.un1_dutycycle_53_8_0 ));
    CascadeMux I__5202 (
            .O(N__26087),
            .I(N__26084));
    InMux I__5201 (
            .O(N__26084),
            .I(N__26081));
    LocalMux I__5200 (
            .O(N__26081),
            .I(N__26078));
    Odrv4 I__5199 (
            .O(N__26078),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    CascadeMux I__5198 (
            .O(N__26075),
            .I(\POWERLED.G_7_i_a5_1_1_cascade_ ));
    InMux I__5197 (
            .O(N__26072),
            .I(N__26069));
    LocalMux I__5196 (
            .O(N__26069),
            .I(\POWERLED.N_11_1 ));
    CascadeMux I__5195 (
            .O(N__26066),
            .I(\POWERLED.N_16_1_cascade_ ));
    InMux I__5194 (
            .O(N__26063),
            .I(N__26060));
    LocalMux I__5193 (
            .O(N__26060),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_9 ));
    InMux I__5192 (
            .O(N__26057),
            .I(\POWERLED.un1_dutycycle_94_cry_9 ));
    InMux I__5191 (
            .O(N__26054),
            .I(\POWERLED.un1_dutycycle_94_cry_10 ));
    CascadeMux I__5190 (
            .O(N__26051),
            .I(N__26047));
    InMux I__5189 (
            .O(N__26050),
            .I(N__26042));
    InMux I__5188 (
            .O(N__26047),
            .I(N__26042));
    LocalMux I__5187 (
            .O(N__26042),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ));
    InMux I__5186 (
            .O(N__26039),
            .I(\POWERLED.un1_dutycycle_94_cry_11 ));
    InMux I__5185 (
            .O(N__26036),
            .I(N__26030));
    InMux I__5184 (
            .O(N__26035),
            .I(N__26030));
    LocalMux I__5183 (
            .O(N__26030),
            .I(N__26027));
    Odrv4 I__5182 (
            .O(N__26027),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    InMux I__5181 (
            .O(N__26024),
            .I(\POWERLED.un1_dutycycle_94_cry_12_cZ0 ));
    InMux I__5180 (
            .O(N__26021),
            .I(N__26012));
    InMux I__5179 (
            .O(N__26020),
            .I(N__26012));
    InMux I__5178 (
            .O(N__26019),
            .I(N__26012));
    LocalMux I__5177 (
            .O(N__26012),
            .I(N__26002));
    InMux I__5176 (
            .O(N__26011),
            .I(N__25993));
    InMux I__5175 (
            .O(N__26010),
            .I(N__25993));
    InMux I__5174 (
            .O(N__26009),
            .I(N__25993));
    InMux I__5173 (
            .O(N__26008),
            .I(N__25993));
    CascadeMux I__5172 (
            .O(N__26007),
            .I(N__25990));
    CascadeMux I__5171 (
            .O(N__26006),
            .I(N__25984));
    CascadeMux I__5170 (
            .O(N__26005),
            .I(N__25980));
    Span4Mux_s3_h I__5169 (
            .O(N__26002),
            .I(N__25977));
    LocalMux I__5168 (
            .O(N__25993),
            .I(N__25974));
    InMux I__5167 (
            .O(N__25990),
            .I(N__25967));
    InMux I__5166 (
            .O(N__25989),
            .I(N__25967));
    InMux I__5165 (
            .O(N__25988),
            .I(N__25967));
    InMux I__5164 (
            .O(N__25987),
            .I(N__25958));
    InMux I__5163 (
            .O(N__25984),
            .I(N__25958));
    InMux I__5162 (
            .O(N__25983),
            .I(N__25958));
    InMux I__5161 (
            .O(N__25980),
            .I(N__25958));
    Odrv4 I__5160 (
            .O(N__25977),
            .I(\POWERLED.N_435_i ));
    Odrv12 I__5159 (
            .O(N__25974),
            .I(\POWERLED.N_435_i ));
    LocalMux I__5158 (
            .O(N__25967),
            .I(\POWERLED.N_435_i ));
    LocalMux I__5157 (
            .O(N__25958),
            .I(\POWERLED.N_435_i ));
    InMux I__5156 (
            .O(N__25949),
            .I(N__25943));
    InMux I__5155 (
            .O(N__25948),
            .I(N__25943));
    LocalMux I__5154 (
            .O(N__25943),
            .I(N__25940));
    Odrv4 I__5153 (
            .O(N__25940),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    InMux I__5152 (
            .O(N__25937),
            .I(\POWERLED.un1_dutycycle_94_cry_13 ));
    InMux I__5151 (
            .O(N__25934),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    InMux I__5150 (
            .O(N__25931),
            .I(N__25925));
    InMux I__5149 (
            .O(N__25930),
            .I(N__25925));
    LocalMux I__5148 (
            .O(N__25925),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    CascadeMux I__5147 (
            .O(N__25922),
            .I(N__25919));
    InMux I__5146 (
            .O(N__25919),
            .I(N__25913));
    InMux I__5145 (
            .O(N__25918),
            .I(N__25913));
    LocalMux I__5144 (
            .O(N__25913),
            .I(N__25910));
    Odrv4 I__5143 (
            .O(N__25910),
            .I(\POWERLED.un1_dutycycle_53_2_1 ));
    CascadeMux I__5142 (
            .O(N__25907),
            .I(N__25904));
    InMux I__5141 (
            .O(N__25904),
            .I(N__25901));
    LocalMux I__5140 (
            .O(N__25901),
            .I(N__25896));
    InMux I__5139 (
            .O(N__25900),
            .I(N__25891));
    InMux I__5138 (
            .O(N__25899),
            .I(N__25891));
    Span4Mux_v I__5137 (
            .O(N__25896),
            .I(N__25888));
    LocalMux I__5136 (
            .O(N__25891),
            .I(N__25885));
    Odrv4 I__5135 (
            .O(N__25888),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_11 ));
    Odrv4 I__5134 (
            .O(N__25885),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_11 ));
    CascadeMux I__5133 (
            .O(N__25880),
            .I(N__25877));
    InMux I__5132 (
            .O(N__25877),
            .I(N__25864));
    InMux I__5131 (
            .O(N__25876),
            .I(N__25861));
    InMux I__5130 (
            .O(N__25875),
            .I(N__25856));
    InMux I__5129 (
            .O(N__25874),
            .I(N__25856));
    InMux I__5128 (
            .O(N__25873),
            .I(N__25853));
    InMux I__5127 (
            .O(N__25872),
            .I(N__25849));
    InMux I__5126 (
            .O(N__25871),
            .I(N__25845));
    InMux I__5125 (
            .O(N__25870),
            .I(N__25842));
    InMux I__5124 (
            .O(N__25869),
            .I(N__25837));
    InMux I__5123 (
            .O(N__25868),
            .I(N__25837));
    CascadeMux I__5122 (
            .O(N__25867),
            .I(N__25832));
    LocalMux I__5121 (
            .O(N__25864),
            .I(N__25823));
    LocalMux I__5120 (
            .O(N__25861),
            .I(N__25823));
    LocalMux I__5119 (
            .O(N__25856),
            .I(N__25823));
    LocalMux I__5118 (
            .O(N__25853),
            .I(N__25823));
    InMux I__5117 (
            .O(N__25852),
            .I(N__25819));
    LocalMux I__5116 (
            .O(N__25849),
            .I(N__25816));
    InMux I__5115 (
            .O(N__25848),
            .I(N__25813));
    LocalMux I__5114 (
            .O(N__25845),
            .I(N__25806));
    LocalMux I__5113 (
            .O(N__25842),
            .I(N__25806));
    LocalMux I__5112 (
            .O(N__25837),
            .I(N__25806));
    InMux I__5111 (
            .O(N__25836),
            .I(N__25799));
    InMux I__5110 (
            .O(N__25835),
            .I(N__25799));
    InMux I__5109 (
            .O(N__25832),
            .I(N__25799));
    Span4Mux_v I__5108 (
            .O(N__25823),
            .I(N__25796));
    InMux I__5107 (
            .O(N__25822),
            .I(N__25793));
    LocalMux I__5106 (
            .O(N__25819),
            .I(dutycycle_RNII6848_0_1));
    Odrv4 I__5105 (
            .O(N__25816),
            .I(dutycycle_RNII6848_0_1));
    LocalMux I__5104 (
            .O(N__25813),
            .I(dutycycle_RNII6848_0_1));
    Odrv4 I__5103 (
            .O(N__25806),
            .I(dutycycle_RNII6848_0_1));
    LocalMux I__5102 (
            .O(N__25799),
            .I(dutycycle_RNII6848_0_1));
    Odrv4 I__5101 (
            .O(N__25796),
            .I(dutycycle_RNII6848_0_1));
    LocalMux I__5100 (
            .O(N__25793),
            .I(dutycycle_RNII6848_0_1));
    InMux I__5099 (
            .O(N__25778),
            .I(N__25775));
    LocalMux I__5098 (
            .O(N__25775),
            .I(N__25772));
    Span4Mux_h I__5097 (
            .O(N__25772),
            .I(N__25769));
    Odrv4 I__5096 (
            .O(N__25769),
            .I(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ));
    InMux I__5095 (
            .O(N__25766),
            .I(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__5094 (
            .O(N__25763),
            .I(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ));
    InMux I__5093 (
            .O(N__25760),
            .I(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ));
    InMux I__5092 (
            .O(N__25757),
            .I(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ));
    InMux I__5091 (
            .O(N__25754),
            .I(N__25751));
    LocalMux I__5090 (
            .O(N__25751),
            .I(N__25748));
    Span12Mux_s8_v I__5089 (
            .O(N__25748),
            .I(N__25745));
    Odrv12 I__5088 (
            .O(N__25745),
            .I(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ));
    InMux I__5087 (
            .O(N__25742),
            .I(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ));
    InMux I__5086 (
            .O(N__25739),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__5085 (
            .O(N__25736),
            .I(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ));
    CascadeMux I__5084 (
            .O(N__25733),
            .I(N__25729));
    InMux I__5083 (
            .O(N__25732),
            .I(N__25724));
    InMux I__5082 (
            .O(N__25729),
            .I(N__25724));
    LocalMux I__5081 (
            .O(N__25724),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ));
    InMux I__5080 (
            .O(N__25721),
            .I(bfn_9_10_0_));
    InMux I__5079 (
            .O(N__25718),
            .I(\POWERLED.un1_dutycycle_94_cry_8 ));
    CascadeMux I__5078 (
            .O(N__25715),
            .I(\POWERLED.g1_0_1_cascade_ ));
    InMux I__5077 (
            .O(N__25712),
            .I(N__25704));
    InMux I__5076 (
            .O(N__25711),
            .I(N__25701));
    InMux I__5075 (
            .O(N__25710),
            .I(N__25696));
    InMux I__5074 (
            .O(N__25709),
            .I(N__25696));
    InMux I__5073 (
            .O(N__25708),
            .I(N__25691));
    InMux I__5072 (
            .O(N__25707),
            .I(N__25691));
    LocalMux I__5071 (
            .O(N__25704),
            .I(N_43));
    LocalMux I__5070 (
            .O(N__25701),
            .I(N_43));
    LocalMux I__5069 (
            .O(N__25696),
            .I(N_43));
    LocalMux I__5068 (
            .O(N__25691),
            .I(N_43));
    InMux I__5067 (
            .O(N__25682),
            .I(N__25679));
    LocalMux I__5066 (
            .O(N__25679),
            .I(\POWERLED.g2_1 ));
    InMux I__5065 (
            .O(N__25676),
            .I(N__25673));
    LocalMux I__5064 (
            .O(N__25673),
            .I(N__25669));
    CascadeMux I__5063 (
            .O(N__25672),
            .I(N__25666));
    Span4Mux_h I__5062 (
            .O(N__25669),
            .I(N__25659));
    InMux I__5061 (
            .O(N__25666),
            .I(N__25656));
    InMux I__5060 (
            .O(N__25665),
            .I(N__25653));
    InMux I__5059 (
            .O(N__25664),
            .I(N__25648));
    InMux I__5058 (
            .O(N__25663),
            .I(N__25648));
    InMux I__5057 (
            .O(N__25662),
            .I(N__25645));
    Span4Mux_h I__5056 (
            .O(N__25659),
            .I(N__25642));
    LocalMux I__5055 (
            .O(N__25656),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__5054 (
            .O(N__25653),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__5053 (
            .O(N__25648),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__5052 (
            .O(N__25645),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__5051 (
            .O(N__25642),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    InMux I__5050 (
            .O(N__25631),
            .I(N__25628));
    LocalMux I__5049 (
            .O(N__25628),
            .I(N__25625));
    Span4Mux_h I__5048 (
            .O(N__25625),
            .I(N__25622));
    Span4Mux_h I__5047 (
            .O(N__25622),
            .I(N__25618));
    InMux I__5046 (
            .O(N__25621),
            .I(N__25615));
    Odrv4 I__5045 (
            .O(N__25618),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    LocalMux I__5044 (
            .O(N__25615),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    InMux I__5043 (
            .O(N__25610),
            .I(N__25607));
    LocalMux I__5042 (
            .O(N__25607),
            .I(N__25603));
    InMux I__5041 (
            .O(N__25606),
            .I(N__25600));
    Span4Mux_s2_h I__5040 (
            .O(N__25603),
            .I(N__25595));
    LocalMux I__5039 (
            .O(N__25600),
            .I(N__25595));
    Span4Mux_v I__5038 (
            .O(N__25595),
            .I(N__25592));
    Span4Mux_h I__5037 (
            .O(N__25592),
            .I(N__25589));
    Odrv4 I__5036 (
            .O(N__25589),
            .I(\PCH_PWRGD.count_0_1 ));
    InMux I__5035 (
            .O(N__25586),
            .I(N__25577));
    CEMux I__5034 (
            .O(N__25585),
            .I(N__25577));
    CascadeMux I__5033 (
            .O(N__25584),
            .I(N__25574));
    CEMux I__5032 (
            .O(N__25583),
            .I(N__25567));
    CEMux I__5031 (
            .O(N__25582),
            .I(N__25563));
    LocalMux I__5030 (
            .O(N__25577),
            .I(N__25557));
    InMux I__5029 (
            .O(N__25574),
            .I(N__25552));
    CEMux I__5028 (
            .O(N__25573),
            .I(N__25552));
    CascadeMux I__5027 (
            .O(N__25572),
            .I(N__25545));
    InMux I__5026 (
            .O(N__25571),
            .I(N__25529));
    CEMux I__5025 (
            .O(N__25570),
            .I(N__25529));
    LocalMux I__5024 (
            .O(N__25567),
            .I(N__25526));
    CEMux I__5023 (
            .O(N__25566),
            .I(N__25523));
    LocalMux I__5022 (
            .O(N__25563),
            .I(N__25520));
    CEMux I__5021 (
            .O(N__25562),
            .I(N__25517));
    InMux I__5020 (
            .O(N__25561),
            .I(N__25512));
    CEMux I__5019 (
            .O(N__25560),
            .I(N__25512));
    Span4Mux_h I__5018 (
            .O(N__25557),
            .I(N__25507));
    LocalMux I__5017 (
            .O(N__25552),
            .I(N__25507));
    InMux I__5016 (
            .O(N__25551),
            .I(N__25498));
    InMux I__5015 (
            .O(N__25550),
            .I(N__25498));
    InMux I__5014 (
            .O(N__25549),
            .I(N__25498));
    InMux I__5013 (
            .O(N__25548),
            .I(N__25498));
    InMux I__5012 (
            .O(N__25545),
            .I(N__25491));
    InMux I__5011 (
            .O(N__25544),
            .I(N__25491));
    InMux I__5010 (
            .O(N__25543),
            .I(N__25491));
    InMux I__5009 (
            .O(N__25542),
            .I(N__25484));
    InMux I__5008 (
            .O(N__25541),
            .I(N__25484));
    InMux I__5007 (
            .O(N__25540),
            .I(N__25484));
    InMux I__5006 (
            .O(N__25539),
            .I(N__25479));
    InMux I__5005 (
            .O(N__25538),
            .I(N__25479));
    InMux I__5004 (
            .O(N__25537),
            .I(N__25470));
    InMux I__5003 (
            .O(N__25536),
            .I(N__25470));
    InMux I__5002 (
            .O(N__25535),
            .I(N__25470));
    InMux I__5001 (
            .O(N__25534),
            .I(N__25470));
    LocalMux I__5000 (
            .O(N__25529),
            .I(N__25464));
    Span4Mux_v I__4999 (
            .O(N__25526),
            .I(N__25461));
    LocalMux I__4998 (
            .O(N__25523),
            .I(N__25452));
    Span4Mux_v I__4997 (
            .O(N__25520),
            .I(N__25452));
    LocalMux I__4996 (
            .O(N__25517),
            .I(N__25452));
    LocalMux I__4995 (
            .O(N__25512),
            .I(N__25452));
    Span4Mux_v I__4994 (
            .O(N__25507),
            .I(N__25447));
    LocalMux I__4993 (
            .O(N__25498),
            .I(N__25447));
    LocalMux I__4992 (
            .O(N__25491),
            .I(N__25438));
    LocalMux I__4991 (
            .O(N__25484),
            .I(N__25438));
    LocalMux I__4990 (
            .O(N__25479),
            .I(N__25438));
    LocalMux I__4989 (
            .O(N__25470),
            .I(N__25438));
    InMux I__4988 (
            .O(N__25469),
            .I(N__25431));
    InMux I__4987 (
            .O(N__25468),
            .I(N__25431));
    InMux I__4986 (
            .O(N__25467),
            .I(N__25431));
    Span12Mux_s4_h I__4985 (
            .O(N__25464),
            .I(N__25428));
    Span4Mux_h I__4984 (
            .O(N__25461),
            .I(N__25417));
    Span4Mux_v I__4983 (
            .O(N__25452),
            .I(N__25417));
    Span4Mux_v I__4982 (
            .O(N__25447),
            .I(N__25417));
    Span4Mux_v I__4981 (
            .O(N__25438),
            .I(N__25417));
    LocalMux I__4980 (
            .O(N__25431),
            .I(N__25417));
    Odrv12 I__4979 (
            .O(N__25428),
            .I(\PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0 ));
    Odrv4 I__4978 (
            .O(N__25417),
            .I(\PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0 ));
    CascadeMux I__4977 (
            .O(N__25412),
            .I(N__25396));
    CascadeMux I__4976 (
            .O(N__25411),
            .I(N__25393));
    CascadeMux I__4975 (
            .O(N__25410),
            .I(N__25387));
    CascadeMux I__4974 (
            .O(N__25409),
            .I(N__25381));
    SRMux I__4973 (
            .O(N__25408),
            .I(N__25377));
    InMux I__4972 (
            .O(N__25407),
            .I(N__25374));
    InMux I__4971 (
            .O(N__25406),
            .I(N__25368));
    SRMux I__4970 (
            .O(N__25405),
            .I(N__25368));
    InMux I__4969 (
            .O(N__25404),
            .I(N__25360));
    SRMux I__4968 (
            .O(N__25403),
            .I(N__25360));
    InMux I__4967 (
            .O(N__25402),
            .I(N__25351));
    InMux I__4966 (
            .O(N__25401),
            .I(N__25351));
    SRMux I__4965 (
            .O(N__25400),
            .I(N__25351));
    InMux I__4964 (
            .O(N__25399),
            .I(N__25351));
    InMux I__4963 (
            .O(N__25396),
            .I(N__25344));
    InMux I__4962 (
            .O(N__25393),
            .I(N__25344));
    InMux I__4961 (
            .O(N__25392),
            .I(N__25344));
    SRMux I__4960 (
            .O(N__25391),
            .I(N__25335));
    InMux I__4959 (
            .O(N__25390),
            .I(N__25335));
    InMux I__4958 (
            .O(N__25387),
            .I(N__25335));
    InMux I__4957 (
            .O(N__25386),
            .I(N__25335));
    InMux I__4956 (
            .O(N__25385),
            .I(N__25326));
    InMux I__4955 (
            .O(N__25384),
            .I(N__25326));
    InMux I__4954 (
            .O(N__25381),
            .I(N__25326));
    InMux I__4953 (
            .O(N__25380),
            .I(N__25326));
    LocalMux I__4952 (
            .O(N__25377),
            .I(N__25323));
    LocalMux I__4951 (
            .O(N__25374),
            .I(N__25320));
    SRMux I__4950 (
            .O(N__25373),
            .I(N__25316));
    LocalMux I__4949 (
            .O(N__25368),
            .I(N__25313));
    InMux I__4948 (
            .O(N__25367),
            .I(N__25307));
    SRMux I__4947 (
            .O(N__25366),
            .I(N__25304));
    SRMux I__4946 (
            .O(N__25365),
            .I(N__25301));
    LocalMux I__4945 (
            .O(N__25360),
            .I(N__25284));
    LocalMux I__4944 (
            .O(N__25351),
            .I(N__25284));
    LocalMux I__4943 (
            .O(N__25344),
            .I(N__25284));
    LocalMux I__4942 (
            .O(N__25335),
            .I(N__25284));
    LocalMux I__4941 (
            .O(N__25326),
            .I(N__25284));
    Span4Mux_v I__4940 (
            .O(N__25323),
            .I(N__25281));
    Span4Mux_v I__4939 (
            .O(N__25320),
            .I(N__25278));
    InMux I__4938 (
            .O(N__25319),
            .I(N__25275));
    LocalMux I__4937 (
            .O(N__25316),
            .I(N__25270));
    Span4Mux_v I__4936 (
            .O(N__25313),
            .I(N__25270));
    InMux I__4935 (
            .O(N__25312),
            .I(N__25267));
    InMux I__4934 (
            .O(N__25311),
            .I(N__25262));
    InMux I__4933 (
            .O(N__25310),
            .I(N__25262));
    LocalMux I__4932 (
            .O(N__25307),
            .I(N__25255));
    LocalMux I__4931 (
            .O(N__25304),
            .I(N__25255));
    LocalMux I__4930 (
            .O(N__25301),
            .I(N__25255));
    InMux I__4929 (
            .O(N__25300),
            .I(N__25252));
    InMux I__4928 (
            .O(N__25299),
            .I(N__25247));
    InMux I__4927 (
            .O(N__25298),
            .I(N__25247));
    InMux I__4926 (
            .O(N__25297),
            .I(N__25240));
    InMux I__4925 (
            .O(N__25296),
            .I(N__25240));
    InMux I__4924 (
            .O(N__25295),
            .I(N__25240));
    Span4Mux_v I__4923 (
            .O(N__25284),
            .I(N__25231));
    Span4Mux_h I__4922 (
            .O(N__25281),
            .I(N__25231));
    Span4Mux_h I__4921 (
            .O(N__25278),
            .I(N__25231));
    LocalMux I__4920 (
            .O(N__25275),
            .I(N__25231));
    Odrv4 I__4919 (
            .O(N__25270),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__4918 (
            .O(N__25267),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__4917 (
            .O(N__25262),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__4916 (
            .O(N__25255),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__4915 (
            .O(N__25252),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__4914 (
            .O(N__25247),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__4913 (
            .O(N__25240),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__4912 (
            .O(N__25231),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    InMux I__4911 (
            .O(N__25214),
            .I(N__25211));
    LocalMux I__4910 (
            .O(N__25211),
            .I(N__25208));
    Span4Mux_v I__4909 (
            .O(N__25208),
            .I(N__25204));
    CascadeMux I__4908 (
            .O(N__25207),
            .I(N__25201));
    Sp12to4 I__4907 (
            .O(N__25204),
            .I(N__25198));
    InMux I__4906 (
            .O(N__25201),
            .I(N__25195));
    Odrv12 I__4905 (
            .O(N__25198),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    LocalMux I__4904 (
            .O(N__25195),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__4903 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__4902 (
            .O(N__25187),
            .I(N__25184));
    Span4Mux_v I__4901 (
            .O(N__25184),
            .I(N__25181));
    Span4Mux_h I__4900 (
            .O(N__25181),
            .I(N__25178));
    Odrv4 I__4899 (
            .O(N__25178),
            .I(\POWERLED.mult1_un124_sum_axb_7_l_fx ));
    InMux I__4898 (
            .O(N__25175),
            .I(N__25169));
    InMux I__4897 (
            .O(N__25174),
            .I(N__25169));
    LocalMux I__4896 (
            .O(N__25169),
            .I(N__25166));
    Span4Mux_v I__4895 (
            .O(N__25166),
            .I(N__25161));
    InMux I__4894 (
            .O(N__25165),
            .I(N__25158));
    CascadeMux I__4893 (
            .O(N__25164),
            .I(N__25155));
    Span4Mux_h I__4892 (
            .O(N__25161),
            .I(N__25147));
    LocalMux I__4891 (
            .O(N__25158),
            .I(N__25147));
    InMux I__4890 (
            .O(N__25155),
            .I(N__25140));
    InMux I__4889 (
            .O(N__25154),
            .I(N__25140));
    InMux I__4888 (
            .O(N__25153),
            .I(N__25140));
    InMux I__4887 (
            .O(N__25152),
            .I(N__25137));
    Odrv4 I__4886 (
            .O(N__25147),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__4885 (
            .O(N__25140),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__4884 (
            .O(N__25137),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    InMux I__4883 (
            .O(N__25130),
            .I(N__25127));
    LocalMux I__4882 (
            .O(N__25127),
            .I(N__25124));
    Span12Mux_s8_v I__4881 (
            .O(N__25124),
            .I(N__25121));
    Odrv12 I__4880 (
            .O(N__25121),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__4879 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__4878 (
            .O(N__25115),
            .I(N__25111));
    InMux I__4877 (
            .O(N__25114),
            .I(N__25108));
    Span12Mux_v I__4876 (
            .O(N__25111),
            .I(N__25101));
    LocalMux I__4875 (
            .O(N__25108),
            .I(N__25101));
    InMux I__4874 (
            .O(N__25107),
            .I(N__25098));
    InMux I__4873 (
            .O(N__25106),
            .I(N__25095));
    Odrv12 I__4872 (
            .O(N__25101),
            .I(N_428));
    LocalMux I__4871 (
            .O(N__25098),
            .I(N_428));
    LocalMux I__4870 (
            .O(N__25095),
            .I(N_428));
    IoInMux I__4869 (
            .O(N__25088),
            .I(N__25085));
    LocalMux I__4868 (
            .O(N__25085),
            .I(N__25081));
    IoInMux I__4867 (
            .O(N__25084),
            .I(N__25078));
    IoSpan4Mux I__4866 (
            .O(N__25081),
            .I(N__25075));
    LocalMux I__4865 (
            .O(N__25078),
            .I(N__25072));
    IoSpan4Mux I__4864 (
            .O(N__25075),
            .I(N__25069));
    Span4Mux_s2_h I__4863 (
            .O(N__25072),
            .I(N__25066));
    Sp12to4 I__4862 (
            .O(N__25069),
            .I(N__25063));
    Span4Mux_v I__4861 (
            .O(N__25066),
            .I(N__25060));
    Odrv12 I__4860 (
            .O(N__25063),
            .I(pch_pwrok));
    Odrv4 I__4859 (
            .O(N__25060),
            .I(pch_pwrok));
    CascadeMux I__4858 (
            .O(N__25055),
            .I(\POWERLED.func_state_RNI12ASZ0Z_1_cascade_ ));
    InMux I__4857 (
            .O(N__25052),
            .I(N__25049));
    LocalMux I__4856 (
            .O(N__25049),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3 ));
    InMux I__4855 (
            .O(N__25046),
            .I(N__25043));
    LocalMux I__4854 (
            .O(N__25043),
            .I(\POWERLED.dutycycle_eena_13 ));
    CascadeMux I__4853 (
            .O(N__25040),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3_cascade_ ));
    InMux I__4852 (
            .O(N__25037),
            .I(N__25031));
    InMux I__4851 (
            .O(N__25036),
            .I(N__25031));
    LocalMux I__4850 (
            .O(N__25031),
            .I(\POWERLED.dutycycle_0_6 ));
    InMux I__4849 (
            .O(N__25028),
            .I(N__25025));
    LocalMux I__4848 (
            .O(N__25025),
            .I(\POWERLED.dutycycle_RNI_13Z0Z_0 ));
    CascadeMux I__4847 (
            .O(N__25022),
            .I(\POWERLED.N_2363_0_cascade_ ));
    InMux I__4846 (
            .O(N__25019),
            .I(N__25016));
    LocalMux I__4845 (
            .O(N__25016),
            .I(\POWERLED.N_12_3_0 ));
    CascadeMux I__4844 (
            .O(N__25013),
            .I(G_11_i_a10_2_1_cascade_));
    CascadeMux I__4843 (
            .O(N__25010),
            .I(N__25007));
    InMux I__4842 (
            .O(N__25007),
            .I(N__25004));
    LocalMux I__4841 (
            .O(N__25004),
            .I(N__25001));
    Span4Mux_h I__4840 (
            .O(N__25001),
            .I(N__24997));
    InMux I__4839 (
            .O(N__25000),
            .I(N__24994));
    Odrv4 I__4838 (
            .O(N__24997),
            .I(\POWERLED.g2_3 ));
    LocalMux I__4837 (
            .O(N__24994),
            .I(\POWERLED.g2_3 ));
    InMux I__4836 (
            .O(N__24989),
            .I(N__24986));
    LocalMux I__4835 (
            .O(N__24986),
            .I(N_28));
    InMux I__4834 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__4833 (
            .O(N__24980),
            .I(N_7));
    CascadeMux I__4832 (
            .O(N__24977),
            .I(N__24973));
    InMux I__4831 (
            .O(N__24976),
            .I(N__24968));
    InMux I__4830 (
            .O(N__24973),
            .I(N__24968));
    LocalMux I__4829 (
            .O(N__24968),
            .I(N__24965));
    Odrv4 I__4828 (
            .O(N__24965),
            .I(N_50));
    CascadeMux I__4827 (
            .O(N__24962),
            .I(N_7_cascade_));
    InMux I__4826 (
            .O(N__24959),
            .I(N__24955));
    InMux I__4825 (
            .O(N__24958),
            .I(N__24952));
    LocalMux I__4824 (
            .O(N__24955),
            .I(N__24949));
    LocalMux I__4823 (
            .O(N__24952),
            .I(\POWERLED.N_2363_0 ));
    Odrv4 I__4822 (
            .O(N__24949),
            .I(\POWERLED.N_2363_0 ));
    InMux I__4821 (
            .O(N__24944),
            .I(N__24941));
    LocalMux I__4820 (
            .O(N__24941),
            .I(N__24937));
    InMux I__4819 (
            .O(N__24940),
            .I(N__24934));
    Odrv4 I__4818 (
            .O(N__24937),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_0 ));
    LocalMux I__4817 (
            .O(N__24934),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_0 ));
    InMux I__4816 (
            .O(N__24929),
            .I(N__24925));
    InMux I__4815 (
            .O(N__24928),
            .I(N__24918));
    LocalMux I__4814 (
            .O(N__24925),
            .I(N__24915));
    InMux I__4813 (
            .O(N__24924),
            .I(N__24912));
    InMux I__4812 (
            .O(N__24923),
            .I(N__24907));
    InMux I__4811 (
            .O(N__24922),
            .I(N__24907));
    InMux I__4810 (
            .O(N__24921),
            .I(N__24904));
    LocalMux I__4809 (
            .O(N__24918),
            .I(N__24901));
    Span4Mux_v I__4808 (
            .O(N__24915),
            .I(N__24898));
    LocalMux I__4807 (
            .O(N__24912),
            .I(N__24891));
    LocalMux I__4806 (
            .O(N__24907),
            .I(N__24891));
    LocalMux I__4805 (
            .O(N__24904),
            .I(N__24891));
    Span4Mux_s3_h I__4804 (
            .O(N__24901),
            .I(N__24884));
    Span4Mux_s3_h I__4803 (
            .O(N__24898),
            .I(N__24884));
    Span4Mux_v I__4802 (
            .O(N__24891),
            .I(N__24884));
    Odrv4 I__4801 (
            .O(N__24884),
            .I(\POWERLED.N_613 ));
    CascadeMux I__4800 (
            .O(N__24881),
            .I(\POWERLED.un1_clk_100khz_51_and_i_3_1_cascade_ ));
    InMux I__4799 (
            .O(N__24878),
            .I(N__24874));
    InMux I__4798 (
            .O(N__24877),
            .I(N__24871));
    LocalMux I__4797 (
            .O(N__24874),
            .I(N__24866));
    LocalMux I__4796 (
            .O(N__24871),
            .I(N__24866));
    Odrv4 I__4795 (
            .O(N__24866),
            .I(\POWERLED.N_252_N ));
    CascadeMux I__4794 (
            .O(N__24863),
            .I(\POWERLED.dutycycle_eena_13_1_cascade_ ));
    CascadeMux I__4793 (
            .O(N__24860),
            .I(\POWERLED.dutycycle_eena_13_cascade_ ));
    InMux I__4792 (
            .O(N__24857),
            .I(N__24854));
    LocalMux I__4791 (
            .O(N__24854),
            .I(N__24851));
    Span4Mux_h I__4790 (
            .O(N__24851),
            .I(N__24848));
    Odrv4 I__4789 (
            .O(N__24848),
            .I(\POWERLED.N_452 ));
    InMux I__4788 (
            .O(N__24845),
            .I(N__24839));
    InMux I__4787 (
            .O(N__24844),
            .I(N__24839));
    LocalMux I__4786 (
            .O(N__24839),
            .I(N__24836));
    Odrv4 I__4785 (
            .O(N__24836),
            .I(\POWERLED.dutycycle_set_1 ));
    InMux I__4784 (
            .O(N__24833),
            .I(N__24830));
    LocalMux I__4783 (
            .O(N__24830),
            .I(\POWERLED.func_state_RNI12ASZ0Z_1 ));
    CascadeMux I__4782 (
            .O(N__24827),
            .I(\POWERLED.dutycycle_e_N_3L4_0_1_cascade_ ));
    InMux I__4781 (
            .O(N__24824),
            .I(N__24821));
    LocalMux I__4780 (
            .O(N__24821),
            .I(\POWERLED.g0_8Z0Z_0 ));
    CascadeMux I__4779 (
            .O(N__24818),
            .I(\POWERLED.N_435_cascade_ ));
    InMux I__4778 (
            .O(N__24815),
            .I(N__24812));
    LocalMux I__4777 (
            .O(N__24812),
            .I(N__24809));
    Odrv4 I__4776 (
            .O(N__24809),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_0 ));
    InMux I__4775 (
            .O(N__24806),
            .I(N__24803));
    LocalMux I__4774 (
            .O(N__24803),
            .I(\POWERLED.func_state_1_m2s2_i_0_0 ));
    CascadeMux I__4773 (
            .O(N__24800),
            .I(\POWERLED.N_423_cascade_ ));
    InMux I__4772 (
            .O(N__24797),
            .I(N__24794));
    LocalMux I__4771 (
            .O(N__24794),
            .I(\POWERLED.N_542 ));
    InMux I__4770 (
            .O(N__24791),
            .I(N__24788));
    LocalMux I__4769 (
            .O(N__24788),
            .I(N__24785));
    Odrv4 I__4768 (
            .O(N__24785),
            .I(\POWERLED.func_stateZ1Z_0 ));
    InMux I__4767 (
            .O(N__24782),
            .I(N__24779));
    LocalMux I__4766 (
            .O(N__24779),
            .I(\POWERLED.g2 ));
    CascadeMux I__4765 (
            .O(N__24776),
            .I(N__24773));
    InMux I__4764 (
            .O(N__24773),
            .I(N__24770));
    LocalMux I__4763 (
            .O(N__24770),
            .I(N__24767));
    Span4Mux_h I__4762 (
            .O(N__24767),
            .I(N__24764));
    Span4Mux_s2_h I__4761 (
            .O(N__24764),
            .I(N__24760));
    InMux I__4760 (
            .O(N__24763),
            .I(N__24757));
    Odrv4 I__4759 (
            .O(N__24760),
            .I(\POWERLED.g0_0_5 ));
    LocalMux I__4758 (
            .O(N__24757),
            .I(\POWERLED.g0_0_5 ));
    InMux I__4757 (
            .O(N__24752),
            .I(N__24748));
    InMux I__4756 (
            .O(N__24751),
            .I(N__24745));
    LocalMux I__4755 (
            .O(N__24748),
            .I(\POWERLED.g2_0 ));
    LocalMux I__4754 (
            .O(N__24745),
            .I(\POWERLED.g2_0 ));
    CascadeMux I__4753 (
            .O(N__24740),
            .I(\POWERLED.g2_cascade_ ));
    InMux I__4752 (
            .O(N__24737),
            .I(N__24731));
    InMux I__4751 (
            .O(N__24736),
            .I(N__24731));
    LocalMux I__4750 (
            .O(N__24731),
            .I(N__24728));
    Span4Mux_h I__4749 (
            .O(N__24728),
            .I(N__24725));
    Odrv4 I__4748 (
            .O(N__24725),
            .I(\POWERLED.N_13_0_0_0 ));
    CascadeMux I__4747 (
            .O(N__24722),
            .I(\POWERLED.func_stateZ0Z_0_cascade_ ));
    InMux I__4746 (
            .O(N__24719),
            .I(N__24714));
    InMux I__4745 (
            .O(N__24718),
            .I(N__24709));
    InMux I__4744 (
            .O(N__24717),
            .I(N__24709));
    LocalMux I__4743 (
            .O(N__24714),
            .I(N__24706));
    LocalMux I__4742 (
            .O(N__24709),
            .I(N__24701));
    Span4Mux_s3_v I__4741 (
            .O(N__24706),
            .I(N__24701));
    Odrv4 I__4740 (
            .O(N__24701),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_0 ));
    InMux I__4739 (
            .O(N__24698),
            .I(N__24684));
    IoInMux I__4738 (
            .O(N__24697),
            .I(N__24680));
    CascadeMux I__4737 (
            .O(N__24696),
            .I(N__24677));
    InMux I__4736 (
            .O(N__24695),
            .I(N__24670));
    InMux I__4735 (
            .O(N__24694),
            .I(N__24670));
    InMux I__4734 (
            .O(N__24693),
            .I(N__24656));
    InMux I__4733 (
            .O(N__24692),
            .I(N__24656));
    CascadeMux I__4732 (
            .O(N__24691),
            .I(N__24650));
    CascadeMux I__4731 (
            .O(N__24690),
            .I(N__24645));
    InMux I__4730 (
            .O(N__24689),
            .I(N__24632));
    InMux I__4729 (
            .O(N__24688),
            .I(N__24632));
    InMux I__4728 (
            .O(N__24687),
            .I(N__24632));
    LocalMux I__4727 (
            .O(N__24684),
            .I(N__24627));
    InMux I__4726 (
            .O(N__24683),
            .I(N__24624));
    LocalMux I__4725 (
            .O(N__24680),
            .I(N__24621));
    InMux I__4724 (
            .O(N__24677),
            .I(N__24617));
    CascadeMux I__4723 (
            .O(N__24676),
            .I(N__24612));
    InMux I__4722 (
            .O(N__24675),
            .I(N__24608));
    LocalMux I__4721 (
            .O(N__24670),
            .I(N__24605));
    InMux I__4720 (
            .O(N__24669),
            .I(N__24602));
    InMux I__4719 (
            .O(N__24668),
            .I(N__24599));
    InMux I__4718 (
            .O(N__24667),
            .I(N__24596));
    InMux I__4717 (
            .O(N__24666),
            .I(N__24591));
    InMux I__4716 (
            .O(N__24665),
            .I(N__24591));
    InMux I__4715 (
            .O(N__24664),
            .I(N__24588));
    InMux I__4714 (
            .O(N__24663),
            .I(N__24581));
    InMux I__4713 (
            .O(N__24662),
            .I(N__24581));
    InMux I__4712 (
            .O(N__24661),
            .I(N__24581));
    LocalMux I__4711 (
            .O(N__24656),
            .I(N__24578));
    InMux I__4710 (
            .O(N__24655),
            .I(N__24565));
    InMux I__4709 (
            .O(N__24654),
            .I(N__24565));
    InMux I__4708 (
            .O(N__24653),
            .I(N__24565));
    InMux I__4707 (
            .O(N__24650),
            .I(N__24565));
    InMux I__4706 (
            .O(N__24649),
            .I(N__24565));
    InMux I__4705 (
            .O(N__24648),
            .I(N__24565));
    InMux I__4704 (
            .O(N__24645),
            .I(N__24556));
    InMux I__4703 (
            .O(N__24644),
            .I(N__24556));
    InMux I__4702 (
            .O(N__24643),
            .I(N__24556));
    InMux I__4701 (
            .O(N__24642),
            .I(N__24556));
    InMux I__4700 (
            .O(N__24641),
            .I(N__24548));
    InMux I__4699 (
            .O(N__24640),
            .I(N__24548));
    InMux I__4698 (
            .O(N__24639),
            .I(N__24548));
    LocalMux I__4697 (
            .O(N__24632),
            .I(N__24545));
    InMux I__4696 (
            .O(N__24631),
            .I(N__24542));
    InMux I__4695 (
            .O(N__24630),
            .I(N__24539));
    Span4Mux_v I__4694 (
            .O(N__24627),
            .I(N__24534));
    LocalMux I__4693 (
            .O(N__24624),
            .I(N__24534));
    IoSpan4Mux I__4692 (
            .O(N__24621),
            .I(N__24531));
    InMux I__4691 (
            .O(N__24620),
            .I(N__24528));
    LocalMux I__4690 (
            .O(N__24617),
            .I(N__24525));
    InMux I__4689 (
            .O(N__24616),
            .I(N__24516));
    InMux I__4688 (
            .O(N__24615),
            .I(N__24516));
    InMux I__4687 (
            .O(N__24612),
            .I(N__24516));
    InMux I__4686 (
            .O(N__24611),
            .I(N__24516));
    LocalMux I__4685 (
            .O(N__24608),
            .I(N__24513));
    Span4Mux_s0_v I__4684 (
            .O(N__24605),
            .I(N__24510));
    LocalMux I__4683 (
            .O(N__24602),
            .I(N__24507));
    LocalMux I__4682 (
            .O(N__24599),
            .I(N__24502));
    LocalMux I__4681 (
            .O(N__24596),
            .I(N__24499));
    LocalMux I__4680 (
            .O(N__24591),
            .I(N__24486));
    LocalMux I__4679 (
            .O(N__24588),
            .I(N__24486));
    LocalMux I__4678 (
            .O(N__24581),
            .I(N__24486));
    Span4Mux_h I__4677 (
            .O(N__24578),
            .I(N__24486));
    LocalMux I__4676 (
            .O(N__24565),
            .I(N__24486));
    LocalMux I__4675 (
            .O(N__24556),
            .I(N__24486));
    InMux I__4674 (
            .O(N__24555),
            .I(N__24483));
    LocalMux I__4673 (
            .O(N__24548),
            .I(N__24476));
    Span4Mux_h I__4672 (
            .O(N__24545),
            .I(N__24476));
    LocalMux I__4671 (
            .O(N__24542),
            .I(N__24476));
    LocalMux I__4670 (
            .O(N__24539),
            .I(N__24471));
    Span4Mux_h I__4669 (
            .O(N__24534),
            .I(N__24471));
    Span4Mux_s2_h I__4668 (
            .O(N__24531),
            .I(N__24466));
    LocalMux I__4667 (
            .O(N__24528),
            .I(N__24466));
    Span4Mux_s2_h I__4666 (
            .O(N__24525),
            .I(N__24461));
    LocalMux I__4665 (
            .O(N__24516),
            .I(N__24461));
    Span4Mux_v I__4664 (
            .O(N__24513),
            .I(N__24454));
    Span4Mux_v I__4663 (
            .O(N__24510),
            .I(N__24454));
    Span4Mux_h I__4662 (
            .O(N__24507),
            .I(N__24454));
    InMux I__4661 (
            .O(N__24506),
            .I(N__24449));
    InMux I__4660 (
            .O(N__24505),
            .I(N__24449));
    Span12Mux_s8_v I__4659 (
            .O(N__24502),
            .I(N__24446));
    Span4Mux_h I__4658 (
            .O(N__24499),
            .I(N__24439));
    Span4Mux_v I__4657 (
            .O(N__24486),
            .I(N__24439));
    LocalMux I__4656 (
            .O(N__24483),
            .I(N__24439));
    Span4Mux_v I__4655 (
            .O(N__24476),
            .I(N__24434));
    Span4Mux_v I__4654 (
            .O(N__24471),
            .I(N__24434));
    Span4Mux_v I__4653 (
            .O(N__24466),
            .I(N__24427));
    Span4Mux_v I__4652 (
            .O(N__24461),
            .I(N__24427));
    Span4Mux_v I__4651 (
            .O(N__24454),
            .I(N__24427));
    LocalMux I__4650 (
            .O(N__24449),
            .I(suswarn_n));
    Odrv12 I__4649 (
            .O(N__24446),
            .I(suswarn_n));
    Odrv4 I__4648 (
            .O(N__24439),
            .I(suswarn_n));
    Odrv4 I__4647 (
            .O(N__24434),
            .I(suswarn_n));
    Odrv4 I__4646 (
            .O(N__24427),
            .I(suswarn_n));
    CascadeMux I__4645 (
            .O(N__24416),
            .I(\POWERLED.N_8_0_cascade_ ));
    InMux I__4644 (
            .O(N__24413),
            .I(N__24410));
    LocalMux I__4643 (
            .O(N__24410),
            .I(N__24407));
    Span4Mux_v I__4642 (
            .O(N__24407),
            .I(N__24404));
    Odrv4 I__4641 (
            .O(N__24404),
            .I(\POWERLED.N_16_2 ));
    CascadeMux I__4640 (
            .O(N__24401),
            .I(\POWERLED.N_423_0_cascade_ ));
    CascadeMux I__4639 (
            .O(N__24398),
            .I(\POWERLED.g1_cascade_ ));
    InMux I__4638 (
            .O(N__24395),
            .I(N__24392));
    LocalMux I__4637 (
            .O(N__24392),
            .I(\POWERLED.g0_0_0 ));
    InMux I__4636 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__4635 (
            .O(N__24386),
            .I(\POWERLED.N_8_0_0 ));
    CascadeMux I__4634 (
            .O(N__24383),
            .I(\POWERLED.g0_0_2_cascade_ ));
    CascadeMux I__4633 (
            .O(N__24380),
            .I(\POWERLED.N_541_cascade_ ));
    InMux I__4632 (
            .O(N__24377),
            .I(N__24373));
    InMux I__4631 (
            .O(N__24376),
            .I(N__24370));
    LocalMux I__4630 (
            .O(N__24373),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__4629 (
            .O(N__24370),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    CascadeMux I__4628 (
            .O(N__24365),
            .I(N__24361));
    InMux I__4627 (
            .O(N__24364),
            .I(N__24358));
    InMux I__4626 (
            .O(N__24361),
            .I(N__24355));
    LocalMux I__4625 (
            .O(N__24358),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__4624 (
            .O(N__24355),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__4623 (
            .O(N__24350),
            .I(N__24346));
    InMux I__4622 (
            .O(N__24349),
            .I(N__24343));
    LocalMux I__4621 (
            .O(N__24346),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__4620 (
            .O(N__24343),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__4619 (
            .O(N__24338),
            .I(N__24335));
    LocalMux I__4618 (
            .O(N__24335),
            .I(N__24332));
    Span4Mux_h I__4617 (
            .O(N__24332),
            .I(N__24329));
    Odrv4 I__4616 (
            .O(N__24329),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11 ));
    CascadeMux I__4615 (
            .O(N__24326),
            .I(\RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ));
    CascadeMux I__4614 (
            .O(N__24323),
            .I(N__24319));
    InMux I__4613 (
            .O(N__24322),
            .I(N__24316));
    InMux I__4612 (
            .O(N__24319),
            .I(N__24313));
    LocalMux I__4611 (
            .O(N__24316),
            .I(\RSMRST_PWRGD.N_264_i ));
    LocalMux I__4610 (
            .O(N__24313),
            .I(\RSMRST_PWRGD.N_264_i ));
    InMux I__4609 (
            .O(N__24308),
            .I(N__24291));
    InMux I__4608 (
            .O(N__24307),
            .I(N__24291));
    InMux I__4607 (
            .O(N__24306),
            .I(N__24291));
    InMux I__4606 (
            .O(N__24305),
            .I(N__24291));
    InMux I__4605 (
            .O(N__24304),
            .I(N__24291));
    CascadeMux I__4604 (
            .O(N__24303),
            .I(N__24288));
    CascadeMux I__4603 (
            .O(N__24302),
            .I(N__24285));
    LocalMux I__4602 (
            .O(N__24291),
            .I(N__24280));
    InMux I__4601 (
            .O(N__24288),
            .I(N__24271));
    InMux I__4600 (
            .O(N__24285),
            .I(N__24271));
    InMux I__4599 (
            .O(N__24284),
            .I(N__24271));
    InMux I__4598 (
            .O(N__24283),
            .I(N__24271));
    Span4Mux_s0_v I__4597 (
            .O(N__24280),
            .I(N__24268));
    LocalMux I__4596 (
            .O(N__24271),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__4595 (
            .O(N__24268),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    InMux I__4594 (
            .O(N__24263),
            .I(N__24251));
    InMux I__4593 (
            .O(N__24262),
            .I(N__24251));
    InMux I__4592 (
            .O(N__24261),
            .I(N__24251));
    InMux I__4591 (
            .O(N__24260),
            .I(N__24251));
    LocalMux I__4590 (
            .O(N__24251),
            .I(N__24248));
    Span4Mux_h I__4589 (
            .O(N__24248),
            .I(N__24239));
    InMux I__4588 (
            .O(N__24247),
            .I(N__24226));
    InMux I__4587 (
            .O(N__24246),
            .I(N__24226));
    InMux I__4586 (
            .O(N__24245),
            .I(N__24226));
    InMux I__4585 (
            .O(N__24244),
            .I(N__24226));
    InMux I__4584 (
            .O(N__24243),
            .I(N__24226));
    InMux I__4583 (
            .O(N__24242),
            .I(N__24226));
    Odrv4 I__4582 (
            .O(N__24239),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__4581 (
            .O(N__24226),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    InMux I__4580 (
            .O(N__24221),
            .I(N__24214));
    InMux I__4579 (
            .O(N__24220),
            .I(N__24214));
    InMux I__4578 (
            .O(N__24219),
            .I(N__24211));
    LocalMux I__4577 (
            .O(N__24214),
            .I(N__24208));
    LocalMux I__4576 (
            .O(N__24211),
            .I(N__24205));
    Span4Mux_s1_v I__4575 (
            .O(N__24208),
            .I(N__24202));
    Odrv4 I__4574 (
            .O(N__24205),
            .I(\RSMRST_PWRGD.N_662 ));
    Odrv4 I__4573 (
            .O(N__24202),
            .I(\RSMRST_PWRGD.N_662 ));
    CascadeMux I__4572 (
            .O(N__24197),
            .I(\RSMRST_PWRGD.N_555_cascade_ ));
    SRMux I__4571 (
            .O(N__24194),
            .I(N__24190));
    SRMux I__4570 (
            .O(N__24193),
            .I(N__24187));
    LocalMux I__4569 (
            .O(N__24190),
            .I(N__24183));
    LocalMux I__4568 (
            .O(N__24187),
            .I(N__24180));
    SRMux I__4567 (
            .O(N__24186),
            .I(N__24177));
    Span4Mux_v I__4566 (
            .O(N__24183),
            .I(N__24170));
    Span4Mux_h I__4565 (
            .O(N__24180),
            .I(N__24170));
    LocalMux I__4564 (
            .O(N__24177),
            .I(N__24170));
    Odrv4 I__4563 (
            .O(N__24170),
            .I(\RSMRST_PWRGD.G_14 ));
    CascadeMux I__4562 (
            .O(N__24167),
            .I(N__24149));
    InMux I__4561 (
            .O(N__24166),
            .I(N__24121));
    InMux I__4560 (
            .O(N__24165),
            .I(N__24121));
    InMux I__4559 (
            .O(N__24164),
            .I(N__24121));
    InMux I__4558 (
            .O(N__24163),
            .I(N__24121));
    InMux I__4557 (
            .O(N__24162),
            .I(N__24114));
    InMux I__4556 (
            .O(N__24161),
            .I(N__24114));
    InMux I__4555 (
            .O(N__24160),
            .I(N__24114));
    InMux I__4554 (
            .O(N__24159),
            .I(N__24105));
    InMux I__4553 (
            .O(N__24158),
            .I(N__24105));
    InMux I__4552 (
            .O(N__24157),
            .I(N__24105));
    InMux I__4551 (
            .O(N__24156),
            .I(N__24105));
    InMux I__4550 (
            .O(N__24155),
            .I(N__24096));
    InMux I__4549 (
            .O(N__24154),
            .I(N__24096));
    InMux I__4548 (
            .O(N__24153),
            .I(N__24096));
    InMux I__4547 (
            .O(N__24152),
            .I(N__24096));
    InMux I__4546 (
            .O(N__24149),
            .I(N__24093));
    InMux I__4545 (
            .O(N__24148),
            .I(N__24084));
    InMux I__4544 (
            .O(N__24147),
            .I(N__24084));
    InMux I__4543 (
            .O(N__24146),
            .I(N__24084));
    InMux I__4542 (
            .O(N__24145),
            .I(N__24084));
    InMux I__4541 (
            .O(N__24144),
            .I(N__24077));
    InMux I__4540 (
            .O(N__24143),
            .I(N__24077));
    InMux I__4539 (
            .O(N__24142),
            .I(N__24077));
    InMux I__4538 (
            .O(N__24141),
            .I(N__24068));
    InMux I__4537 (
            .O(N__24140),
            .I(N__24068));
    InMux I__4536 (
            .O(N__24139),
            .I(N__24068));
    InMux I__4535 (
            .O(N__24138),
            .I(N__24068));
    InMux I__4534 (
            .O(N__24137),
            .I(N__24059));
    InMux I__4533 (
            .O(N__24136),
            .I(N__24059));
    InMux I__4532 (
            .O(N__24135),
            .I(N__24059));
    InMux I__4531 (
            .O(N__24134),
            .I(N__24059));
    InMux I__4530 (
            .O(N__24133),
            .I(N__24054));
    InMux I__4529 (
            .O(N__24132),
            .I(N__24054));
    InMux I__4528 (
            .O(N__24131),
            .I(N__24049));
    InMux I__4527 (
            .O(N__24130),
            .I(N__24049));
    LocalMux I__4526 (
            .O(N__24121),
            .I(N__24044));
    LocalMux I__4525 (
            .O(N__24114),
            .I(N__24041));
    LocalMux I__4524 (
            .O(N__24105),
            .I(N__24032));
    LocalMux I__4523 (
            .O(N__24096),
            .I(N__24029));
    LocalMux I__4522 (
            .O(N__24093),
            .I(N__24025));
    LocalMux I__4521 (
            .O(N__24084),
            .I(N__24022));
    LocalMux I__4520 (
            .O(N__24077),
            .I(N__24019));
    LocalMux I__4519 (
            .O(N__24068),
            .I(N__24016));
    LocalMux I__4518 (
            .O(N__24059),
            .I(N__24013));
    LocalMux I__4517 (
            .O(N__24054),
            .I(N__24010));
    LocalMux I__4516 (
            .O(N__24049),
            .I(N__24007));
    CEMux I__4515 (
            .O(N__24048),
            .I(N__23966));
    CEMux I__4514 (
            .O(N__24047),
            .I(N__23966));
    Glb2LocalMux I__4513 (
            .O(N__24044),
            .I(N__23966));
    Glb2LocalMux I__4512 (
            .O(N__24041),
            .I(N__23966));
    CEMux I__4511 (
            .O(N__24040),
            .I(N__23966));
    CEMux I__4510 (
            .O(N__24039),
            .I(N__23966));
    CEMux I__4509 (
            .O(N__24038),
            .I(N__23966));
    CEMux I__4508 (
            .O(N__24037),
            .I(N__23966));
    CEMux I__4507 (
            .O(N__24036),
            .I(N__23966));
    CEMux I__4506 (
            .O(N__24035),
            .I(N__23966));
    Glb2LocalMux I__4505 (
            .O(N__24032),
            .I(N__23966));
    Glb2LocalMux I__4504 (
            .O(N__24029),
            .I(N__23966));
    CEMux I__4503 (
            .O(N__24028),
            .I(N__23966));
    Glb2LocalMux I__4502 (
            .O(N__24025),
            .I(N__23966));
    Glb2LocalMux I__4501 (
            .O(N__24022),
            .I(N__23966));
    Glb2LocalMux I__4500 (
            .O(N__24019),
            .I(N__23966));
    Glb2LocalMux I__4499 (
            .O(N__24016),
            .I(N__23966));
    Glb2LocalMux I__4498 (
            .O(N__24013),
            .I(N__23966));
    Glb2LocalMux I__4497 (
            .O(N__24010),
            .I(N__23966));
    Glb2LocalMux I__4496 (
            .O(N__24007),
            .I(N__23966));
    GlobalMux I__4495 (
            .O(N__23966),
            .I(N__23963));
    gio2CtrlBuf I__4494 (
            .O(N__23963),
            .I(N_92_g));
    CascadeMux I__4493 (
            .O(N__23960),
            .I(\RSMRST_PWRGD.G_14_cascade_ ));
    CEMux I__4492 (
            .O(N__23957),
            .I(N__23954));
    LocalMux I__4491 (
            .O(N__23954),
            .I(N__23951));
    Span4Mux_h I__4490 (
            .O(N__23951),
            .I(N__23948));
    Odrv4 I__4489 (
            .O(N__23948),
            .I(\RSMRST_PWRGD.N_92_1 ));
    InMux I__4488 (
            .O(N__23945),
            .I(N__23939));
    InMux I__4487 (
            .O(N__23944),
            .I(N__23939));
    LocalMux I__4486 (
            .O(N__23939),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    InMux I__4485 (
            .O(N__23936),
            .I(\POWERLED.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__4484 (
            .O(N__23933),
            .I(bfn_8_16_0_));
    InMux I__4483 (
            .O(N__23930),
            .I(N__23927));
    LocalMux I__4482 (
            .O(N__23927),
            .I(N__23924));
    Span4Mux_s2_v I__4481 (
            .O(N__23924),
            .I(N__23921));
    Odrv4 I__4480 (
            .O(N__23921),
            .I(\POWERLED.un1_count_clk_2_axb_10 ));
    InMux I__4479 (
            .O(N__23918),
            .I(\POWERLED.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__4478 (
            .O(N__23915),
            .I(\POWERLED.un1_count_clk_2_cry_10 ));
    InMux I__4477 (
            .O(N__23912),
            .I(\POWERLED.un1_count_clk_2_cry_11 ));
    InMux I__4476 (
            .O(N__23909),
            .I(N__23903));
    InMux I__4475 (
            .O(N__23908),
            .I(N__23903));
    LocalMux I__4474 (
            .O(N__23903),
            .I(N__23900));
    Odrv4 I__4473 (
            .O(N__23900),
            .I(\POWERLED.count_clk_1_13 ));
    InMux I__4472 (
            .O(N__23897),
            .I(\POWERLED.un1_count_clk_2_cry_12_cZ0 ));
    InMux I__4471 (
            .O(N__23894),
            .I(\POWERLED.un1_count_clk_2_cry_13 ));
    InMux I__4470 (
            .O(N__23891),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    InMux I__4469 (
            .O(N__23888),
            .I(N__23882));
    InMux I__4468 (
            .O(N__23887),
            .I(N__23882));
    LocalMux I__4467 (
            .O(N__23882),
            .I(N__23879));
    Odrv4 I__4466 (
            .O(N__23879),
            .I(\POWERLED.count_clk_1_15 ));
    InMux I__4465 (
            .O(N__23876),
            .I(N__23873));
    LocalMux I__4464 (
            .O(N__23873),
            .I(\POWERLED.un1_count_clk_2_axb_14 ));
    InMux I__4463 (
            .O(N__23870),
            .I(N__23867));
    LocalMux I__4462 (
            .O(N__23867),
            .I(N__23864));
    Odrv4 I__4461 (
            .O(N__23864),
            .I(\POWERLED.count_clk_0_4 ));
    InMux I__4460 (
            .O(N__23861),
            .I(N__23855));
    InMux I__4459 (
            .O(N__23860),
            .I(N__23855));
    LocalMux I__4458 (
            .O(N__23855),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    InMux I__4457 (
            .O(N__23852),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    InMux I__4456 (
            .O(N__23849),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    InMux I__4455 (
            .O(N__23846),
            .I(N__23843));
    LocalMux I__4454 (
            .O(N__23843),
            .I(N__23839));
    InMux I__4453 (
            .O(N__23842),
            .I(N__23836));
    Span4Mux_h I__4452 (
            .O(N__23839),
            .I(N__23833));
    LocalMux I__4451 (
            .O(N__23836),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    Odrv4 I__4450 (
            .O(N__23833),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    InMux I__4449 (
            .O(N__23828),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__4448 (
            .O(N__23825),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__4447 (
            .O(N__23822),
            .I(N__23818));
    InMux I__4446 (
            .O(N__23821),
            .I(N__23815));
    LocalMux I__4445 (
            .O(N__23818),
            .I(N__23812));
    LocalMux I__4444 (
            .O(N__23815),
            .I(N__23809));
    Span12Mux_s7_h I__4443 (
            .O(N__23812),
            .I(N__23806));
    Span4Mux_h I__4442 (
            .O(N__23809),
            .I(N__23803));
    Odrv12 I__4441 (
            .O(N__23806),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    Odrv4 I__4440 (
            .O(N__23803),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    InMux I__4439 (
            .O(N__23798),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    InMux I__4438 (
            .O(N__23795),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__4437 (
            .O(N__23792),
            .I(N__23784));
    InMux I__4436 (
            .O(N__23791),
            .I(N__23784));
    InMux I__4435 (
            .O(N__23790),
            .I(N__23779));
    InMux I__4434 (
            .O(N__23789),
            .I(N__23779));
    LocalMux I__4433 (
            .O(N__23784),
            .I(N__23776));
    LocalMux I__4432 (
            .O(N__23779),
            .I(N__23773));
    Odrv4 I__4431 (
            .O(N__23776),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_6 ));
    Odrv4 I__4430 (
            .O(N__23773),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_6 ));
    InMux I__4429 (
            .O(N__23768),
            .I(N__23765));
    LocalMux I__4428 (
            .O(N__23765),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_8 ));
    InMux I__4427 (
            .O(N__23762),
            .I(N__23756));
    InMux I__4426 (
            .O(N__23761),
            .I(N__23756));
    LocalMux I__4425 (
            .O(N__23756),
            .I(\POWERLED.dutycycleZ1Z_14 ));
    CascadeMux I__4424 (
            .O(N__23753),
            .I(\POWERLED.dutycycleZ0Z_10_cascade_ ));
    InMux I__4423 (
            .O(N__23750),
            .I(N__23746));
    InMux I__4422 (
            .O(N__23749),
            .I(N__23743));
    LocalMux I__4421 (
            .O(N__23746),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_13 ));
    LocalMux I__4420 (
            .O(N__23743),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_13 ));
    CascadeMux I__4419 (
            .O(N__23738),
            .I(N__23735));
    InMux I__4418 (
            .O(N__23735),
            .I(N__23732));
    LocalMux I__4417 (
            .O(N__23732),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_15 ));
    InMux I__4416 (
            .O(N__23729),
            .I(N__23726));
    LocalMux I__4415 (
            .O(N__23726),
            .I(\POWERLED.count_clk_0_13 ));
    InMux I__4414 (
            .O(N__23723),
            .I(N__23720));
    LocalMux I__4413 (
            .O(N__23720),
            .I(N__23717));
    Span12Mux_s3_v I__4412 (
            .O(N__23717),
            .I(N__23714));
    Odrv12 I__4411 (
            .O(N__23714),
            .I(\POWERLED.N_492 ));
    CascadeMux I__4410 (
            .O(N__23711),
            .I(\POWERLED.count_clk_en_cascade_ ));
    InMux I__4409 (
            .O(N__23708),
            .I(N__23705));
    LocalMux I__4408 (
            .O(N__23705),
            .I(\POWERLED.count_clk_0_2 ));
    InMux I__4407 (
            .O(N__23702),
            .I(N__23699));
    LocalMux I__4406 (
            .O(N__23699),
            .I(\POWERLED.count_clk_0_15 ));
    CascadeMux I__4405 (
            .O(N__23696),
            .I(\POWERLED.dutycycle_RNI_15Z0Z_3_cascade_ ));
    CascadeMux I__4404 (
            .O(N__23693),
            .I(N__23690));
    InMux I__4403 (
            .O(N__23690),
            .I(N__23687));
    LocalMux I__4402 (
            .O(N__23687),
            .I(\POWERLED.dutycycle_RNIZ0Z_15 ));
    CascadeMux I__4401 (
            .O(N__23684),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_6_cascade_ ));
    CascadeMux I__4400 (
            .O(N__23681),
            .I(N__23678));
    InMux I__4399 (
            .O(N__23678),
            .I(N__23675));
    LocalMux I__4398 (
            .O(N__23675),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_10 ));
    InMux I__4397 (
            .O(N__23672),
            .I(N__23669));
    LocalMux I__4396 (
            .O(N__23669),
            .I(\POWERLED.N_4_0 ));
    CascadeMux I__4395 (
            .O(N__23666),
            .I(N__23663));
    InMux I__4394 (
            .O(N__23663),
            .I(N__23660));
    LocalMux I__4393 (
            .O(N__23660),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_13 ));
    CascadeMux I__4392 (
            .O(N__23657),
            .I(\POWERLED.un1_dutycycle_53_12_1_0_cascade_ ));
    CascadeMux I__4391 (
            .O(N__23654),
            .I(N__23651));
    InMux I__4390 (
            .O(N__23651),
            .I(N__23645));
    InMux I__4389 (
            .O(N__23650),
            .I(N__23645));
    LocalMux I__4388 (
            .O(N__23645),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    InMux I__4387 (
            .O(N__23642),
            .I(N__23636));
    InMux I__4386 (
            .O(N__23641),
            .I(N__23636));
    LocalMux I__4385 (
            .O(N__23636),
            .I(N__23633));
    Odrv4 I__4384 (
            .O(N__23633),
            .I(\POWERLED.dutycycle_RNIT70K5Z0Z_8 ));
    CascadeMux I__4383 (
            .O(N__23630),
            .I(\POWERLED.dutycycleZ0Z_3_cascade_ ));
    CascadeMux I__4382 (
            .O(N__23627),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8_cascade_ ));
    CascadeMux I__4381 (
            .O(N__23624),
            .I(\POWERLED.N_6_3_cascade_ ));
    InMux I__4380 (
            .O(N__23621),
            .I(N__23618));
    LocalMux I__4379 (
            .O(N__23618),
            .I(\POWERLED.g0_9_1_0 ));
    CascadeMux I__4378 (
            .O(N__23615),
            .I(\POWERLED.N_9_1_cascade_ ));
    CascadeMux I__4377 (
            .O(N__23612),
            .I(\POWERLED.un1_m2_e_1_cascade_ ));
    InMux I__4376 (
            .O(N__23609),
            .I(N__23606));
    LocalMux I__4375 (
            .O(N__23606),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_8 ));
    InMux I__4374 (
            .O(N__23603),
            .I(N__23597));
    InMux I__4373 (
            .O(N__23602),
            .I(N__23597));
    LocalMux I__4372 (
            .O(N__23597),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__4371 (
            .O(N__23594),
            .I(\POWERLED.dutycycleZ0Z_7_cascade_ ));
    CascadeMux I__4370 (
            .O(N__23591),
            .I(\POWERLED.un1_dutycycle_53_56_a1_2_cascade_ ));
    CascadeMux I__4369 (
            .O(N__23588),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_8_cascade_ ));
    InMux I__4368 (
            .O(N__23585),
            .I(N__23582));
    LocalMux I__4367 (
            .O(N__23582),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_8 ));
    InMux I__4366 (
            .O(N__23579),
            .I(N__23576));
    LocalMux I__4365 (
            .O(N__23576),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_8 ));
    InMux I__4364 (
            .O(N__23573),
            .I(N__23567));
    InMux I__4363 (
            .O(N__23572),
            .I(N__23567));
    LocalMux I__4362 (
            .O(N__23567),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    CascadeMux I__4361 (
            .O(N__23564),
            .I(N__23561));
    InMux I__4360 (
            .O(N__23561),
            .I(N__23555));
    InMux I__4359 (
            .O(N__23560),
            .I(N__23555));
    LocalMux I__4358 (
            .O(N__23555),
            .I(N_16_0));
    InMux I__4357 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__4356 (
            .O(N__23549),
            .I(N__23546));
    Odrv4 I__4355 (
            .O(N__23546),
            .I(\POWERLED.g0_0_1 ));
    CascadeMux I__4354 (
            .O(N__23543),
            .I(\POWERLED.N_598_cascade_ ));
    CascadeMux I__4353 (
            .O(N__23540),
            .I(\POWERLED.N_450_cascade_ ));
    InMux I__4352 (
            .O(N__23537),
            .I(N__23534));
    LocalMux I__4351 (
            .O(N__23534),
            .I(\POWERLED.dutycycle_RNI5FJ65Z0Z_13 ));
    CascadeMux I__4350 (
            .O(N__23531),
            .I(N__23528));
    InMux I__4349 (
            .O(N__23528),
            .I(N__23522));
    InMux I__4348 (
            .O(N__23527),
            .I(N__23522));
    LocalMux I__4347 (
            .O(N__23522),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    CascadeMux I__4346 (
            .O(N__23519),
            .I(\POWERLED.dutycycle_RNI5FJ65Z0Z_13_cascade_ ));
    CascadeMux I__4345 (
            .O(N__23516),
            .I(\POWERLED.dutycycleZ0Z_11_cascade_ ));
    InMux I__4344 (
            .O(N__23513),
            .I(N__23509));
    InMux I__4343 (
            .O(N__23512),
            .I(N__23506));
    LocalMux I__4342 (
            .O(N__23509),
            .I(\POWERLED.N_2336_i ));
    LocalMux I__4341 (
            .O(N__23506),
            .I(\POWERLED.N_2336_i ));
    InMux I__4340 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__4339 (
            .O(N__23498),
            .I(\POWERLED.N_449 ));
    InMux I__4338 (
            .O(N__23495),
            .I(N__23492));
    LocalMux I__4337 (
            .O(N__23492),
            .I(G_11_i_a10_0_1));
    CascadeMux I__4336 (
            .O(N__23489),
            .I(N_8_3_cascade_));
    InMux I__4335 (
            .O(N__23486),
            .I(N__23483));
    LocalMux I__4334 (
            .O(N__23483),
            .I(\POWERLED.N_10_1 ));
    InMux I__4333 (
            .O(N__23480),
            .I(N__23477));
    LocalMux I__4332 (
            .O(N__23477),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_1 ));
    InMux I__4331 (
            .O(N__23474),
            .I(N__23468));
    InMux I__4330 (
            .O(N__23473),
            .I(N__23468));
    LocalMux I__4329 (
            .O(N__23468),
            .I(\POWERLED.dutycycle_0_5 ));
    CascadeMux I__4328 (
            .O(N__23465),
            .I(N__23461));
    InMux I__4327 (
            .O(N__23464),
            .I(N__23456));
    InMux I__4326 (
            .O(N__23461),
            .I(N__23456));
    LocalMux I__4325 (
            .O(N__23456),
            .I(\POWERLED.g0_i_o4_2 ));
    CascadeMux I__4324 (
            .O(N__23453),
            .I(\POWERLED.dutycycleZ1Z_5_cascade_ ));
    InMux I__4323 (
            .O(N__23450),
            .I(N__23441));
    InMux I__4322 (
            .O(N__23449),
            .I(N__23441));
    InMux I__4321 (
            .O(N__23448),
            .I(N__23441));
    LocalMux I__4320 (
            .O(N__23441),
            .I(\POWERLED.N_546 ));
    CascadeMux I__4319 (
            .O(N__23438),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3_cascade_ ));
    CascadeMux I__4318 (
            .O(N__23435),
            .I(N__23432));
    InMux I__4317 (
            .O(N__23432),
            .I(N__23429));
    LocalMux I__4316 (
            .O(N__23429),
            .I(N__23426));
    Odrv4 I__4315 (
            .O(N__23426),
            .I(\POWERLED.dutycycle_RNIZ0Z_5 ));
    InMux I__4314 (
            .O(N__23423),
            .I(N__23417));
    InMux I__4313 (
            .O(N__23422),
            .I(N__23414));
    InMux I__4312 (
            .O(N__23421),
            .I(N__23409));
    InMux I__4311 (
            .O(N__23420),
            .I(N__23409));
    LocalMux I__4310 (
            .O(N__23417),
            .I(N__23404));
    LocalMux I__4309 (
            .O(N__23414),
            .I(N__23404));
    LocalMux I__4308 (
            .O(N__23409),
            .I(\POWERLED.N_612 ));
    Odrv12 I__4307 (
            .O(N__23404),
            .I(\POWERLED.N_612 ));
    CascadeMux I__4306 (
            .O(N__23399),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_0_cascade_ ));
    CascadeMux I__4305 (
            .O(N__23396),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_0_cascade_ ));
    CascadeMux I__4304 (
            .O(N__23393),
            .I(\POWERLED.N_676_cascade_ ));
    CascadeMux I__4303 (
            .O(N__23390),
            .I(G_11_i_a10_0_1_cascade_));
    InMux I__4302 (
            .O(N__23387),
            .I(N__23384));
    LocalMux I__4301 (
            .O(N__23384),
            .I(G_11_i_2));
    CascadeMux I__4300 (
            .O(N__23381),
            .I(N_9_2_cascade_));
    InMux I__4299 (
            .O(N__23378),
            .I(N__23375));
    LocalMux I__4298 (
            .O(N__23375),
            .I(N_8_3));
    CascadeMux I__4297 (
            .O(N__23372),
            .I(\POWERLED.N_413_N_cascade_ ));
    InMux I__4296 (
            .O(N__23369),
            .I(N__23363));
    InMux I__4295 (
            .O(N__23368),
            .I(N__23363));
    LocalMux I__4294 (
            .O(N__23363),
            .I(\POWERLED.dutycycle_eena ));
    InMux I__4293 (
            .O(N__23360),
            .I(N__23356));
    InMux I__4292 (
            .O(N__23359),
            .I(N__23353));
    LocalMux I__4291 (
            .O(N__23356),
            .I(N__23348));
    LocalMux I__4290 (
            .O(N__23353),
            .I(N__23348));
    Odrv4 I__4289 (
            .O(N__23348),
            .I(\POWERLED.N_413_N ));
    CascadeMux I__4288 (
            .O(N__23345),
            .I(\POWERLED.N_430_cascade_ ));
    CascadeMux I__4287 (
            .O(N__23342),
            .I(N__23339));
    InMux I__4286 (
            .O(N__23339),
            .I(N__23333));
    InMux I__4285 (
            .O(N__23338),
            .I(N__23333));
    LocalMux I__4284 (
            .O(N__23333),
            .I(\POWERLED.dutycycle_eena_1 ));
    InMux I__4283 (
            .O(N__23330),
            .I(N__23321));
    InMux I__4282 (
            .O(N__23329),
            .I(N__23321));
    InMux I__4281 (
            .O(N__23328),
            .I(N__23321));
    LocalMux I__4280 (
            .O(N__23321),
            .I(SUSWARN_N_fast));
    CascadeMux I__4279 (
            .O(N__23318),
            .I(N__23315));
    InMux I__4278 (
            .O(N__23315),
            .I(N__23312));
    LocalMux I__4277 (
            .O(N__23312),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m0 ));
    CascadeMux I__4276 (
            .O(N__23309),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m1_ns_1_cascade_ ));
    InMux I__4275 (
            .O(N__23306),
            .I(N__23303));
    LocalMux I__4274 (
            .O(N__23303),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m1 ));
    CascadeMux I__4273 (
            .O(N__23300),
            .I(N__23297));
    InMux I__4272 (
            .O(N__23297),
            .I(N__23294));
    LocalMux I__4271 (
            .O(N__23294),
            .I(\COUNTER.tmp_0_fast_RNI0RLUZ0Z1 ));
    InMux I__4270 (
            .O(N__23291),
            .I(bfn_8_3_0_));
    InMux I__4269 (
            .O(N__23288),
            .I(N__23284));
    InMux I__4268 (
            .O(N__23287),
            .I(N__23281));
    LocalMux I__4267 (
            .O(N__23284),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__4266 (
            .O(N__23281),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    CascadeMux I__4265 (
            .O(N__23276),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    InMux I__4264 (
            .O(N__23273),
            .I(N__23269));
    InMux I__4263 (
            .O(N__23272),
            .I(N__23266));
    LocalMux I__4262 (
            .O(N__23269),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__4261 (
            .O(N__23266),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__4260 (
            .O(N__23261),
            .I(bfn_8_2_0_));
    InMux I__4259 (
            .O(N__23258),
            .I(N__23254));
    InMux I__4258 (
            .O(N__23257),
            .I(N__23251));
    LocalMux I__4257 (
            .O(N__23254),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__4256 (
            .O(N__23251),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__4255 (
            .O(N__23246),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__4254 (
            .O(N__23243),
            .I(N__23239));
    InMux I__4253 (
            .O(N__23242),
            .I(N__23236));
    LocalMux I__4252 (
            .O(N__23239),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    LocalMux I__4251 (
            .O(N__23236),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__4250 (
            .O(N__23231),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__4249 (
            .O(N__23228),
            .I(N__23224));
    InMux I__4248 (
            .O(N__23227),
            .I(N__23221));
    LocalMux I__4247 (
            .O(N__23224),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__4246 (
            .O(N__23221),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__4245 (
            .O(N__23216),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    InMux I__4244 (
            .O(N__23213),
            .I(N__23209));
    InMux I__4243 (
            .O(N__23212),
            .I(N__23206));
    LocalMux I__4242 (
            .O(N__23209),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__4241 (
            .O(N__23206),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__4240 (
            .O(N__23201),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__4239 (
            .O(N__23198),
            .I(N__23194));
    InMux I__4238 (
            .O(N__23197),
            .I(N__23191));
    LocalMux I__4237 (
            .O(N__23194),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__4236 (
            .O(N__23191),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__4235 (
            .O(N__23186),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__4234 (
            .O(N__23183),
            .I(N__23179));
    InMux I__4233 (
            .O(N__23182),
            .I(N__23176));
    LocalMux I__4232 (
            .O(N__23179),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__4231 (
            .O(N__23176),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__4230 (
            .O(N__23171),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    CascadeMux I__4229 (
            .O(N__23168),
            .I(N__23164));
    InMux I__4228 (
            .O(N__23167),
            .I(N__23160));
    InMux I__4227 (
            .O(N__23164),
            .I(N__23155));
    InMux I__4226 (
            .O(N__23163),
            .I(N__23155));
    LocalMux I__4225 (
            .O(N__23160),
            .I(N__23152));
    LocalMux I__4224 (
            .O(N__23155),
            .I(N__23149));
    Span4Mux_h I__4223 (
            .O(N__23152),
            .I(N__23142));
    Span4Mux_h I__4222 (
            .O(N__23149),
            .I(N__23142));
    InMux I__4221 (
            .O(N__23148),
            .I(N__23139));
    InMux I__4220 (
            .O(N__23147),
            .I(N__23136));
    IoSpan4Mux I__4219 (
            .O(N__23142),
            .I(N__23131));
    LocalMux I__4218 (
            .O(N__23139),
            .I(N__23126));
    LocalMux I__4217 (
            .O(N__23136),
            .I(N__23126));
    IoInMux I__4216 (
            .O(N__23135),
            .I(N__23123));
    InMux I__4215 (
            .O(N__23134),
            .I(N__23120));
    Span4Mux_s3_v I__4214 (
            .O(N__23131),
            .I(N__23115));
    Span4Mux_s3_v I__4213 (
            .O(N__23126),
            .I(N__23115));
    LocalMux I__4212 (
            .O(N__23123),
            .I(N__23112));
    LocalMux I__4211 (
            .O(N__23120),
            .I(N__23109));
    Span4Mux_v I__4210 (
            .O(N__23115),
            .I(N__23106));
    Span12Mux_s4_h I__4209 (
            .O(N__23112),
            .I(N__23103));
    Span4Mux_h I__4208 (
            .O(N__23109),
            .I(N__23100));
    Odrv4 I__4207 (
            .O(N__23106),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4206 (
            .O(N__23103),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4205 (
            .O(N__23100),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4204 (
            .O(N__23093),
            .I(N__23089));
    InMux I__4203 (
            .O(N__23092),
            .I(N__23086));
    InMux I__4202 (
            .O(N__23089),
            .I(N__23083));
    LocalMux I__4201 (
            .O(N__23086),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__4200 (
            .O(N__23083),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    CascadeMux I__4199 (
            .O(N__23078),
            .I(N__23074));
    InMux I__4198 (
            .O(N__23077),
            .I(N__23071));
    InMux I__4197 (
            .O(N__23074),
            .I(N__23068));
    LocalMux I__4196 (
            .O(N__23071),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__4195 (
            .O(N__23068),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    InMux I__4194 (
            .O(N__23063),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__4193 (
            .O(N__23060),
            .I(N__23056));
    InMux I__4192 (
            .O(N__23059),
            .I(N__23053));
    LocalMux I__4191 (
            .O(N__23056),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__4190 (
            .O(N__23053),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__4189 (
            .O(N__23048),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    InMux I__4188 (
            .O(N__23045),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__4187 (
            .O(N__23042),
            .I(N__23038));
    InMux I__4186 (
            .O(N__23041),
            .I(N__23035));
    LocalMux I__4185 (
            .O(N__23038),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__4184 (
            .O(N__23035),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__4183 (
            .O(N__23030),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__4182 (
            .O(N__23027),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__4181 (
            .O(N__23024),
            .I(N__23020));
    InMux I__4180 (
            .O(N__23023),
            .I(N__23017));
    LocalMux I__4179 (
            .O(N__23020),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__4178 (
            .O(N__23017),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__4177 (
            .O(N__23012),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__4176 (
            .O(N__23009),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    CascadeMux I__4175 (
            .O(N__23006),
            .I(N__23003));
    InMux I__4174 (
            .O(N__23003),
            .I(N__22999));
    InMux I__4173 (
            .O(N__23002),
            .I(N__22996));
    LocalMux I__4172 (
            .O(N__22999),
            .I(N__22993));
    LocalMux I__4171 (
            .O(N__22996),
            .I(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ));
    Odrv4 I__4170 (
            .O(N__22993),
            .I(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ));
    InMux I__4169 (
            .O(N__22988),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__4168 (
            .O(N__22985),
            .I(N__22982));
    InMux I__4167 (
            .O(N__22982),
            .I(N__22979));
    LocalMux I__4166 (
            .O(N__22979),
            .I(\POWERLED.mult1_un47_sum_axb_4 ));
    CascadeMux I__4165 (
            .O(N__22976),
            .I(N__22973));
    InMux I__4164 (
            .O(N__22973),
            .I(N__22970));
    LocalMux I__4163 (
            .O(N__22970),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__4162 (
            .O(N__22967),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__4161 (
            .O(N__22964),
            .I(N__22961));
    InMux I__4160 (
            .O(N__22961),
            .I(N__22958));
    LocalMux I__4159 (
            .O(N__22958),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__4158 (
            .O(N__22955),
            .I(N__22952));
    InMux I__4157 (
            .O(N__22952),
            .I(N__22949));
    LocalMux I__4156 (
            .O(N__22949),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__4155 (
            .O(N__22946),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__4154 (
            .O(N__22943),
            .I(N__22940));
    LocalMux I__4153 (
            .O(N__22940),
            .I(N__22937));
    Odrv4 I__4152 (
            .O(N__22937),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_5 ));
    InMux I__4151 (
            .O(N__22934),
            .I(N__22927));
    InMux I__4150 (
            .O(N__22933),
            .I(N__22927));
    InMux I__4149 (
            .O(N__22932),
            .I(N__22924));
    LocalMux I__4148 (
            .O(N__22927),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__4147 (
            .O(N__22924),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    InMux I__4146 (
            .O(N__22919),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    CascadeMux I__4145 (
            .O(N__22916),
            .I(N__22913));
    InMux I__4144 (
            .O(N__22913),
            .I(N__22910));
    LocalMux I__4143 (
            .O(N__22910),
            .I(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__4142 (
            .O(N__22907),
            .I(\POWERLED.mult1_un47_sum_cry_6 ));
    CascadeMux I__4141 (
            .O(N__22904),
            .I(N__22901));
    InMux I__4140 (
            .O(N__22901),
            .I(N__22893));
    InMux I__4139 (
            .O(N__22900),
            .I(N__22893));
    InMux I__4138 (
            .O(N__22899),
            .I(N__22890));
    InMux I__4137 (
            .O(N__22898),
            .I(N__22887));
    LocalMux I__4136 (
            .O(N__22893),
            .I(N__22882));
    LocalMux I__4135 (
            .O(N__22890),
            .I(N__22882));
    LocalMux I__4134 (
            .O(N__22887),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    Odrv4 I__4133 (
            .O(N__22882),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__4132 (
            .O(N__22877),
            .I(N__22874));
    InMux I__4131 (
            .O(N__22874),
            .I(N__22864));
    InMux I__4130 (
            .O(N__22873),
            .I(N__22864));
    InMux I__4129 (
            .O(N__22872),
            .I(N__22864));
    InMux I__4128 (
            .O(N__22871),
            .I(N__22861));
    LocalMux I__4127 (
            .O(N__22864),
            .I(N__22856));
    LocalMux I__4126 (
            .O(N__22861),
            .I(N__22856));
    Odrv4 I__4125 (
            .O(N__22856),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    CascadeMux I__4124 (
            .O(N__22853),
            .I(N__22850));
    InMux I__4123 (
            .O(N__22850),
            .I(N__22847));
    LocalMux I__4122 (
            .O(N__22847),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    InMux I__4121 (
            .O(N__22844),
            .I(N__22839));
    InMux I__4120 (
            .O(N__22843),
            .I(N__22836));
    InMux I__4119 (
            .O(N__22842),
            .I(N__22833));
    LocalMux I__4118 (
            .O(N__22839),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__4117 (
            .O(N__22836),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__4116 (
            .O(N__22833),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    CascadeMux I__4115 (
            .O(N__22826),
            .I(N__22823));
    InMux I__4114 (
            .O(N__22823),
            .I(N__22820));
    LocalMux I__4113 (
            .O(N__22820),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    CascadeMux I__4112 (
            .O(N__22817),
            .I(N__22814));
    InMux I__4111 (
            .O(N__22814),
            .I(N__22811));
    LocalMux I__4110 (
            .O(N__22811),
            .I(N__22808));
    Span4Mux_s3_v I__4109 (
            .O(N__22808),
            .I(N__22805));
    Odrv4 I__4108 (
            .O(N__22805),
            .I(\POWERLED.un1_dutycycle_53_i_28 ));
    CascadeMux I__4107 (
            .O(N__22802),
            .I(N__22798));
    CascadeMux I__4106 (
            .O(N__22801),
            .I(N__22794));
    InMux I__4105 (
            .O(N__22798),
            .I(N__22787));
    InMux I__4104 (
            .O(N__22797),
            .I(N__22787));
    InMux I__4103 (
            .O(N__22794),
            .I(N__22787));
    LocalMux I__4102 (
            .O(N__22787),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    CascadeMux I__4101 (
            .O(N__22784),
            .I(N__22781));
    InMux I__4100 (
            .O(N__22781),
            .I(N__22778));
    LocalMux I__4099 (
            .O(N__22778),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_14 ));
    InMux I__4098 (
            .O(N__22775),
            .I(N__22772));
    LocalMux I__4097 (
            .O(N__22772),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__4096 (
            .O(N__22769),
            .I(N__22763));
    InMux I__4095 (
            .O(N__22768),
            .I(N__22763));
    LocalMux I__4094 (
            .O(N__22763),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__4093 (
            .O(N__22760),
            .I(N__22755));
    CascadeMux I__4092 (
            .O(N__22759),
            .I(N__22752));
    InMux I__4091 (
            .O(N__22758),
            .I(N__22745));
    InMux I__4090 (
            .O(N__22755),
            .I(N__22745));
    InMux I__4089 (
            .O(N__22752),
            .I(N__22745));
    LocalMux I__4088 (
            .O(N__22745),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    InMux I__4087 (
            .O(N__22742),
            .I(N__22739));
    LocalMux I__4086 (
            .O(N__22739),
            .I(N__22735));
    InMux I__4085 (
            .O(N__22738),
            .I(N__22732));
    Span4Mux_v I__4084 (
            .O(N__22735),
            .I(N__22729));
    LocalMux I__4083 (
            .O(N__22732),
            .I(N__22726));
    Odrv4 I__4082 (
            .O(N__22729),
            .I(\POWERLED.mult1_un75_sum ));
    Odrv4 I__4081 (
            .O(N__22726),
            .I(\POWERLED.mult1_un75_sum ));
    InMux I__4080 (
            .O(N__22721),
            .I(\POWERLED.un1_dutycycle_53_cry_9 ));
    InMux I__4079 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__4078 (
            .O(N__22715),
            .I(N__22711));
    InMux I__4077 (
            .O(N__22714),
            .I(N__22708));
    Odrv4 I__4076 (
            .O(N__22711),
            .I(\POWERLED.mult1_un68_sum ));
    LocalMux I__4075 (
            .O(N__22708),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__4074 (
            .O(N__22703),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    InMux I__4073 (
            .O(N__22700),
            .I(N__22697));
    LocalMux I__4072 (
            .O(N__22697),
            .I(N__22693));
    InMux I__4071 (
            .O(N__22696),
            .I(N__22690));
    Odrv4 I__4070 (
            .O(N__22693),
            .I(\POWERLED.mult1_un61_sum ));
    LocalMux I__4069 (
            .O(N__22690),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__4068 (
            .O(N__22685),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    CascadeMux I__4067 (
            .O(N__22682),
            .I(N__22679));
    InMux I__4066 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__4065 (
            .O(N__22676),
            .I(N__22673));
    Odrv4 I__4064 (
            .O(N__22673),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    CascadeMux I__4063 (
            .O(N__22670),
            .I(N__22667));
    InMux I__4062 (
            .O(N__22667),
            .I(N__22663));
    InMux I__4061 (
            .O(N__22666),
            .I(N__22660));
    LocalMux I__4060 (
            .O(N__22663),
            .I(N__22657));
    LocalMux I__4059 (
            .O(N__22660),
            .I(\POWERLED.mult1_un54_sum ));
    Odrv4 I__4058 (
            .O(N__22657),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__4057 (
            .O(N__22652),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__4056 (
            .O(N__22649),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    InMux I__4055 (
            .O(N__22646),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    InMux I__4054 (
            .O(N__22643),
            .I(bfn_7_13_0_));
    InMux I__4053 (
            .O(N__22640),
            .I(\POWERLED.CO2 ));
    InMux I__4052 (
            .O(N__22637),
            .I(N__22634));
    LocalMux I__4051 (
            .O(N__22634),
            .I(N__22631));
    Span4Mux_v I__4050 (
            .O(N__22631),
            .I(N__22628));
    Odrv4 I__4049 (
            .O(N__22628),
            .I(\POWERLED.dutycycle_RNIZ0Z_2 ));
    InMux I__4048 (
            .O(N__22625),
            .I(N__22622));
    LocalMux I__4047 (
            .O(N__22622),
            .I(N__22618));
    InMux I__4046 (
            .O(N__22621),
            .I(N__22615));
    Span12Mux_s10_v I__4045 (
            .O(N__22618),
            .I(N__22612));
    LocalMux I__4044 (
            .O(N__22615),
            .I(N__22609));
    Odrv12 I__4043 (
            .O(N__22612),
            .I(\POWERLED.mult1_un131_sum ));
    Odrv4 I__4042 (
            .O(N__22609),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__4041 (
            .O(N__22604),
            .I(\POWERLED.un1_dutycycle_53_cry_1 ));
    InMux I__4040 (
            .O(N__22601),
            .I(N__22598));
    LocalMux I__4039 (
            .O(N__22598),
            .I(N__22595));
    Span4Mux_h I__4038 (
            .O(N__22595),
            .I(N__22592));
    Span4Mux_v I__4037 (
            .O(N__22592),
            .I(N__22589));
    Odrv4 I__4036 (
            .O(N__22589),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_2 ));
    InMux I__4035 (
            .O(N__22586),
            .I(N__22582));
    InMux I__4034 (
            .O(N__22585),
            .I(N__22579));
    LocalMux I__4033 (
            .O(N__22582),
            .I(N__22574));
    LocalMux I__4032 (
            .O(N__22579),
            .I(N__22574));
    Span12Mux_s6_h I__4031 (
            .O(N__22574),
            .I(N__22571));
    Odrv12 I__4030 (
            .O(N__22571),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__4029 (
            .O(N__22568),
            .I(\POWERLED.un1_dutycycle_53_cry_2 ));
    InMux I__4028 (
            .O(N__22565),
            .I(N__22562));
    LocalMux I__4027 (
            .O(N__22562),
            .I(N__22559));
    Span4Mux_v I__4026 (
            .O(N__22559),
            .I(N__22556));
    Odrv4 I__4025 (
            .O(N__22556),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_3 ));
    CascadeMux I__4024 (
            .O(N__22553),
            .I(N__22549));
    CascadeMux I__4023 (
            .O(N__22552),
            .I(N__22546));
    InMux I__4022 (
            .O(N__22549),
            .I(N__22543));
    InMux I__4021 (
            .O(N__22546),
            .I(N__22540));
    LocalMux I__4020 (
            .O(N__22543),
            .I(N__22537));
    LocalMux I__4019 (
            .O(N__22540),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_3 ));
    Odrv4 I__4018 (
            .O(N__22537),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_3 ));
    InMux I__4017 (
            .O(N__22532),
            .I(N__22528));
    InMux I__4016 (
            .O(N__22531),
            .I(N__22525));
    LocalMux I__4015 (
            .O(N__22528),
            .I(N__22522));
    LocalMux I__4014 (
            .O(N__22525),
            .I(N__22519));
    Span4Mux_h I__4013 (
            .O(N__22522),
            .I(N__22514));
    Span4Mux_v I__4012 (
            .O(N__22519),
            .I(N__22514));
    Odrv4 I__4011 (
            .O(N__22514),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__4010 (
            .O(N__22511),
            .I(\POWERLED.un1_dutycycle_53_cry_3 ));
    InMux I__4009 (
            .O(N__22508),
            .I(N__22504));
    InMux I__4008 (
            .O(N__22507),
            .I(N__22501));
    LocalMux I__4007 (
            .O(N__22504),
            .I(N__22498));
    LocalMux I__4006 (
            .O(N__22501),
            .I(N__22495));
    Odrv12 I__4005 (
            .O(N__22498),
            .I(\POWERLED.mult1_un110_sum ));
    Odrv4 I__4004 (
            .O(N__22495),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__4003 (
            .O(N__22490),
            .I(\POWERLED.un1_dutycycle_53_cry_4 ));
    InMux I__4002 (
            .O(N__22487),
            .I(N__22483));
    InMux I__4001 (
            .O(N__22486),
            .I(N__22480));
    LocalMux I__4000 (
            .O(N__22483),
            .I(N__22475));
    LocalMux I__3999 (
            .O(N__22480),
            .I(N__22475));
    Span4Mux_v I__3998 (
            .O(N__22475),
            .I(N__22472));
    Span4Mux_h I__3997 (
            .O(N__22472),
            .I(N__22469));
    Odrv4 I__3996 (
            .O(N__22469),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__3995 (
            .O(N__22466),
            .I(\POWERLED.un1_dutycycle_53_cry_5 ));
    InMux I__3994 (
            .O(N__22463),
            .I(N__22459));
    InMux I__3993 (
            .O(N__22462),
            .I(N__22456));
    LocalMux I__3992 (
            .O(N__22459),
            .I(N__22451));
    LocalMux I__3991 (
            .O(N__22456),
            .I(N__22451));
    Span4Mux_v I__3990 (
            .O(N__22451),
            .I(N__22448));
    Span4Mux_h I__3989 (
            .O(N__22448),
            .I(N__22445));
    Odrv4 I__3988 (
            .O(N__22445),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__3987 (
            .O(N__22442),
            .I(\POWERLED.un1_dutycycle_53_cry_6 ));
    CascadeMux I__3986 (
            .O(N__22439),
            .I(N__22436));
    InMux I__3985 (
            .O(N__22436),
            .I(N__22433));
    LocalMux I__3984 (
            .O(N__22433),
            .I(N__22430));
    Odrv4 I__3983 (
            .O(N__22430),
            .I(\POWERLED.dutycycle_RNIZ0Z_11 ));
    InMux I__3982 (
            .O(N__22427),
            .I(N__22424));
    LocalMux I__3981 (
            .O(N__22424),
            .I(N__22420));
    InMux I__3980 (
            .O(N__22423),
            .I(N__22417));
    Span4Mux_v I__3979 (
            .O(N__22420),
            .I(N__22412));
    LocalMux I__3978 (
            .O(N__22417),
            .I(N__22412));
    Odrv4 I__3977 (
            .O(N__22412),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__3976 (
            .O(N__22409),
            .I(bfn_7_12_0_));
    InMux I__3975 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__3974 (
            .O(N__22403),
            .I(N__22400));
    Odrv4 I__3973 (
            .O(N__22400),
            .I(\POWERLED.dutycycle_RNIZ0Z_12 ));
    InMux I__3972 (
            .O(N__22397),
            .I(N__22393));
    InMux I__3971 (
            .O(N__22396),
            .I(N__22390));
    LocalMux I__3970 (
            .O(N__22393),
            .I(N__22385));
    LocalMux I__3969 (
            .O(N__22390),
            .I(N__22385));
    Span4Mux_v I__3968 (
            .O(N__22385),
            .I(N__22382));
    Odrv4 I__3967 (
            .O(N__22382),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__3966 (
            .O(N__22379),
            .I(\POWERLED.un1_dutycycle_53_cry_8 ));
    CascadeMux I__3965 (
            .O(N__22376),
            .I(\POWERLED.N_9_i_1_cascade_ ));
    CascadeMux I__3964 (
            .O(N__22373),
            .I(\POWERLED.dutycycle_RNIZ0Z_8_cascade_ ));
    InMux I__3963 (
            .O(N__22370),
            .I(N__22367));
    LocalMux I__3962 (
            .O(N__22367),
            .I(N__22364));
    Span4Mux_h I__3961 (
            .O(N__22364),
            .I(N__22361));
    Odrv4 I__3960 (
            .O(N__22361),
            .I(\POWERLED.un1_clk_100khz_32_and_i_0_a2_0_0_0 ));
    CascadeMux I__3959 (
            .O(N__22358),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_6_cascade_ ));
    InMux I__3958 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__3957 (
            .O(N__22352),
            .I(\POWERLED.un2_count_clk_17_0_0_a2_0_3 ));
    InMux I__3956 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__3955 (
            .O(N__22346),
            .I(N__22342));
    InMux I__3954 (
            .O(N__22345),
            .I(N__22339));
    Span4Mux_v I__3953 (
            .O(N__22342),
            .I(N__22336));
    LocalMux I__3952 (
            .O(N__22339),
            .I(N__22333));
    Odrv4 I__3951 (
            .O(N__22336),
            .I(\POWERLED.un1_dutycycle_53_axb_0 ));
    Odrv12 I__3950 (
            .O(N__22333),
            .I(\POWERLED.un1_dutycycle_53_axb_0 ));
    CascadeMux I__3949 (
            .O(N__22328),
            .I(N__22325));
    InMux I__3948 (
            .O(N__22325),
            .I(N__22322));
    LocalMux I__3947 (
            .O(N__22322),
            .I(N__22319));
    Odrv4 I__3946 (
            .O(N__22319),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    InMux I__3945 (
            .O(N__22316),
            .I(N__22313));
    LocalMux I__3944 (
            .O(N__22313),
            .I(N__22310));
    Span4Mux_v I__3943 (
            .O(N__22310),
            .I(N__22306));
    InMux I__3942 (
            .O(N__22309),
            .I(N__22303));
    Span4Mux_h I__3941 (
            .O(N__22306),
            .I(N__22300));
    LocalMux I__3940 (
            .O(N__22303),
            .I(N__22297));
    Odrv4 I__3939 (
            .O(N__22300),
            .I(\POWERLED.mult1_un138_sum ));
    Odrv4 I__3938 (
            .O(N__22297),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__3937 (
            .O(N__22292),
            .I(\POWERLED.un1_dutycycle_53_cry_0 ));
    InMux I__3936 (
            .O(N__22289),
            .I(N__22283));
    InMux I__3935 (
            .O(N__22288),
            .I(N__22283));
    LocalMux I__3934 (
            .O(N__22283),
            .I(N__22280));
    Odrv12 I__3933 (
            .O(N__22280),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_0 ));
    CascadeMux I__3932 (
            .O(N__22277),
            .I(\POWERLED.un2_count_clk_17_0_0_a2_0_4_cascade_ ));
    InMux I__3931 (
            .O(N__22274),
            .I(N__22270));
    InMux I__3930 (
            .O(N__22273),
            .I(N__22267));
    LocalMux I__3929 (
            .O(N__22270),
            .I(\POWERLED.N_604 ));
    LocalMux I__3928 (
            .O(N__22267),
            .I(\POWERLED.N_604 ));
    InMux I__3927 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__3926 (
            .O(N__22259),
            .I(\POWERLED.func_state_RNI1O2V5Z0Z_1 ));
    CascadeMux I__3925 (
            .O(N__22256),
            .I(N__22253));
    InMux I__3924 (
            .O(N__22253),
            .I(N__22250));
    LocalMux I__3923 (
            .O(N__22250),
            .I(N__22247));
    Span4Mux_h I__3922 (
            .O(N__22247),
            .I(N__22244));
    Odrv4 I__3921 (
            .O(N__22244),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__3920 (
            .O(N__22241),
            .I(N__22237));
    CascadeMux I__3919 (
            .O(N__22240),
            .I(N__22233));
    LocalMux I__3918 (
            .O(N__22237),
            .I(N__22229));
    InMux I__3917 (
            .O(N__22236),
            .I(N__22226));
    InMux I__3916 (
            .O(N__22233),
            .I(N__22221));
    InMux I__3915 (
            .O(N__22232),
            .I(N__22221));
    Span4Mux_v I__3914 (
            .O(N__22229),
            .I(N__22218));
    LocalMux I__3913 (
            .O(N__22226),
            .I(N__22213));
    LocalMux I__3912 (
            .O(N__22221),
            .I(N__22213));
    Span4Mux_v I__3911 (
            .O(N__22218),
            .I(N__22209));
    Span4Mux_v I__3910 (
            .O(N__22213),
            .I(N__22206));
    InMux I__3909 (
            .O(N__22212),
            .I(N__22203));
    Odrv4 I__3908 (
            .O(N__22209),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    Odrv4 I__3907 (
            .O(N__22206),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__3906 (
            .O(N__22203),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__3905 (
            .O(N__22196),
            .I(N__22193));
    InMux I__3904 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__3903 (
            .O(N__22190),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__3902 (
            .O(N__22187),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    CascadeMux I__3901 (
            .O(N__22184),
            .I(N__22180));
    InMux I__3900 (
            .O(N__22183),
            .I(N__22172));
    InMux I__3899 (
            .O(N__22180),
            .I(N__22172));
    InMux I__3898 (
            .O(N__22179),
            .I(N__22172));
    LocalMux I__3897 (
            .O(N__22172),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    CascadeMux I__3896 (
            .O(N__22169),
            .I(N__22166));
    InMux I__3895 (
            .O(N__22166),
            .I(N__22163));
    LocalMux I__3894 (
            .O(N__22163),
            .I(N__22160));
    Span4Mux_v I__3893 (
            .O(N__22160),
            .I(N__22157));
    Odrv4 I__3892 (
            .O(N__22157),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__3891 (
            .O(N__22154),
            .I(N__22151));
    LocalMux I__3890 (
            .O(N__22151),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__3889 (
            .O(N__22148),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__3888 (
            .O(N__22145),
            .I(N__22142));
    LocalMux I__3887 (
            .O(N__22142),
            .I(N__22139));
    Odrv12 I__3886 (
            .O(N__22139),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__3885 (
            .O(N__22136),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    InMux I__3884 (
            .O(N__22133),
            .I(N__22130));
    LocalMux I__3883 (
            .O(N__22130),
            .I(N__22126));
    CascadeMux I__3882 (
            .O(N__22129),
            .I(N__22123));
    Span4Mux_v I__3881 (
            .O(N__22126),
            .I(N__22117));
    InMux I__3880 (
            .O(N__22123),
            .I(N__22110));
    InMux I__3879 (
            .O(N__22122),
            .I(N__22110));
    InMux I__3878 (
            .O(N__22121),
            .I(N__22110));
    InMux I__3877 (
            .O(N__22120),
            .I(N__22107));
    Odrv4 I__3876 (
            .O(N__22117),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__3875 (
            .O(N__22110),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__3874 (
            .O(N__22107),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__3873 (
            .O(N__22100),
            .I(N__22097));
    InMux I__3872 (
            .O(N__22097),
            .I(N__22094));
    LocalMux I__3871 (
            .O(N__22094),
            .I(\POWERLED.mult1_un152_sum_i ));
    InMux I__3870 (
            .O(N__22091),
            .I(N__22088));
    LocalMux I__3869 (
            .O(N__22088),
            .I(N__22085));
    Odrv12 I__3868 (
            .O(N__22085),
            .I(\POWERLED.un1_dutycycle_53_axb_4_1 ));
    InMux I__3867 (
            .O(N__22082),
            .I(N__22079));
    LocalMux I__3866 (
            .O(N__22079),
            .I(N__22076));
    Odrv4 I__3865 (
            .O(N__22076),
            .I(\POWERLED.g0_7_a2_2 ));
    CascadeMux I__3864 (
            .O(N__22073),
            .I(N__22070));
    InMux I__3863 (
            .O(N__22070),
            .I(N__22067));
    LocalMux I__3862 (
            .O(N__22067),
            .I(N__22064));
    Span4Mux_s3_v I__3861 (
            .O(N__22064),
            .I(N__22061));
    Odrv4 I__3860 (
            .O(N__22061),
            .I(\POWERLED.mult1_un145_sum_i ));
    CascadeMux I__3859 (
            .O(N__22058),
            .I(\POWERLED.N_672_cascade_ ));
    InMux I__3858 (
            .O(N__22055),
            .I(N__22049));
    InMux I__3857 (
            .O(N__22054),
            .I(N__22049));
    LocalMux I__3856 (
            .O(N__22049),
            .I(dutycycle_RNI_1_5));
    InMux I__3855 (
            .O(N__22046),
            .I(N__22043));
    LocalMux I__3854 (
            .O(N__22043),
            .I(POWERLED_un1_dutycycle_172_m1));
    CascadeMux I__3853 (
            .O(N__22040),
            .I(dutycycle_RNI_3_1_cascade_));
    InMux I__3852 (
            .O(N__22037),
            .I(N__22034));
    LocalMux I__3851 (
            .O(N__22034),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__3850 (
            .O(N__22031),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__3849 (
            .O(N__22028),
            .I(N__22025));
    LocalMux I__3848 (
            .O(N__22025),
            .I(N__22022));
    Odrv12 I__3847 (
            .O(N__22022),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    CascadeMux I__3846 (
            .O(N__22019),
            .I(N__22016));
    InMux I__3845 (
            .O(N__22016),
            .I(N__22013));
    LocalMux I__3844 (
            .O(N__22013),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__3843 (
            .O(N__22010),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    CascadeMux I__3842 (
            .O(N__22007),
            .I(N__22004));
    InMux I__3841 (
            .O(N__22004),
            .I(N__22001));
    LocalMux I__3840 (
            .O(N__22001),
            .I(N__21998));
    Span4Mux_v I__3839 (
            .O(N__21998),
            .I(N__21995));
    Odrv4 I__3838 (
            .O(N__21995),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__3837 (
            .O(N__21992),
            .I(N__21989));
    LocalMux I__3836 (
            .O(N__21989),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__3835 (
            .O(N__21986),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__3834 (
            .O(N__21983),
            .I(N__21980));
    LocalMux I__3833 (
            .O(N__21980),
            .I(N__21977));
    Odrv12 I__3832 (
            .O(N__21977),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    CascadeMux I__3831 (
            .O(N__21974),
            .I(\POWERLED.dutycycle_cascade_ ));
    CascadeMux I__3830 (
            .O(N__21971),
            .I(N__21968));
    InMux I__3829 (
            .O(N__21968),
            .I(N__21965));
    LocalMux I__3828 (
            .O(N__21965),
            .I(\POWERLED.dutycycle_1_0_0 ));
    CascadeMux I__3827 (
            .O(N__21962),
            .I(\POWERLED.dutycycle_1_0_0_cascade_ ));
    InMux I__3826 (
            .O(N__21959),
            .I(N__21953));
    InMux I__3825 (
            .O(N__21958),
            .I(N__21953));
    LocalMux I__3824 (
            .O(N__21953),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    CascadeMux I__3823 (
            .O(N__21950),
            .I(\POWERLED.dutycycle_1_0_1_cascade_ ));
    CascadeMux I__3822 (
            .O(N__21947),
            .I(dutycycle_RNII6848_0_1_cascade_));
    InMux I__3821 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__3820 (
            .O(N__21941),
            .I(\POWERLED.dutycycle_eena_0 ));
    InMux I__3819 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__3818 (
            .O(N__21935),
            .I(\POWERLED.dutycycle_1_0_1 ));
    CascadeMux I__3817 (
            .O(N__21932),
            .I(\POWERLED.dutycycle_eena_0_cascade_ ));
    InMux I__3816 (
            .O(N__21929),
            .I(N__21923));
    InMux I__3815 (
            .O(N__21928),
            .I(N__21923));
    LocalMux I__3814 (
            .O(N__21923),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    CascadeMux I__3813 (
            .O(N__21920),
            .I(N__21917));
    InMux I__3812 (
            .O(N__21917),
            .I(N__21914));
    LocalMux I__3811 (
            .O(N__21914),
            .I(N__21911));
    Span12Mux_s6_h I__3810 (
            .O(N__21911),
            .I(N__21908));
    Odrv12 I__3809 (
            .O(N__21908),
            .I(\POWERLED.N_15 ));
    CascadeMux I__3808 (
            .O(N__21905),
            .I(\POWERLED.un1_dutycycle_172_m1_ns_1_cascade_ ));
    InMux I__3807 (
            .O(N__21902),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__3806 (
            .O(N__21899),
            .I(N__21896));
    InMux I__3805 (
            .O(N__21896),
            .I(N__21887));
    InMux I__3804 (
            .O(N__21895),
            .I(N__21887));
    InMux I__3803 (
            .O(N__21894),
            .I(N__21887));
    LocalMux I__3802 (
            .O(N__21887),
            .I(N__21884));
    Span12Mux_s7_v I__3801 (
            .O(N__21884),
            .I(N__21879));
    InMux I__3800 (
            .O(N__21883),
            .I(N__21876));
    InMux I__3799 (
            .O(N__21882),
            .I(N__21873));
    Odrv12 I__3798 (
            .O(N__21879),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3797 (
            .O(N__21876),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3796 (
            .O(N__21873),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    CascadeMux I__3795 (
            .O(N__21866),
            .I(N__21862));
    InMux I__3794 (
            .O(N__21865),
            .I(N__21854));
    InMux I__3793 (
            .O(N__21862),
            .I(N__21854));
    InMux I__3792 (
            .O(N__21861),
            .I(N__21854));
    LocalMux I__3791 (
            .O(N__21854),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    InMux I__3790 (
            .O(N__21851),
            .I(N__21845));
    InMux I__3789 (
            .O(N__21850),
            .I(N__21845));
    LocalMux I__3788 (
            .O(N__21845),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    CascadeMux I__3787 (
            .O(N__21842),
            .I(\POWERLED.dutycycleZ0Z_0_cascade_ ));
    CascadeMux I__3786 (
            .O(N__21839),
            .I(\POWERLED.un1_dutycycle_53_axb_3_1_cascade_ ));
    CascadeMux I__3785 (
            .O(N__21836),
            .I(\POWERLED.un1_dutycycle_53_axb_3_cascade_ ));
    InMux I__3784 (
            .O(N__21833),
            .I(N__21830));
    LocalMux I__3783 (
            .O(N__21830),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10 ));
    CascadeMux I__3782 (
            .O(N__21827),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12_cascade_ ));
    InMux I__3781 (
            .O(N__21824),
            .I(N__21821));
    LocalMux I__3780 (
            .O(N__21821),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9 ));
    InMux I__3779 (
            .O(N__21818),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    InMux I__3778 (
            .O(N__21815),
            .I(N__21812));
    LocalMux I__3777 (
            .O(N__21812),
            .I(N__21809));
    Span4Mux_s3_v I__3776 (
            .O(N__21809),
            .I(N__21806));
    Span4Mux_v I__3775 (
            .O(N__21806),
            .I(N__21803));
    Odrv4 I__3774 (
            .O(N__21803),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__3773 (
            .O(N__21800),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    CascadeMux I__3772 (
            .O(N__21797),
            .I(N__21794));
    InMux I__3771 (
            .O(N__21794),
            .I(N__21791));
    LocalMux I__3770 (
            .O(N__21791),
            .I(N__21788));
    Span4Mux_s3_v I__3769 (
            .O(N__21788),
            .I(N__21785));
    Span4Mux_v I__3768 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__3767 (
            .O(N__21782),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__3766 (
            .O(N__21779),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__3765 (
            .O(N__21776),
            .I(N__21773));
    LocalMux I__3764 (
            .O(N__21773),
            .I(N__21770));
    Span4Mux_s3_v I__3763 (
            .O(N__21770),
            .I(N__21767));
    Span4Mux_v I__3762 (
            .O(N__21767),
            .I(N__21764));
    Odrv4 I__3761 (
            .O(N__21764),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__3760 (
            .O(N__21761),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    CascadeMux I__3759 (
            .O(N__21758),
            .I(N__21755));
    InMux I__3758 (
            .O(N__21755),
            .I(N__21752));
    LocalMux I__3757 (
            .O(N__21752),
            .I(N__21749));
    Span4Mux_s3_v I__3756 (
            .O(N__21749),
            .I(N__21746));
    Span4Mux_v I__3755 (
            .O(N__21746),
            .I(N__21743));
    Odrv4 I__3754 (
            .O(N__21743),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    InMux I__3753 (
            .O(N__21740),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__3752 (
            .O(N__21737),
            .I(N__21734));
    LocalMux I__3751 (
            .O(N__21734),
            .I(N__21731));
    Span4Mux_h I__3750 (
            .O(N__21731),
            .I(N__21728));
    Span4Mux_v I__3749 (
            .O(N__21728),
            .I(N__21725));
    Odrv4 I__3748 (
            .O(N__21725),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    CascadeMux I__3747 (
            .O(N__21722),
            .I(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1_cascade_ ));
    CascadeMux I__3746 (
            .O(N__21719),
            .I(N__21699));
    CascadeMux I__3745 (
            .O(N__21718),
            .I(N__21695));
    InMux I__3744 (
            .O(N__21717),
            .I(N__21682));
    InMux I__3743 (
            .O(N__21716),
            .I(N__21682));
    InMux I__3742 (
            .O(N__21715),
            .I(N__21682));
    InMux I__3741 (
            .O(N__21714),
            .I(N__21682));
    InMux I__3740 (
            .O(N__21713),
            .I(N__21682));
    InMux I__3739 (
            .O(N__21712),
            .I(N__21673));
    InMux I__3738 (
            .O(N__21711),
            .I(N__21673));
    InMux I__3737 (
            .O(N__21710),
            .I(N__21673));
    InMux I__3736 (
            .O(N__21709),
            .I(N__21673));
    InMux I__3735 (
            .O(N__21708),
            .I(N__21670));
    InMux I__3734 (
            .O(N__21707),
            .I(N__21661));
    InMux I__3733 (
            .O(N__21706),
            .I(N__21661));
    InMux I__3732 (
            .O(N__21705),
            .I(N__21661));
    InMux I__3731 (
            .O(N__21704),
            .I(N__21661));
    InMux I__3730 (
            .O(N__21703),
            .I(N__21652));
    InMux I__3729 (
            .O(N__21702),
            .I(N__21652));
    InMux I__3728 (
            .O(N__21699),
            .I(N__21652));
    InMux I__3727 (
            .O(N__21698),
            .I(N__21652));
    InMux I__3726 (
            .O(N__21695),
            .I(N__21649));
    CascadeMux I__3725 (
            .O(N__21694),
            .I(N__21640));
    CascadeMux I__3724 (
            .O(N__21693),
            .I(N__21637));
    LocalMux I__3723 (
            .O(N__21682),
            .I(N__21629));
    LocalMux I__3722 (
            .O(N__21673),
            .I(N__21624));
    LocalMux I__3721 (
            .O(N__21670),
            .I(N__21624));
    LocalMux I__3720 (
            .O(N__21661),
            .I(N__21621));
    LocalMux I__3719 (
            .O(N__21652),
            .I(N__21616));
    LocalMux I__3718 (
            .O(N__21649),
            .I(N__21616));
    InMux I__3717 (
            .O(N__21648),
            .I(N__21613));
    InMux I__3716 (
            .O(N__21647),
            .I(N__21610));
    InMux I__3715 (
            .O(N__21646),
            .I(N__21607));
    InMux I__3714 (
            .O(N__21645),
            .I(N__21604));
    InMux I__3713 (
            .O(N__21644),
            .I(N__21593));
    InMux I__3712 (
            .O(N__21643),
            .I(N__21593));
    InMux I__3711 (
            .O(N__21640),
            .I(N__21593));
    InMux I__3710 (
            .O(N__21637),
            .I(N__21593));
    InMux I__3709 (
            .O(N__21636),
            .I(N__21593));
    InMux I__3708 (
            .O(N__21635),
            .I(N__21584));
    InMux I__3707 (
            .O(N__21634),
            .I(N__21584));
    InMux I__3706 (
            .O(N__21633),
            .I(N__21584));
    InMux I__3705 (
            .O(N__21632),
            .I(N__21584));
    Span4Mux_s1_v I__3704 (
            .O(N__21629),
            .I(N__21577));
    Span4Mux_v I__3703 (
            .O(N__21624),
            .I(N__21577));
    Span4Mux_v I__3702 (
            .O(N__21621),
            .I(N__21577));
    Span4Mux_h I__3701 (
            .O(N__21616),
            .I(N__21574));
    LocalMux I__3700 (
            .O(N__21613),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__3699 (
            .O(N__21610),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__3698 (
            .O(N__21607),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__3697 (
            .O(N__21604),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__3696 (
            .O(N__21593),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__3695 (
            .O(N__21584),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__3694 (
            .O(N__21577),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__3693 (
            .O(N__21574),
            .I(\VPP_VDDQ.N_1_i ));
    CascadeMux I__3692 (
            .O(N__21557),
            .I(\VPP_VDDQ.N_664_cascade_ ));
    CascadeMux I__3691 (
            .O(N__21554),
            .I(\VPP_VDDQ.m4_0_0_cascade_ ));
    InMux I__3690 (
            .O(N__21551),
            .I(N__21533));
    InMux I__3689 (
            .O(N__21550),
            .I(N__21524));
    InMux I__3688 (
            .O(N__21549),
            .I(N__21524));
    InMux I__3687 (
            .O(N__21548),
            .I(N__21524));
    InMux I__3686 (
            .O(N__21547),
            .I(N__21524));
    CascadeMux I__3685 (
            .O(N__21546),
            .I(N__21519));
    InMux I__3684 (
            .O(N__21545),
            .I(N__21513));
    InMux I__3683 (
            .O(N__21544),
            .I(N__21504));
    InMux I__3682 (
            .O(N__21543),
            .I(N__21504));
    InMux I__3681 (
            .O(N__21542),
            .I(N__21504));
    InMux I__3680 (
            .O(N__21541),
            .I(N__21504));
    InMux I__3679 (
            .O(N__21540),
            .I(N__21497));
    InMux I__3678 (
            .O(N__21539),
            .I(N__21497));
    InMux I__3677 (
            .O(N__21538),
            .I(N__21497));
    InMux I__3676 (
            .O(N__21537),
            .I(N__21492));
    InMux I__3675 (
            .O(N__21536),
            .I(N__21492));
    LocalMux I__3674 (
            .O(N__21533),
            .I(N__21475));
    LocalMux I__3673 (
            .O(N__21524),
            .I(N__21475));
    InMux I__3672 (
            .O(N__21523),
            .I(N__21466));
    InMux I__3671 (
            .O(N__21522),
            .I(N__21466));
    InMux I__3670 (
            .O(N__21519),
            .I(N__21466));
    InMux I__3669 (
            .O(N__21518),
            .I(N__21466));
    InMux I__3668 (
            .O(N__21517),
            .I(N__21461));
    InMux I__3667 (
            .O(N__21516),
            .I(N__21461));
    LocalMux I__3666 (
            .O(N__21513),
            .I(N__21456));
    LocalMux I__3665 (
            .O(N__21504),
            .I(N__21456));
    LocalMux I__3664 (
            .O(N__21497),
            .I(N__21451));
    LocalMux I__3663 (
            .O(N__21492),
            .I(N__21451));
    InMux I__3662 (
            .O(N__21491),
            .I(N__21440));
    InMux I__3661 (
            .O(N__21490),
            .I(N__21440));
    InMux I__3660 (
            .O(N__21489),
            .I(N__21440));
    InMux I__3659 (
            .O(N__21488),
            .I(N__21440));
    InMux I__3658 (
            .O(N__21487),
            .I(N__21440));
    InMux I__3657 (
            .O(N__21486),
            .I(N__21429));
    InMux I__3656 (
            .O(N__21485),
            .I(N__21429));
    InMux I__3655 (
            .O(N__21484),
            .I(N__21429));
    InMux I__3654 (
            .O(N__21483),
            .I(N__21429));
    InMux I__3653 (
            .O(N__21482),
            .I(N__21429));
    InMux I__3652 (
            .O(N__21481),
            .I(N__21422));
    InMux I__3651 (
            .O(N__21480),
            .I(N__21419));
    Span4Mux_h I__3650 (
            .O(N__21475),
            .I(N__21414));
    LocalMux I__3649 (
            .O(N__21466),
            .I(N__21414));
    LocalMux I__3648 (
            .O(N__21461),
            .I(N__21409));
    Span4Mux_h I__3647 (
            .O(N__21456),
            .I(N__21409));
    Span4Mux_v I__3646 (
            .O(N__21451),
            .I(N__21402));
    LocalMux I__3645 (
            .O(N__21440),
            .I(N__21402));
    LocalMux I__3644 (
            .O(N__21429),
            .I(N__21402));
    InMux I__3643 (
            .O(N__21428),
            .I(N__21397));
    InMux I__3642 (
            .O(N__21427),
            .I(N__21397));
    InMux I__3641 (
            .O(N__21426),
            .I(N__21394));
    InMux I__3640 (
            .O(N__21425),
            .I(N__21391));
    LocalMux I__3639 (
            .O(N__21422),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__3638 (
            .O(N__21419),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__3637 (
            .O(N__21414),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__3636 (
            .O(N__21409),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__3635 (
            .O(N__21402),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__3634 (
            .O(N__21397),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__3633 (
            .O(N__21394),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__3632 (
            .O(N__21391),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    InMux I__3631 (
            .O(N__21374),
            .I(N__21364));
    InMux I__3630 (
            .O(N__21373),
            .I(N__21364));
    InMux I__3629 (
            .O(N__21372),
            .I(N__21364));
    InMux I__3628 (
            .O(N__21371),
            .I(N__21361));
    LocalMux I__3627 (
            .O(N__21364),
            .I(N__21358));
    LocalMux I__3626 (
            .O(N__21361),
            .I(N__21355));
    Odrv4 I__3625 (
            .O(N__21358),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ));
    Odrv4 I__3624 (
            .O(N__21355),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ));
    CascadeMux I__3623 (
            .O(N__21350),
            .I(N__21345));
    CascadeMux I__3622 (
            .O(N__21349),
            .I(N__21341));
    CascadeMux I__3621 (
            .O(N__21348),
            .I(N__21338));
    InMux I__3620 (
            .O(N__21345),
            .I(N__21329));
    InMux I__3619 (
            .O(N__21344),
            .I(N__21329));
    InMux I__3618 (
            .O(N__21341),
            .I(N__21329));
    InMux I__3617 (
            .O(N__21338),
            .I(N__21322));
    InMux I__3616 (
            .O(N__21337),
            .I(N__21322));
    InMux I__3615 (
            .O(N__21336),
            .I(N__21322));
    LocalMux I__3614 (
            .O(N__21329),
            .I(N__21317));
    LocalMux I__3613 (
            .O(N__21322),
            .I(N__21317));
    Span4Mux_s1_v I__3612 (
            .O(N__21317),
            .I(N__21314));
    Span4Mux_v I__3611 (
            .O(N__21314),
            .I(N__21310));
    InMux I__3610 (
            .O(N__21313),
            .I(N__21307));
    Span4Mux_h I__3609 (
            .O(N__21310),
            .I(N__21301));
    LocalMux I__3608 (
            .O(N__21307),
            .I(N__21301));
    InMux I__3607 (
            .O(N__21306),
            .I(N__21298));
    Span4Mux_v I__3606 (
            .O(N__21301),
            .I(N__21295));
    LocalMux I__3605 (
            .O(N__21298),
            .I(N__21292));
    Span4Mux_v I__3604 (
            .O(N__21295),
            .I(N__21289));
    Span12Mux_v I__3603 (
            .O(N__21292),
            .I(N__21286));
    Sp12to4 I__3602 (
            .O(N__21289),
            .I(N__21283));
    Odrv12 I__3601 (
            .O(N__21286),
            .I(vddq_ok));
    Odrv12 I__3600 (
            .O(N__21283),
            .I(vddq_ok));
    CascadeMux I__3599 (
            .O(N__21278),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    InMux I__3598 (
            .O(N__21275),
            .I(N__21269));
    InMux I__3597 (
            .O(N__21274),
            .I(N__21269));
    LocalMux I__3596 (
            .O(N__21269),
            .I(\VPP_VDDQ.N_664 ));
    InMux I__3595 (
            .O(N__21266),
            .I(N__21263));
    LocalMux I__3594 (
            .O(N__21263),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    InMux I__3593 (
            .O(N__21260),
            .I(N__21257));
    LocalMux I__3592 (
            .O(N__21257),
            .I(\VPP_VDDQ.N_53 ));
    InMux I__3591 (
            .O(N__21254),
            .I(N__21251));
    LocalMux I__3590 (
            .O(N__21251),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    CascadeMux I__3589 (
            .O(N__21248),
            .I(N__21242));
    CascadeMux I__3588 (
            .O(N__21247),
            .I(N__21239));
    InMux I__3587 (
            .O(N__21246),
            .I(N__21234));
    InMux I__3586 (
            .O(N__21245),
            .I(N__21231));
    InMux I__3585 (
            .O(N__21242),
            .I(N__21228));
    InMux I__3584 (
            .O(N__21239),
            .I(N__21225));
    InMux I__3583 (
            .O(N__21238),
            .I(N__21222));
    InMux I__3582 (
            .O(N__21237),
            .I(N__21219));
    LocalMux I__3581 (
            .O(N__21234),
            .I(N__21216));
    LocalMux I__3580 (
            .O(N__21231),
            .I(N__21203));
    LocalMux I__3579 (
            .O(N__21228),
            .I(N__21200));
    LocalMux I__3578 (
            .O(N__21225),
            .I(N__21196));
    LocalMux I__3577 (
            .O(N__21222),
            .I(N__21193));
    LocalMux I__3576 (
            .O(N__21219),
            .I(N__21190));
    Glb2LocalMux I__3575 (
            .O(N__21216),
            .I(N__21155));
    CEMux I__3574 (
            .O(N__21215),
            .I(N__21155));
    CEMux I__3573 (
            .O(N__21214),
            .I(N__21155));
    CEMux I__3572 (
            .O(N__21213),
            .I(N__21155));
    CEMux I__3571 (
            .O(N__21212),
            .I(N__21155));
    CEMux I__3570 (
            .O(N__21211),
            .I(N__21155));
    CEMux I__3569 (
            .O(N__21210),
            .I(N__21155));
    CEMux I__3568 (
            .O(N__21209),
            .I(N__21155));
    CEMux I__3567 (
            .O(N__21208),
            .I(N__21155));
    CEMux I__3566 (
            .O(N__21207),
            .I(N__21155));
    CEMux I__3565 (
            .O(N__21206),
            .I(N__21155));
    Glb2LocalMux I__3564 (
            .O(N__21203),
            .I(N__21155));
    Glb2LocalMux I__3563 (
            .O(N__21200),
            .I(N__21155));
    CEMux I__3562 (
            .O(N__21199),
            .I(N__21155));
    Glb2LocalMux I__3561 (
            .O(N__21196),
            .I(N__21155));
    Glb2LocalMux I__3560 (
            .O(N__21193),
            .I(N__21155));
    Glb2LocalMux I__3559 (
            .O(N__21190),
            .I(N__21155));
    GlobalMux I__3558 (
            .O(N__21155),
            .I(N__21152));
    gio2CtrlBuf I__3557 (
            .O(N__21152),
            .I(N_557_g));
    CascadeMux I__3556 (
            .O(N__21149),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_ ));
    CascadeMux I__3555 (
            .O(N__21146),
            .I(N__21143));
    InMux I__3554 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__3553 (
            .O(N__21140),
            .I(N__21137));
    Odrv4 I__3552 (
            .O(N__21137),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__3551 (
            .O(N__21134),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    CascadeMux I__3550 (
            .O(N__21131),
            .I(N__21128));
    InMux I__3549 (
            .O(N__21128),
            .I(N__21125));
    LocalMux I__3548 (
            .O(N__21125),
            .I(N__21122));
    Odrv4 I__3547 (
            .O(N__21122),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__3546 (
            .O(N__21119),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__3545 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__3544 (
            .O(N__21113),
            .I(N__21110));
    Odrv4 I__3543 (
            .O(N__21110),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__3542 (
            .O(N__21107),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__3541 (
            .O(N__21104),
            .I(N__21101));
    LocalMux I__3540 (
            .O(N__21101),
            .I(N__21098));
    Odrv4 I__3539 (
            .O(N__21098),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    InMux I__3538 (
            .O(N__21095),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__3537 (
            .O(N__21092),
            .I(N__21089));
    LocalMux I__3536 (
            .O(N__21089),
            .I(N__21086));
    Odrv4 I__3535 (
            .O(N__21086),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__3534 (
            .O(N__21083),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__3533 (
            .O(N__21080),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    CascadeMux I__3532 (
            .O(N__21077),
            .I(N__21074));
    InMux I__3531 (
            .O(N__21074),
            .I(N__21071));
    LocalMux I__3530 (
            .O(N__21071),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    CascadeMux I__3529 (
            .O(N__21068),
            .I(\VPP_VDDQ.N_53_cascade_ ));
    CascadeMux I__3528 (
            .O(N__21065),
            .I(N__21044));
    CascadeMux I__3527 (
            .O(N__21064),
            .I(N__21041));
    CascadeMux I__3526 (
            .O(N__21063),
            .I(N__21038));
    CascadeMux I__3525 (
            .O(N__21062),
            .I(N__21035));
    CascadeMux I__3524 (
            .O(N__21061),
            .I(N__21032));
    CascadeMux I__3523 (
            .O(N__21060),
            .I(N__21029));
    CascadeMux I__3522 (
            .O(N__21059),
            .I(N__21025));
    CascadeMux I__3521 (
            .O(N__21058),
            .I(N__21022));
    InMux I__3520 (
            .O(N__21057),
            .I(N__21019));
    CascadeMux I__3519 (
            .O(N__21056),
            .I(N__21016));
    CascadeMux I__3518 (
            .O(N__21055),
            .I(N__21012));
    CascadeMux I__3517 (
            .O(N__21054),
            .I(N__21009));
    CascadeMux I__3516 (
            .O(N__21053),
            .I(N__21005));
    CascadeMux I__3515 (
            .O(N__21052),
            .I(N__21001));
    CascadeMux I__3514 (
            .O(N__21051),
            .I(N__20994));
    CascadeMux I__3513 (
            .O(N__21050),
            .I(N__20991));
    CascadeMux I__3512 (
            .O(N__21049),
            .I(N__20988));
    CascadeMux I__3511 (
            .O(N__21048),
            .I(N__20983));
    InMux I__3510 (
            .O(N__21047),
            .I(N__20970));
    InMux I__3509 (
            .O(N__21044),
            .I(N__20970));
    InMux I__3508 (
            .O(N__21041),
            .I(N__20970));
    InMux I__3507 (
            .O(N__21038),
            .I(N__20970));
    InMux I__3506 (
            .O(N__21035),
            .I(N__20970));
    InMux I__3505 (
            .O(N__21032),
            .I(N__20961));
    InMux I__3504 (
            .O(N__21029),
            .I(N__20961));
    InMux I__3503 (
            .O(N__21028),
            .I(N__20961));
    InMux I__3502 (
            .O(N__21025),
            .I(N__20961));
    InMux I__3501 (
            .O(N__21022),
            .I(N__20958));
    LocalMux I__3500 (
            .O(N__21019),
            .I(N__20954));
    InMux I__3499 (
            .O(N__21016),
            .I(N__20947));
    InMux I__3498 (
            .O(N__21015),
            .I(N__20947));
    InMux I__3497 (
            .O(N__21012),
            .I(N__20947));
    InMux I__3496 (
            .O(N__21009),
            .I(N__20936));
    InMux I__3495 (
            .O(N__21008),
            .I(N__20936));
    InMux I__3494 (
            .O(N__21005),
            .I(N__20936));
    InMux I__3493 (
            .O(N__21004),
            .I(N__20936));
    InMux I__3492 (
            .O(N__21001),
            .I(N__20936));
    InMux I__3491 (
            .O(N__21000),
            .I(N__20927));
    InMux I__3490 (
            .O(N__20999),
            .I(N__20927));
    InMux I__3489 (
            .O(N__20998),
            .I(N__20927));
    InMux I__3488 (
            .O(N__20997),
            .I(N__20927));
    InMux I__3487 (
            .O(N__20994),
            .I(N__20924));
    InMux I__3486 (
            .O(N__20991),
            .I(N__20915));
    InMux I__3485 (
            .O(N__20988),
            .I(N__20915));
    InMux I__3484 (
            .O(N__20987),
            .I(N__20915));
    InMux I__3483 (
            .O(N__20986),
            .I(N__20915));
    InMux I__3482 (
            .O(N__20983),
            .I(N__20912));
    InMux I__3481 (
            .O(N__20982),
            .I(N__20909));
    CascadeMux I__3480 (
            .O(N__20981),
            .I(N__20906));
    LocalMux I__3479 (
            .O(N__20970),
            .I(N__20899));
    LocalMux I__3478 (
            .O(N__20961),
            .I(N__20899));
    LocalMux I__3477 (
            .O(N__20958),
            .I(N__20899));
    CascadeMux I__3476 (
            .O(N__20957),
            .I(N__20896));
    Span4Mux_h I__3475 (
            .O(N__20954),
            .I(N__20890));
    LocalMux I__3474 (
            .O(N__20947),
            .I(N__20890));
    LocalMux I__3473 (
            .O(N__20936),
            .I(N__20885));
    LocalMux I__3472 (
            .O(N__20927),
            .I(N__20885));
    LocalMux I__3471 (
            .O(N__20924),
            .I(N__20876));
    LocalMux I__3470 (
            .O(N__20915),
            .I(N__20876));
    LocalMux I__3469 (
            .O(N__20912),
            .I(N__20876));
    LocalMux I__3468 (
            .O(N__20909),
            .I(N__20876));
    InMux I__3467 (
            .O(N__20906),
            .I(N__20873));
    Span4Mux_v I__3466 (
            .O(N__20899),
            .I(N__20870));
    InMux I__3465 (
            .O(N__20896),
            .I(N__20865));
    InMux I__3464 (
            .O(N__20895),
            .I(N__20865));
    Span4Mux_v I__3463 (
            .O(N__20890),
            .I(N__20858));
    Span4Mux_h I__3462 (
            .O(N__20885),
            .I(N__20858));
    Span4Mux_v I__3461 (
            .O(N__20876),
            .I(N__20858));
    LocalMux I__3460 (
            .O(N__20873),
            .I(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1 ));
    Odrv4 I__3459 (
            .O(N__20870),
            .I(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1 ));
    LocalMux I__3458 (
            .O(N__20865),
            .I(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1 ));
    Odrv4 I__3457 (
            .O(N__20858),
            .I(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1 ));
    InMux I__3456 (
            .O(N__20849),
            .I(N__20846));
    LocalMux I__3455 (
            .O(N__20846),
            .I(\POWERLED.un79_clk_100khzlto15_3 ));
    InMux I__3454 (
            .O(N__20843),
            .I(N__20838));
    InMux I__3453 (
            .O(N__20842),
            .I(N__20835));
    InMux I__3452 (
            .O(N__20841),
            .I(N__20832));
    LocalMux I__3451 (
            .O(N__20838),
            .I(N__20829));
    LocalMux I__3450 (
            .O(N__20835),
            .I(N__20824));
    LocalMux I__3449 (
            .O(N__20832),
            .I(N__20824));
    Span4Mux_v I__3448 (
            .O(N__20829),
            .I(N__20820));
    Span4Mux_v I__3447 (
            .O(N__20824),
            .I(N__20817));
    InMux I__3446 (
            .O(N__20823),
            .I(N__20814));
    Odrv4 I__3445 (
            .O(N__20820),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv4 I__3444 (
            .O(N__20817),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__3443 (
            .O(N__20814),
            .I(\POWERLED.countZ0Z_15 ));
    InMux I__3442 (
            .O(N__20807),
            .I(N__20803));
    InMux I__3441 (
            .O(N__20806),
            .I(N__20799));
    LocalMux I__3440 (
            .O(N__20803),
            .I(N__20796));
    CascadeMux I__3439 (
            .O(N__20802),
            .I(N__20793));
    LocalMux I__3438 (
            .O(N__20799),
            .I(N__20790));
    Span4Mux_v I__3437 (
            .O(N__20796),
            .I(N__20787));
    InMux I__3436 (
            .O(N__20793),
            .I(N__20784));
    Odrv12 I__3435 (
            .O(N__20790),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__3434 (
            .O(N__20787),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__3433 (
            .O(N__20784),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__3432 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__3431 (
            .O(N__20774),
            .I(N__20771));
    Span4Mux_s3_v I__3430 (
            .O(N__20771),
            .I(N__20768));
    Span4Mux_h I__3429 (
            .O(N__20768),
            .I(N__20765));
    Odrv4 I__3428 (
            .O(N__20765),
            .I(\POWERLED.g1_i_o4_5 ));
    InMux I__3427 (
            .O(N__20762),
            .I(N__20759));
    LocalMux I__3426 (
            .O(N__20759),
            .I(N__20756));
    Span4Mux_v I__3425 (
            .O(N__20756),
            .I(N__20751));
    CascadeMux I__3424 (
            .O(N__20755),
            .I(N__20748));
    CascadeMux I__3423 (
            .O(N__20754),
            .I(N__20744));
    Span4Mux_v I__3422 (
            .O(N__20751),
            .I(N__20741));
    InMux I__3421 (
            .O(N__20748),
            .I(N__20736));
    InMux I__3420 (
            .O(N__20747),
            .I(N__20736));
    InMux I__3419 (
            .O(N__20744),
            .I(N__20733));
    Odrv4 I__3418 (
            .O(N__20741),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__3417 (
            .O(N__20736),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__3416 (
            .O(N__20733),
            .I(\POWERLED.countZ0Z_7 ));
    InMux I__3415 (
            .O(N__20726),
            .I(N__20720));
    InMux I__3414 (
            .O(N__20725),
            .I(N__20720));
    LocalMux I__3413 (
            .O(N__20720),
            .I(\POWERLED.count_1_7 ));
    InMux I__3412 (
            .O(N__20717),
            .I(N__20714));
    LocalMux I__3411 (
            .O(N__20714),
            .I(N__20711));
    Odrv4 I__3410 (
            .O(N__20711),
            .I(\POWERLED.count_0_7 ));
    InMux I__3409 (
            .O(N__20708),
            .I(N__20705));
    LocalMux I__3408 (
            .O(N__20705),
            .I(N__20702));
    Odrv12 I__3407 (
            .O(N__20702),
            .I(\POWERLED.N_6 ));
    InMux I__3406 (
            .O(N__20699),
            .I(N__20696));
    LocalMux I__3405 (
            .O(N__20696),
            .I(N__20693));
    Span4Mux_v I__3404 (
            .O(N__20693),
            .I(N__20690));
    Odrv4 I__3403 (
            .O(N__20690),
            .I(\POWERLED.count_clk_0_6 ));
    InMux I__3402 (
            .O(N__20687),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__3401 (
            .O(N__20684),
            .I(N__20681));
    InMux I__3400 (
            .O(N__20681),
            .I(N__20677));
    CascadeMux I__3399 (
            .O(N__20680),
            .I(N__20673));
    LocalMux I__3398 (
            .O(N__20677),
            .I(N__20669));
    InMux I__3397 (
            .O(N__20676),
            .I(N__20664));
    InMux I__3396 (
            .O(N__20673),
            .I(N__20664));
    InMux I__3395 (
            .O(N__20672),
            .I(N__20661));
    Odrv4 I__3394 (
            .O(N__20669),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__3393 (
            .O(N__20664),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__3392 (
            .O(N__20661),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__3391 (
            .O(N__20654),
            .I(\POWERLED.mult1_un61_sum_s_8_cascade_ ));
    CascadeMux I__3390 (
            .O(N__20651),
            .I(N__20647));
    CascadeMux I__3389 (
            .O(N__20650),
            .I(N__20643));
    InMux I__3388 (
            .O(N__20647),
            .I(N__20636));
    InMux I__3387 (
            .O(N__20646),
            .I(N__20636));
    InMux I__3386 (
            .O(N__20643),
            .I(N__20636));
    LocalMux I__3385 (
            .O(N__20636),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__3384 (
            .O(N__20633),
            .I(N__20630));
    LocalMux I__3383 (
            .O(N__20630),
            .I(N__20626));
    CascadeMux I__3382 (
            .O(N__20629),
            .I(N__20623));
    Span4Mux_v I__3381 (
            .O(N__20626),
            .I(N__20620));
    InMux I__3380 (
            .O(N__20623),
            .I(N__20617));
    Odrv4 I__3379 (
            .O(N__20620),
            .I(\POWERLED.mult1_un82_sum_i_8 ));
    LocalMux I__3378 (
            .O(N__20617),
            .I(\POWERLED.mult1_un82_sum_i_8 ));
    InMux I__3377 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__3376 (
            .O(N__20609),
            .I(N__20606));
    Span4Mux_h I__3375 (
            .O(N__20606),
            .I(N__20603));
    Odrv4 I__3374 (
            .O(N__20603),
            .I(\POWERLED.count_RNICOIT_0Z0Z_12 ));
    InMux I__3373 (
            .O(N__20600),
            .I(N__20597));
    LocalMux I__3372 (
            .O(N__20597),
            .I(\POWERLED.count_0_13 ));
    CascadeMux I__3371 (
            .O(N__20594),
            .I(N__20591));
    InMux I__3370 (
            .O(N__20591),
            .I(N__20585));
    InMux I__3369 (
            .O(N__20590),
            .I(N__20585));
    LocalMux I__3368 (
            .O(N__20585),
            .I(\POWERLED.count_1_13 ));
    InMux I__3367 (
            .O(N__20582),
            .I(N__20579));
    LocalMux I__3366 (
            .O(N__20579),
            .I(N__20575));
    CascadeMux I__3365 (
            .O(N__20578),
            .I(N__20572));
    Span4Mux_v I__3364 (
            .O(N__20575),
            .I(N__20569));
    InMux I__3363 (
            .O(N__20572),
            .I(N__20566));
    Odrv4 I__3362 (
            .O(N__20569),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__3361 (
            .O(N__20566),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__3360 (
            .O(N__20561),
            .I(N__20554));
    InMux I__3359 (
            .O(N__20560),
            .I(N__20554));
    InMux I__3358 (
            .O(N__20559),
            .I(N__20551));
    LocalMux I__3357 (
            .O(N__20554),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__3356 (
            .O(N__20551),
            .I(\POWERLED.countZ0Z_12 ));
    CascadeMux I__3355 (
            .O(N__20546),
            .I(\POWERLED.countZ0Z_13_cascade_ ));
    CascadeMux I__3354 (
            .O(N__20543),
            .I(N__20539));
    CascadeMux I__3353 (
            .O(N__20542),
            .I(N__20536));
    InMux I__3352 (
            .O(N__20539),
            .I(N__20527));
    InMux I__3351 (
            .O(N__20536),
            .I(N__20527));
    InMux I__3350 (
            .O(N__20535),
            .I(N__20527));
    InMux I__3349 (
            .O(N__20534),
            .I(N__20524));
    LocalMux I__3348 (
            .O(N__20527),
            .I(\POWERLED.count_1_12 ));
    LocalMux I__3347 (
            .O(N__20524),
            .I(\POWERLED.count_1_12 ));
    InMux I__3346 (
            .O(N__20519),
            .I(N__20514));
    CascadeMux I__3345 (
            .O(N__20518),
            .I(N__20511));
    InMux I__3344 (
            .O(N__20517),
            .I(N__20508));
    LocalMux I__3343 (
            .O(N__20514),
            .I(N__20505));
    InMux I__3342 (
            .O(N__20511),
            .I(N__20502));
    LocalMux I__3341 (
            .O(N__20508),
            .I(N__20499));
    Span4Mux_v I__3340 (
            .O(N__20505),
            .I(N__20494));
    LocalMux I__3339 (
            .O(N__20502),
            .I(N__20494));
    Odrv4 I__3338 (
            .O(N__20499),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__3337 (
            .O(N__20494),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__3336 (
            .O(N__20489),
            .I(N__20486));
    LocalMux I__3335 (
            .O(N__20486),
            .I(N__20480));
    CascadeMux I__3334 (
            .O(N__20485),
            .I(N__20477));
    InMux I__3333 (
            .O(N__20484),
            .I(N__20474));
    CascadeMux I__3332 (
            .O(N__20483),
            .I(N__20471));
    Span4Mux_v I__3331 (
            .O(N__20480),
            .I(N__20468));
    InMux I__3330 (
            .O(N__20477),
            .I(N__20465));
    LocalMux I__3329 (
            .O(N__20474),
            .I(N__20462));
    InMux I__3328 (
            .O(N__20471),
            .I(N__20459));
    Odrv4 I__3327 (
            .O(N__20468),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__3326 (
            .O(N__20465),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__3325 (
            .O(N__20462),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__3324 (
            .O(N__20459),
            .I(\POWERLED.countZ0Z_9 ));
    CascadeMux I__3323 (
            .O(N__20450),
            .I(\POWERLED.un79_clk_100khzlto15_3_cascade_ ));
    InMux I__3322 (
            .O(N__20447),
            .I(N__20444));
    LocalMux I__3321 (
            .O(N__20444),
            .I(N__20441));
    Odrv12 I__3320 (
            .O(N__20441),
            .I(\POWERLED.un79_clk_100khzlto15_6 ));
    CascadeMux I__3319 (
            .O(N__20438),
            .I(N__20435));
    InMux I__3318 (
            .O(N__20435),
            .I(N__20432));
    LocalMux I__3317 (
            .O(N__20432),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__3316 (
            .O(N__20429),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__3315 (
            .O(N__20426),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__3314 (
            .O(N__20423),
            .I(N__20418));
    InMux I__3313 (
            .O(N__20422),
            .I(N__20413));
    InMux I__3312 (
            .O(N__20421),
            .I(N__20410));
    InMux I__3311 (
            .O(N__20418),
            .I(N__20405));
    InMux I__3310 (
            .O(N__20417),
            .I(N__20405));
    InMux I__3309 (
            .O(N__20416),
            .I(N__20402));
    LocalMux I__3308 (
            .O(N__20413),
            .I(N__20399));
    LocalMux I__3307 (
            .O(N__20410),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3306 (
            .O(N__20405),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3305 (
            .O(N__20402),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    Odrv4 I__3304 (
            .O(N__20399),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    InMux I__3303 (
            .O(N__20390),
            .I(N__20387));
    LocalMux I__3302 (
            .O(N__20387),
            .I(\POWERLED.mult1_un54_sum_i ));
    CascadeMux I__3301 (
            .O(N__20384),
            .I(N__20381));
    InMux I__3300 (
            .O(N__20381),
            .I(N__20378));
    LocalMux I__3299 (
            .O(N__20378),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__3298 (
            .O(N__20375),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    InMux I__3297 (
            .O(N__20372),
            .I(N__20369));
    LocalMux I__3296 (
            .O(N__20369),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__3295 (
            .O(N__20366),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    CascadeMux I__3294 (
            .O(N__20363),
            .I(N__20360));
    InMux I__3293 (
            .O(N__20360),
            .I(N__20357));
    LocalMux I__3292 (
            .O(N__20357),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__3291 (
            .O(N__20354),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    InMux I__3290 (
            .O(N__20351),
            .I(N__20348));
    LocalMux I__3289 (
            .O(N__20348),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    InMux I__3288 (
            .O(N__20345),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    CascadeMux I__3287 (
            .O(N__20342),
            .I(N__20339));
    InMux I__3286 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__3285 (
            .O(N__20336),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__3284 (
            .O(N__20333),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__3283 (
            .O(N__20330),
            .I(N__20326));
    CascadeMux I__3282 (
            .O(N__20329),
            .I(N__20322));
    InMux I__3281 (
            .O(N__20326),
            .I(N__20315));
    InMux I__3280 (
            .O(N__20325),
            .I(N__20315));
    InMux I__3279 (
            .O(N__20322),
            .I(N__20315));
    LocalMux I__3278 (
            .O(N__20315),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    InMux I__3277 (
            .O(N__20312),
            .I(N__20309));
    LocalMux I__3276 (
            .O(N__20309),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__3275 (
            .O(N__20306),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__3274 (
            .O(N__20303),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    CascadeMux I__3273 (
            .O(N__20300),
            .I(N__20297));
    InMux I__3272 (
            .O(N__20297),
            .I(N__20287));
    InMux I__3271 (
            .O(N__20296),
            .I(N__20287));
    InMux I__3270 (
            .O(N__20295),
            .I(N__20287));
    InMux I__3269 (
            .O(N__20294),
            .I(N__20284));
    LocalMux I__3268 (
            .O(N__20287),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__3267 (
            .O(N__20284),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    CascadeMux I__3266 (
            .O(N__20279),
            .I(\POWERLED.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__3265 (
            .O(N__20276),
            .I(N__20273));
    InMux I__3264 (
            .O(N__20273),
            .I(N__20270));
    LocalMux I__3263 (
            .O(N__20270),
            .I(N__20267));
    Odrv4 I__3262 (
            .O(N__20267),
            .I(\POWERLED.mult1_un75_sum_i_8 ));
    InMux I__3261 (
            .O(N__20264),
            .I(N__20261));
    LocalMux I__3260 (
            .O(N__20261),
            .I(N__20258));
    Odrv12 I__3259 (
            .O(N__20258),
            .I(\POWERLED.mult1_un61_sum_i ));
    CascadeMux I__3258 (
            .O(N__20255),
            .I(N__20252));
    InMux I__3257 (
            .O(N__20252),
            .I(N__20249));
    LocalMux I__3256 (
            .O(N__20249),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__3255 (
            .O(N__20246),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    CascadeMux I__3254 (
            .O(N__20243),
            .I(N__20240));
    InMux I__3253 (
            .O(N__20240),
            .I(N__20237));
    LocalMux I__3252 (
            .O(N__20237),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__3251 (
            .O(N__20234),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    InMux I__3250 (
            .O(N__20231),
            .I(N__20228));
    LocalMux I__3249 (
            .O(N__20228),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__3248 (
            .O(N__20225),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__3247 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__3246 (
            .O(N__20219),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__3245 (
            .O(N__20216),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    CascadeMux I__3244 (
            .O(N__20213),
            .I(N__20210));
    InMux I__3243 (
            .O(N__20210),
            .I(N__20207));
    LocalMux I__3242 (
            .O(N__20207),
            .I(N__20204));
    Odrv12 I__3241 (
            .O(N__20204),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__3240 (
            .O(N__20201),
            .I(N__20198));
    LocalMux I__3239 (
            .O(N__20198),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__3238 (
            .O(N__20195),
            .I(N__20192));
    LocalMux I__3237 (
            .O(N__20192),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__3236 (
            .O(N__20189),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    CascadeMux I__3235 (
            .O(N__20186),
            .I(N__20183));
    InMux I__3234 (
            .O(N__20183),
            .I(N__20180));
    LocalMux I__3233 (
            .O(N__20180),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__3232 (
            .O(N__20177),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__3231 (
            .O(N__20174),
            .I(N__20171));
    LocalMux I__3230 (
            .O(N__20171),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__3229 (
            .O(N__20168),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    CascadeMux I__3228 (
            .O(N__20165),
            .I(N__20162));
    InMux I__3227 (
            .O(N__20162),
            .I(N__20159));
    LocalMux I__3226 (
            .O(N__20159),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__3225 (
            .O(N__20156),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    CascadeMux I__3224 (
            .O(N__20153),
            .I(N__20149));
    InMux I__3223 (
            .O(N__20152),
            .I(N__20141));
    InMux I__3222 (
            .O(N__20149),
            .I(N__20141));
    InMux I__3221 (
            .O(N__20148),
            .I(N__20141));
    LocalMux I__3220 (
            .O(N__20141),
            .I(G_2161));
    InMux I__3219 (
            .O(N__20138),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__3218 (
            .O(N__20135),
            .I(N__20132));
    InMux I__3217 (
            .O(N__20132),
            .I(N__20129));
    LocalMux I__3216 (
            .O(N__20129),
            .I(N__20126));
    Span4Mux_v I__3215 (
            .O(N__20126),
            .I(N__20123));
    Odrv4 I__3214 (
            .O(N__20123),
            .I(\POWERLED.mult1_un166_sum_i_8 ));
    InMux I__3213 (
            .O(N__20120),
            .I(N__20117));
    LocalMux I__3212 (
            .O(N__20117),
            .I(N__20114));
    Span4Mux_h I__3211 (
            .O(N__20114),
            .I(N__20111));
    Odrv4 I__3210 (
            .O(N__20111),
            .I(\POWERLED.mult1_un145_sum_i_8 ));
    CascadeMux I__3209 (
            .O(N__20108),
            .I(N__20105));
    InMux I__3208 (
            .O(N__20105),
            .I(N__20102));
    LocalMux I__3207 (
            .O(N__20102),
            .I(\COUNTER.un4_counter_4_and ));
    CascadeMux I__3206 (
            .O(N__20099),
            .I(N__20096));
    InMux I__3205 (
            .O(N__20096),
            .I(N__20093));
    LocalMux I__3204 (
            .O(N__20093),
            .I(N__20090));
    Odrv4 I__3203 (
            .O(N__20090),
            .I(\COUNTER.un4_counter_5_and ));
    CascadeMux I__3202 (
            .O(N__20087),
            .I(N__20084));
    InMux I__3201 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__3200 (
            .O(N__20081),
            .I(N__20078));
    Odrv4 I__3199 (
            .O(N__20078),
            .I(\COUNTER.un4_counter_6_and ));
    CascadeMux I__3198 (
            .O(N__20075),
            .I(N__20072));
    InMux I__3197 (
            .O(N__20072),
            .I(N__20069));
    LocalMux I__3196 (
            .O(N__20069),
            .I(N__20066));
    Span4Mux_h I__3195 (
            .O(N__20066),
            .I(N__20063));
    Odrv4 I__3194 (
            .O(N__20063),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__3193 (
            .O(N__20060),
            .I(bfn_6_6_0_));
    CascadeMux I__3192 (
            .O(N__20057),
            .I(N__20054));
    InMux I__3191 (
            .O(N__20054),
            .I(N__20051));
    LocalMux I__3190 (
            .O(N__20051),
            .I(\POWERLED.mult1_un159_sum_i ));
    CascadeMux I__3189 (
            .O(N__20048),
            .I(N__20043));
    CEMux I__3188 (
            .O(N__20047),
            .I(N__20036));
    CEMux I__3187 (
            .O(N__20046),
            .I(N__20031));
    InMux I__3186 (
            .O(N__20043),
            .I(N__20018));
    CEMux I__3185 (
            .O(N__20042),
            .I(N__20018));
    InMux I__3184 (
            .O(N__20041),
            .I(N__20013));
    CEMux I__3183 (
            .O(N__20040),
            .I(N__20013));
    CascadeMux I__3182 (
            .O(N__20039),
            .I(N__20010));
    LocalMux I__3181 (
            .O(N__20036),
            .I(N__20005));
    CEMux I__3180 (
            .O(N__20035),
            .I(N__20002));
    CEMux I__3179 (
            .O(N__20034),
            .I(N__19999));
    LocalMux I__3178 (
            .O(N__20031),
            .I(N__19996));
    InMux I__3177 (
            .O(N__20030),
            .I(N__19989));
    InMux I__3176 (
            .O(N__20029),
            .I(N__19989));
    InMux I__3175 (
            .O(N__20028),
            .I(N__19989));
    InMux I__3174 (
            .O(N__20027),
            .I(N__19984));
    InMux I__3173 (
            .O(N__20026),
            .I(N__19984));
    InMux I__3172 (
            .O(N__20025),
            .I(N__19981));
    InMux I__3171 (
            .O(N__20024),
            .I(N__19974));
    CEMux I__3170 (
            .O(N__20023),
            .I(N__19974));
    LocalMux I__3169 (
            .O(N__20018),
            .I(N__19971));
    LocalMux I__3168 (
            .O(N__20013),
            .I(N__19968));
    InMux I__3167 (
            .O(N__20010),
            .I(N__19961));
    InMux I__3166 (
            .O(N__20009),
            .I(N__19961));
    InMux I__3165 (
            .O(N__20008),
            .I(N__19961));
    Span4Mux_v I__3164 (
            .O(N__20005),
            .I(N__19954));
    LocalMux I__3163 (
            .O(N__20002),
            .I(N__19954));
    LocalMux I__3162 (
            .O(N__19999),
            .I(N__19949));
    Span4Mux_s0_v I__3161 (
            .O(N__19996),
            .I(N__19940));
    LocalMux I__3160 (
            .O(N__19989),
            .I(N__19940));
    LocalMux I__3159 (
            .O(N__19984),
            .I(N__19940));
    LocalMux I__3158 (
            .O(N__19981),
            .I(N__19940));
    InMux I__3157 (
            .O(N__19980),
            .I(N__19935));
    InMux I__3156 (
            .O(N__19979),
            .I(N__19935));
    LocalMux I__3155 (
            .O(N__19974),
            .I(N__19931));
    Span4Mux_s2_v I__3154 (
            .O(N__19971),
            .I(N__19924));
    Span4Mux_s2_v I__3153 (
            .O(N__19968),
            .I(N__19924));
    LocalMux I__3152 (
            .O(N__19961),
            .I(N__19924));
    InMux I__3151 (
            .O(N__19960),
            .I(N__19919));
    InMux I__3150 (
            .O(N__19959),
            .I(N__19919));
    Span4Mux_h I__3149 (
            .O(N__19954),
            .I(N__19916));
    InMux I__3148 (
            .O(N__19953),
            .I(N__19913));
    InMux I__3147 (
            .O(N__19952),
            .I(N__19910));
    Span4Mux_v I__3146 (
            .O(N__19949),
            .I(N__19903));
    Span4Mux_v I__3145 (
            .O(N__19940),
            .I(N__19903));
    LocalMux I__3144 (
            .O(N__19935),
            .I(N__19903));
    InMux I__3143 (
            .O(N__19934),
            .I(N__19900));
    Span4Mux_h I__3142 (
            .O(N__19931),
            .I(N__19893));
    Span4Mux_v I__3141 (
            .O(N__19924),
            .I(N__19893));
    LocalMux I__3140 (
            .O(N__19919),
            .I(N__19893));
    Odrv4 I__3139 (
            .O(N__19916),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    LocalMux I__3138 (
            .O(N__19913),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    LocalMux I__3137 (
            .O(N__19910),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    Odrv4 I__3136 (
            .O(N__19903),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    LocalMux I__3135 (
            .O(N__19900),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    Odrv4 I__3134 (
            .O(N__19893),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    CascadeMux I__3133 (
            .O(N__19880),
            .I(\VPP_VDDQ.count_2_1_11_cascade_ ));
    InMux I__3132 (
            .O(N__19877),
            .I(N__19874));
    LocalMux I__3131 (
            .O(N__19874),
            .I(\VPP_VDDQ.count_2_0_11 ));
    InMux I__3130 (
            .O(N__19871),
            .I(N__19867));
    InMux I__3129 (
            .O(N__19870),
            .I(N__19864));
    LocalMux I__3128 (
            .O(N__19867),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    LocalMux I__3127 (
            .O(N__19864),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    SRMux I__3126 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__3125 (
            .O(N__19856),
            .I(N__19853));
    Span4Mux_s2_v I__3124 (
            .O(N__19853),
            .I(N__19850));
    Span4Mux_h I__3123 (
            .O(N__19850),
            .I(N__19847));
    Odrv4 I__3122 (
            .O(N__19847),
            .I(\VPP_VDDQ.N_60_i ));
    CascadeMux I__3121 (
            .O(N__19844),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_ ));
    InMux I__3120 (
            .O(N__19841),
            .I(N__19835));
    InMux I__3119 (
            .O(N__19840),
            .I(N__19835));
    LocalMux I__3118 (
            .O(N__19835),
            .I(N__19831));
    InMux I__3117 (
            .O(N__19834),
            .I(N__19828));
    Odrv4 I__3116 (
            .O(N__19831),
            .I(\VPP_VDDQ.N_60 ));
    LocalMux I__3115 (
            .O(N__19828),
            .I(\VPP_VDDQ.N_60 ));
    CascadeMux I__3114 (
            .O(N__19823),
            .I(\VPP_VDDQ.N_60_cascade_ ));
    CascadeMux I__3113 (
            .O(N__19820),
            .I(N__19816));
    InMux I__3112 (
            .O(N__19819),
            .I(N__19811));
    InMux I__3111 (
            .O(N__19816),
            .I(N__19811));
    LocalMux I__3110 (
            .O(N__19811),
            .I(N__19808));
    Odrv4 I__3109 (
            .O(N__19808),
            .I(\VPP_VDDQ.delayed_vddq_ok_en ));
    CascadeMux I__3108 (
            .O(N__19805),
            .I(N__19802));
    InMux I__3107 (
            .O(N__19802),
            .I(N__19799));
    LocalMux I__3106 (
            .O(N__19799),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__3105 (
            .O(N__19796),
            .I(N__19793));
    InMux I__3104 (
            .O(N__19793),
            .I(N__19790));
    LocalMux I__3103 (
            .O(N__19790),
            .I(\COUNTER.un4_counter_1_and ));
    CascadeMux I__3102 (
            .O(N__19787),
            .I(N__19784));
    InMux I__3101 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__3100 (
            .O(N__19781),
            .I(\COUNTER.un4_counter_2_and ));
    CascadeMux I__3099 (
            .O(N__19778),
            .I(N__19775));
    InMux I__3098 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__3097 (
            .O(N__19772),
            .I(\COUNTER.un4_counter_3_and ));
    IoInMux I__3096 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__3095 (
            .O(N__19766),
            .I(N__19763));
    Span4Mux_s2_h I__3094 (
            .O(N__19763),
            .I(N__19759));
    InMux I__3093 (
            .O(N__19762),
            .I(N__19756));
    Sp12to4 I__3092 (
            .O(N__19759),
            .I(N__19753));
    LocalMux I__3091 (
            .O(N__19756),
            .I(N__19750));
    Span12Mux_s11_v I__3090 (
            .O(N__19753),
            .I(N__19747));
    Span12Mux_s11_v I__3089 (
            .O(N__19750),
            .I(N__19744));
    Odrv12 I__3088 (
            .O(N__19747),
            .I(v1p8a_ok));
    Odrv12 I__3087 (
            .O(N__19744),
            .I(v1p8a_ok));
    InMux I__3086 (
            .O(N__19739),
            .I(N__19736));
    LocalMux I__3085 (
            .O(N__19736),
            .I(N__19733));
    Span4Mux_v I__3084 (
            .O(N__19733),
            .I(N__19730));
    Span4Mux_h I__3083 (
            .O(N__19730),
            .I(N__19727));
    Odrv4 I__3082 (
            .O(N__19727),
            .I(v5a_ok));
    IoInMux I__3081 (
            .O(N__19724),
            .I(N__19721));
    LocalMux I__3080 (
            .O(N__19721),
            .I(N__19717));
    InMux I__3079 (
            .O(N__19720),
            .I(N__19714));
    IoSpan4Mux I__3078 (
            .O(N__19717),
            .I(N__19711));
    LocalMux I__3077 (
            .O(N__19714),
            .I(N__19707));
    IoSpan4Mux I__3076 (
            .O(N__19711),
            .I(N__19704));
    IoInMux I__3075 (
            .O(N__19710),
            .I(N__19701));
    Span4Mux_s2_v I__3074 (
            .O(N__19707),
            .I(N__19698));
    IoSpan4Mux I__3073 (
            .O(N__19704),
            .I(N__19693));
    LocalMux I__3072 (
            .O(N__19701),
            .I(N__19693));
    Sp12to4 I__3071 (
            .O(N__19698),
            .I(N__19690));
    IoSpan4Mux I__3070 (
            .O(N__19693),
            .I(N__19687));
    Span12Mux_s11_h I__3069 (
            .O(N__19690),
            .I(N__19684));
    IoSpan4Mux I__3068 (
            .O(N__19687),
            .I(N__19681));
    Span12Mux_v I__3067 (
            .O(N__19684),
            .I(N__19678));
    IoSpan4Mux I__3066 (
            .O(N__19681),
            .I(N__19675));
    Odrv12 I__3065 (
            .O(N__19678),
            .I(v33a_ok));
    Odrv4 I__3064 (
            .O(N__19675),
            .I(v33a_ok));
    CascadeMux I__3063 (
            .O(N__19670),
            .I(N__19666));
    InMux I__3062 (
            .O(N__19669),
            .I(N__19661));
    InMux I__3061 (
            .O(N__19666),
            .I(N__19661));
    LocalMux I__3060 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_v I__3059 (
            .O(N__19658),
            .I(N__19655));
    Sp12to4 I__3058 (
            .O(N__19655),
            .I(N__19652));
    Span12Mux_s8_h I__3057 (
            .O(N__19652),
            .I(N__19649));
    Odrv12 I__3056 (
            .O(N__19649),
            .I(slp_susn));
    IoInMux I__3055 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__3054 (
            .O(N__19643),
            .I(N__19640));
    Span4Mux_s3_h I__3053 (
            .O(N__19640),
            .I(N__19637));
    Span4Mux_v I__3052 (
            .O(N__19637),
            .I(N__19634));
    Span4Mux_v I__3051 (
            .O(N__19634),
            .I(N__19631));
    Odrv4 I__3050 (
            .O(N__19631),
            .I(v33a_enn));
    CascadeMux I__3049 (
            .O(N__19628),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ));
    CascadeMux I__3048 (
            .O(N__19625),
            .I(\VPP_VDDQ.count_2_1_1_cascade_ ));
    InMux I__3047 (
            .O(N__19622),
            .I(N__19618));
    InMux I__3046 (
            .O(N__19621),
            .I(N__19615));
    LocalMux I__3045 (
            .O(N__19618),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    LocalMux I__3044 (
            .O(N__19615),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    InMux I__3043 (
            .O(N__19610),
            .I(N__19607));
    LocalMux I__3042 (
            .O(N__19607),
            .I(\VPP_VDDQ.count_2_1_1 ));
    CascadeMux I__3041 (
            .O(N__19604),
            .I(N__19600));
    CascadeMux I__3040 (
            .O(N__19603),
            .I(N__19596));
    InMux I__3039 (
            .O(N__19600),
            .I(N__19592));
    InMux I__3038 (
            .O(N__19599),
            .I(N__19589));
    InMux I__3037 (
            .O(N__19596),
            .I(N__19584));
    InMux I__3036 (
            .O(N__19595),
            .I(N__19584));
    LocalMux I__3035 (
            .O(N__19592),
            .I(N__19581));
    LocalMux I__3034 (
            .O(N__19589),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__3033 (
            .O(N__19584),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    Odrv4 I__3032 (
            .O(N__19581),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    InMux I__3031 (
            .O(N__19574),
            .I(N__19571));
    LocalMux I__3030 (
            .O(N__19571),
            .I(\VPP_VDDQ.un9_clk_100khz_1 ));
    InMux I__3029 (
            .O(N__19568),
            .I(N__19565));
    LocalMux I__3028 (
            .O(N__19565),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1 ));
    InMux I__3027 (
            .O(N__19562),
            .I(N__19556));
    InMux I__3026 (
            .O(N__19561),
            .I(N__19556));
    LocalMux I__3025 (
            .O(N__19556),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    InMux I__3024 (
            .O(N__19553),
            .I(N__19547));
    InMux I__3023 (
            .O(N__19552),
            .I(N__19547));
    LocalMux I__3022 (
            .O(N__19547),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ));
    InMux I__3021 (
            .O(N__19544),
            .I(N__19538));
    InMux I__3020 (
            .O(N__19543),
            .I(N__19538));
    LocalMux I__3019 (
            .O(N__19538),
            .I(\VPP_VDDQ.delayed_vddq_okZ0 ));
    CascadeMux I__3018 (
            .O(N__19535),
            .I(VPP_VDDQ_delayed_vddq_ok_cascade_));
    IoInMux I__3017 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__3016 (
            .O(N__19529),
            .I(vccst_pwrgd));
    InMux I__3015 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__3014 (
            .O(N__19523),
            .I(N__19519));
    InMux I__3013 (
            .O(N__19522),
            .I(N__19516));
    Odrv4 I__3012 (
            .O(N__19519),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    LocalMux I__3011 (
            .O(N__19516),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    InMux I__3010 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__3009 (
            .O(N__19508),
            .I(\VPP_VDDQ.un9_clk_100khz_9 ));
    CascadeMux I__3008 (
            .O(N__19505),
            .I(\VPP_VDDQ.un9_clk_100khz_0_cascade_ ));
    InMux I__3007 (
            .O(N__19502),
            .I(N__19499));
    LocalMux I__3006 (
            .O(N__19499),
            .I(N__19496));
    Odrv4 I__3005 (
            .O(N__19496),
            .I(\VPP_VDDQ.un9_clk_100khz_13 ));
    InMux I__3004 (
            .O(N__19493),
            .I(N__19487));
    InMux I__3003 (
            .O(N__19492),
            .I(N__19487));
    LocalMux I__3002 (
            .O(N__19487),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ));
    CascadeMux I__3001 (
            .O(N__19484),
            .I(\VPP_VDDQ.N_1_i_cascade_ ));
    InMux I__3000 (
            .O(N__19481),
            .I(N__19478));
    LocalMux I__2999 (
            .O(N__19478),
            .I(\VPP_VDDQ.count_2_1_6 ));
    CascadeMux I__2998 (
            .O(N__19475),
            .I(\VPP_VDDQ.count_2_1_6_cascade_ ));
    InMux I__2997 (
            .O(N__19472),
            .I(N__19466));
    InMux I__2996 (
            .O(N__19471),
            .I(N__19466));
    LocalMux I__2995 (
            .O(N__19466),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    InMux I__2994 (
            .O(N__19463),
            .I(N__19460));
    LocalMux I__2993 (
            .O(N__19460),
            .I(\VPP_VDDQ.un1_count_2_1_axb_6 ));
    CascadeMux I__2992 (
            .O(N__19457),
            .I(N__19453));
    InMux I__2991 (
            .O(N__19456),
            .I(N__19448));
    InMux I__2990 (
            .O(N__19453),
            .I(N__19448));
    LocalMux I__2989 (
            .O(N__19448),
            .I(\POWERLED.count_1_9 ));
    InMux I__2988 (
            .O(N__19445),
            .I(N__19442));
    LocalMux I__2987 (
            .O(N__19442),
            .I(\POWERLED.count_0_9 ));
    InMux I__2986 (
            .O(N__19439),
            .I(N__19436));
    LocalMux I__2985 (
            .O(N__19436),
            .I(N__19431));
    InMux I__2984 (
            .O(N__19435),
            .I(N__19428));
    InMux I__2983 (
            .O(N__19434),
            .I(N__19425));
    Odrv4 I__2982 (
            .O(N__19431),
            .I(\POWERLED.count_1_10 ));
    LocalMux I__2981 (
            .O(N__19428),
            .I(\POWERLED.count_1_10 ));
    LocalMux I__2980 (
            .O(N__19425),
            .I(\POWERLED.count_1_10 ));
    InMux I__2979 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__2978 (
            .O(N__19415),
            .I(\POWERLED.count_0_10 ));
    InMux I__2977 (
            .O(N__19412),
            .I(N__19407));
    InMux I__2976 (
            .O(N__19411),
            .I(N__19404));
    CascadeMux I__2975 (
            .O(N__19410),
            .I(N__19401));
    LocalMux I__2974 (
            .O(N__19407),
            .I(N__19398));
    LocalMux I__2973 (
            .O(N__19404),
            .I(N__19395));
    InMux I__2972 (
            .O(N__19401),
            .I(N__19392));
    Span4Mux_h I__2971 (
            .O(N__19398),
            .I(N__19389));
    Span4Mux_v I__2970 (
            .O(N__19395),
            .I(N__19384));
    LocalMux I__2969 (
            .O(N__19392),
            .I(N__19384));
    Odrv4 I__2968 (
            .O(N__19389),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__2967 (
            .O(N__19384),
            .I(\POWERLED.countZ0Z_6 ));
    InMux I__2966 (
            .O(N__19379),
            .I(N__19374));
    InMux I__2965 (
            .O(N__19378),
            .I(N__19369));
    InMux I__2964 (
            .O(N__19377),
            .I(N__19369));
    LocalMux I__2963 (
            .O(N__19374),
            .I(N__19366));
    LocalMux I__2962 (
            .O(N__19369),
            .I(N__19363));
    Odrv12 I__2961 (
            .O(N__19366),
            .I(\POWERLED.count_1_6 ));
    Odrv4 I__2960 (
            .O(N__19363),
            .I(\POWERLED.count_1_6 ));
    InMux I__2959 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__2958 (
            .O(N__19355),
            .I(\POWERLED.count_0_6 ));
    InMux I__2957 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__2956 (
            .O(N__19349),
            .I(N__19344));
    InMux I__2955 (
            .O(N__19348),
            .I(N__19341));
    InMux I__2954 (
            .O(N__19347),
            .I(N__19338));
    Span4Mux_s3_v I__2953 (
            .O(N__19344),
            .I(N__19335));
    LocalMux I__2952 (
            .O(N__19341),
            .I(N__19330));
    LocalMux I__2951 (
            .O(N__19338),
            .I(N__19330));
    Odrv4 I__2950 (
            .O(N__19335),
            .I(\POWERLED.count_1_8 ));
    Odrv4 I__2949 (
            .O(N__19330),
            .I(\POWERLED.count_1_8 ));
    InMux I__2948 (
            .O(N__19325),
            .I(N__19322));
    LocalMux I__2947 (
            .O(N__19322),
            .I(N__19319));
    Odrv4 I__2946 (
            .O(N__19319),
            .I(\POWERLED.count_0_8 ));
    InMux I__2945 (
            .O(N__19316),
            .I(N__19312));
    InMux I__2944 (
            .O(N__19315),
            .I(N__19309));
    LocalMux I__2943 (
            .O(N__19312),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    LocalMux I__2942 (
            .O(N__19309),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    InMux I__2941 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__2940 (
            .O(N__19301),
            .I(\VPP_VDDQ.count_2_0_3 ));
    CascadeMux I__2939 (
            .O(N__19298),
            .I(\VPP_VDDQ.count_2_1_3_cascade_ ));
    InMux I__2938 (
            .O(N__19295),
            .I(N__19291));
    InMux I__2937 (
            .O(N__19294),
            .I(N__19288));
    LocalMux I__2936 (
            .O(N__19291),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    LocalMux I__2935 (
            .O(N__19288),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    InMux I__2934 (
            .O(N__19283),
            .I(bfn_5_14_0_));
    InMux I__2933 (
            .O(N__19280),
            .I(N__19277));
    LocalMux I__2932 (
            .O(N__19277),
            .I(N__19273));
    CascadeMux I__2931 (
            .O(N__19276),
            .I(N__19269));
    Span4Mux_v I__2930 (
            .O(N__19273),
            .I(N__19266));
    InMux I__2929 (
            .O(N__19272),
            .I(N__19263));
    InMux I__2928 (
            .O(N__19269),
            .I(N__19260));
    Odrv4 I__2927 (
            .O(N__19266),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__2926 (
            .O(N__19263),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__2925 (
            .O(N__19260),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__2924 (
            .O(N__19253),
            .I(\POWERLED.un1_count_cry_9 ));
    InMux I__2923 (
            .O(N__19250),
            .I(N__19246));
    CascadeMux I__2922 (
            .O(N__19249),
            .I(N__19242));
    LocalMux I__2921 (
            .O(N__19246),
            .I(N__19239));
    InMux I__2920 (
            .O(N__19245),
            .I(N__19236));
    InMux I__2919 (
            .O(N__19242),
            .I(N__19233));
    Odrv12 I__2918 (
            .O(N__19239),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__2917 (
            .O(N__19236),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__2916 (
            .O(N__19233),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__2915 (
            .O(N__19226),
            .I(N__19222));
    CascadeMux I__2914 (
            .O(N__19225),
            .I(N__19219));
    LocalMux I__2913 (
            .O(N__19222),
            .I(N__19215));
    InMux I__2912 (
            .O(N__19219),
            .I(N__19210));
    InMux I__2911 (
            .O(N__19218),
            .I(N__19210));
    Odrv4 I__2910 (
            .O(N__19215),
            .I(\POWERLED.count_1_11 ));
    LocalMux I__2909 (
            .O(N__19210),
            .I(\POWERLED.count_1_11 ));
    InMux I__2908 (
            .O(N__19205),
            .I(\POWERLED.un1_count_cry_10 ));
    InMux I__2907 (
            .O(N__19202),
            .I(\POWERLED.un1_count_cry_11 ));
    InMux I__2906 (
            .O(N__19199),
            .I(\POWERLED.un1_count_cry_12 ));
    CascadeMux I__2905 (
            .O(N__19196),
            .I(N__19193));
    InMux I__2904 (
            .O(N__19193),
            .I(N__19187));
    InMux I__2903 (
            .O(N__19192),
            .I(N__19187));
    LocalMux I__2902 (
            .O(N__19187),
            .I(\POWERLED.count_1_14 ));
    InMux I__2901 (
            .O(N__19184),
            .I(\POWERLED.un1_count_cry_13 ));
    InMux I__2900 (
            .O(N__19181),
            .I(N__19176));
    InMux I__2899 (
            .O(N__19180),
            .I(N__19167));
    InMux I__2898 (
            .O(N__19179),
            .I(N__19167));
    LocalMux I__2897 (
            .O(N__19176),
            .I(N__19164));
    InMux I__2896 (
            .O(N__19175),
            .I(N__19151));
    InMux I__2895 (
            .O(N__19174),
            .I(N__19151));
    InMux I__2894 (
            .O(N__19173),
            .I(N__19151));
    InMux I__2893 (
            .O(N__19172),
            .I(N__19151));
    LocalMux I__2892 (
            .O(N__19167),
            .I(N__19148));
    Span4Mux_v I__2891 (
            .O(N__19164),
            .I(N__19138));
    InMux I__2890 (
            .O(N__19163),
            .I(N__19131));
    InMux I__2889 (
            .O(N__19162),
            .I(N__19131));
    InMux I__2888 (
            .O(N__19161),
            .I(N__19131));
    InMux I__2887 (
            .O(N__19160),
            .I(N__19128));
    LocalMux I__2886 (
            .O(N__19151),
            .I(N__19123));
    Span4Mux_v I__2885 (
            .O(N__19148),
            .I(N__19123));
    InMux I__2884 (
            .O(N__19147),
            .I(N__19114));
    InMux I__2883 (
            .O(N__19146),
            .I(N__19114));
    InMux I__2882 (
            .O(N__19145),
            .I(N__19114));
    InMux I__2881 (
            .O(N__19144),
            .I(N__19114));
    InMux I__2880 (
            .O(N__19143),
            .I(N__19107));
    InMux I__2879 (
            .O(N__19142),
            .I(N__19107));
    InMux I__2878 (
            .O(N__19141),
            .I(N__19107));
    Odrv4 I__2877 (
            .O(N__19138),
            .I(\POWERLED.count_0_sqmuxa ));
    LocalMux I__2876 (
            .O(N__19131),
            .I(\POWERLED.count_0_sqmuxa ));
    LocalMux I__2875 (
            .O(N__19128),
            .I(\POWERLED.count_0_sqmuxa ));
    Odrv4 I__2874 (
            .O(N__19123),
            .I(\POWERLED.count_0_sqmuxa ));
    LocalMux I__2873 (
            .O(N__19114),
            .I(\POWERLED.count_0_sqmuxa ));
    LocalMux I__2872 (
            .O(N__19107),
            .I(\POWERLED.count_0_sqmuxa ));
    InMux I__2871 (
            .O(N__19094),
            .I(\POWERLED.un1_count_cry_14 ));
    CascadeMux I__2870 (
            .O(N__19091),
            .I(N__19088));
    InMux I__2869 (
            .O(N__19088),
            .I(N__19084));
    InMux I__2868 (
            .O(N__19087),
            .I(N__19081));
    LocalMux I__2867 (
            .O(N__19084),
            .I(N__19078));
    LocalMux I__2866 (
            .O(N__19081),
            .I(\POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ));
    Odrv4 I__2865 (
            .O(N__19078),
            .I(\POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ));
    CascadeMux I__2864 (
            .O(N__19073),
            .I(N__19070));
    InMux I__2863 (
            .O(N__19070),
            .I(N__19067));
    LocalMux I__2862 (
            .O(N__19067),
            .I(\POWERLED.un1_count_axb_12 ));
    InMux I__2861 (
            .O(N__19064),
            .I(N__19061));
    LocalMux I__2860 (
            .O(N__19061),
            .I(N__19054));
    InMux I__2859 (
            .O(N__19060),
            .I(N__19047));
    InMux I__2858 (
            .O(N__19059),
            .I(N__19047));
    InMux I__2857 (
            .O(N__19058),
            .I(N__19047));
    InMux I__2856 (
            .O(N__19057),
            .I(N__19044));
    Odrv12 I__2855 (
            .O(N__19054),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2854 (
            .O(N__19047),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2853 (
            .O(N__19044),
            .I(\POWERLED.countZ0Z_0 ));
    CascadeMux I__2852 (
            .O(N__19037),
            .I(N__19033));
    InMux I__2851 (
            .O(N__19036),
            .I(N__19030));
    InMux I__2850 (
            .O(N__19033),
            .I(N__19027));
    LocalMux I__2849 (
            .O(N__19030),
            .I(\POWERLED.un1_count_axb_1 ));
    LocalMux I__2848 (
            .O(N__19027),
            .I(\POWERLED.un1_count_axb_1 ));
    CascadeMux I__2847 (
            .O(N__19022),
            .I(N__19019));
    InMux I__2846 (
            .O(N__19019),
            .I(N__19016));
    LocalMux I__2845 (
            .O(N__19016),
            .I(\POWERLED.un1_count_axb_2 ));
    InMux I__2844 (
            .O(N__19013),
            .I(N__19001));
    InMux I__2843 (
            .O(N__19012),
            .I(N__19001));
    InMux I__2842 (
            .O(N__19011),
            .I(N__19001));
    InMux I__2841 (
            .O(N__19010),
            .I(N__19001));
    LocalMux I__2840 (
            .O(N__19001),
            .I(\POWERLED.count_1_2 ));
    InMux I__2839 (
            .O(N__18998),
            .I(\POWERLED.un1_count_cry_1 ));
    InMux I__2838 (
            .O(N__18995),
            .I(N__18991));
    CascadeMux I__2837 (
            .O(N__18994),
            .I(N__18987));
    LocalMux I__2836 (
            .O(N__18991),
            .I(N__18984));
    InMux I__2835 (
            .O(N__18990),
            .I(N__18981));
    InMux I__2834 (
            .O(N__18987),
            .I(N__18978));
    Odrv4 I__2833 (
            .O(N__18984),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__2832 (
            .O(N__18981),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__2831 (
            .O(N__18978),
            .I(\POWERLED.countZ0Z_3 ));
    InMux I__2830 (
            .O(N__18971),
            .I(N__18965));
    InMux I__2829 (
            .O(N__18970),
            .I(N__18965));
    LocalMux I__2828 (
            .O(N__18965),
            .I(\POWERLED.un1_count_cry_2_c_RNICZ0Z419 ));
    InMux I__2827 (
            .O(N__18962),
            .I(\POWERLED.un1_count_cry_2 ));
    CascadeMux I__2826 (
            .O(N__18959),
            .I(N__18956));
    InMux I__2825 (
            .O(N__18956),
            .I(N__18953));
    LocalMux I__2824 (
            .O(N__18953),
            .I(\POWERLED.un1_count_axb_4 ));
    CascadeMux I__2823 (
            .O(N__18950),
            .I(N__18947));
    InMux I__2822 (
            .O(N__18947),
            .I(N__18935));
    InMux I__2821 (
            .O(N__18946),
            .I(N__18935));
    InMux I__2820 (
            .O(N__18945),
            .I(N__18935));
    InMux I__2819 (
            .O(N__18944),
            .I(N__18935));
    LocalMux I__2818 (
            .O(N__18935),
            .I(\POWERLED.count_1_4 ));
    InMux I__2817 (
            .O(N__18932),
            .I(\POWERLED.un1_count_cry_3 ));
    CascadeMux I__2816 (
            .O(N__18929),
            .I(N__18926));
    InMux I__2815 (
            .O(N__18926),
            .I(N__18923));
    LocalMux I__2814 (
            .O(N__18923),
            .I(N__18920));
    Odrv4 I__2813 (
            .O(N__18920),
            .I(\POWERLED.un1_count_axb_5 ));
    InMux I__2812 (
            .O(N__18917),
            .I(N__18912));
    InMux I__2811 (
            .O(N__18916),
            .I(N__18907));
    InMux I__2810 (
            .O(N__18915),
            .I(N__18907));
    LocalMux I__2809 (
            .O(N__18912),
            .I(N__18904));
    LocalMux I__2808 (
            .O(N__18907),
            .I(N__18901));
    Odrv12 I__2807 (
            .O(N__18904),
            .I(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ));
    Odrv4 I__2806 (
            .O(N__18901),
            .I(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ));
    InMux I__2805 (
            .O(N__18896),
            .I(\POWERLED.un1_count_cry_4 ));
    InMux I__2804 (
            .O(N__18893),
            .I(\POWERLED.un1_count_cry_5 ));
    InMux I__2803 (
            .O(N__18890),
            .I(\POWERLED.un1_count_cry_6 ));
    InMux I__2802 (
            .O(N__18887),
            .I(\POWERLED.un1_count_cry_7 ));
    CascadeMux I__2801 (
            .O(N__18884),
            .I(N__18881));
    InMux I__2800 (
            .O(N__18881),
            .I(N__18878));
    LocalMux I__2799 (
            .O(N__18878),
            .I(N__18875));
    Odrv12 I__2798 (
            .O(N__18875),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__2797 (
            .O(N__18872),
            .I(N__18869));
    LocalMux I__2796 (
            .O(N__18869),
            .I(N__18866));
    Odrv12 I__2795 (
            .O(N__18866),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__2794 (
            .O(N__18863),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__2793 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__2792 (
            .O(N__18857),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__2791 (
            .O(N__18854),
            .I(N__18851));
    LocalMux I__2790 (
            .O(N__18851),
            .I(N__18848));
    Odrv4 I__2789 (
            .O(N__18848),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__2788 (
            .O(N__18845),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    CascadeMux I__2787 (
            .O(N__18842),
            .I(N__18839));
    InMux I__2786 (
            .O(N__18839),
            .I(N__18836));
    LocalMux I__2785 (
            .O(N__18836),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    CascadeMux I__2784 (
            .O(N__18833),
            .I(N__18830));
    InMux I__2783 (
            .O(N__18830),
            .I(N__18827));
    LocalMux I__2782 (
            .O(N__18827),
            .I(N__18824));
    Odrv4 I__2781 (
            .O(N__18824),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__2780 (
            .O(N__18821),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__2779 (
            .O(N__18818),
            .I(N__18815));
    LocalMux I__2778 (
            .O(N__18815),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    CascadeMux I__2777 (
            .O(N__18812),
            .I(N__18809));
    InMux I__2776 (
            .O(N__18809),
            .I(N__18806));
    LocalMux I__2775 (
            .O(N__18806),
            .I(N__18803));
    Odrv12 I__2774 (
            .O(N__18803),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__2773 (
            .O(N__18800),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    CascadeMux I__2772 (
            .O(N__18797),
            .I(N__18794));
    InMux I__2771 (
            .O(N__18794),
            .I(N__18791));
    LocalMux I__2770 (
            .O(N__18791),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__2769 (
            .O(N__18788),
            .I(N__18785));
    LocalMux I__2768 (
            .O(N__18785),
            .I(N__18782));
    Odrv4 I__2767 (
            .O(N__18782),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__2766 (
            .O(N__18779),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__2765 (
            .O(N__18776),
            .I(N__18773));
    LocalMux I__2764 (
            .O(N__18773),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__2763 (
            .O(N__18770),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    CascadeMux I__2762 (
            .O(N__18767),
            .I(N__18763));
    InMux I__2761 (
            .O(N__18766),
            .I(N__18755));
    InMux I__2760 (
            .O(N__18763),
            .I(N__18755));
    InMux I__2759 (
            .O(N__18762),
            .I(N__18755));
    LocalMux I__2758 (
            .O(N__18755),
            .I(N__18750));
    InMux I__2757 (
            .O(N__18754),
            .I(N__18747));
    InMux I__2756 (
            .O(N__18753),
            .I(N__18744));
    Odrv4 I__2755 (
            .O(N__18750),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2754 (
            .O(N__18747),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2753 (
            .O(N__18744),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__2752 (
            .O(N__18737),
            .I(N__18733));
    InMux I__2751 (
            .O(N__18736),
            .I(N__18727));
    InMux I__2750 (
            .O(N__18733),
            .I(N__18720));
    InMux I__2749 (
            .O(N__18732),
            .I(N__18720));
    InMux I__2748 (
            .O(N__18731),
            .I(N__18720));
    InMux I__2747 (
            .O(N__18730),
            .I(N__18717));
    LocalMux I__2746 (
            .O(N__18727),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2745 (
            .O(N__18720),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2744 (
            .O(N__18717),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__2743 (
            .O(N__18710),
            .I(N__18706));
    InMux I__2742 (
            .O(N__18709),
            .I(N__18698));
    InMux I__2741 (
            .O(N__18706),
            .I(N__18698));
    InMux I__2740 (
            .O(N__18705),
            .I(N__18698));
    LocalMux I__2739 (
            .O(N__18698),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__2738 (
            .O(N__18695),
            .I(N__18690));
    InMux I__2737 (
            .O(N__18694),
            .I(N__18687));
    CascadeMux I__2736 (
            .O(N__18693),
            .I(N__18684));
    LocalMux I__2735 (
            .O(N__18690),
            .I(N__18679));
    LocalMux I__2734 (
            .O(N__18687),
            .I(N__18676));
    InMux I__2733 (
            .O(N__18684),
            .I(N__18671));
    InMux I__2732 (
            .O(N__18683),
            .I(N__18671));
    InMux I__2731 (
            .O(N__18682),
            .I(N__18668));
    Odrv4 I__2730 (
            .O(N__18679),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    Odrv12 I__2729 (
            .O(N__18676),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2728 (
            .O(N__18671),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2727 (
            .O(N__18668),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    InMux I__2726 (
            .O(N__18659),
            .I(N__18656));
    LocalMux I__2725 (
            .O(N__18656),
            .I(\POWERLED.mult1_un124_sum_i_8 ));
    CascadeMux I__2724 (
            .O(N__18653),
            .I(N__18650));
    InMux I__2723 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__2722 (
            .O(N__18647),
            .I(N__18644));
    Odrv4 I__2721 (
            .O(N__18644),
            .I(\POWERLED.mult1_un75_sum_i ));
    InMux I__2720 (
            .O(N__18641),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    InMux I__2719 (
            .O(N__18638),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__2718 (
            .O(N__18635),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__2717 (
            .O(N__18632),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    InMux I__2716 (
            .O(N__18629),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__2715 (
            .O(N__18626),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    CascadeMux I__2714 (
            .O(N__18623),
            .I(N__18619));
    InMux I__2713 (
            .O(N__18622),
            .I(N__18611));
    InMux I__2712 (
            .O(N__18619),
            .I(N__18611));
    InMux I__2711 (
            .O(N__18618),
            .I(N__18611));
    LocalMux I__2710 (
            .O(N__18611),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    CascadeMux I__2709 (
            .O(N__18608),
            .I(N__18604));
    InMux I__2708 (
            .O(N__18607),
            .I(N__18596));
    InMux I__2707 (
            .O(N__18604),
            .I(N__18596));
    InMux I__2706 (
            .O(N__18603),
            .I(N__18596));
    LocalMux I__2705 (
            .O(N__18596),
            .I(N__18592));
    InMux I__2704 (
            .O(N__18595),
            .I(N__18589));
    Span4Mux_v I__2703 (
            .O(N__18592),
            .I(N__18584));
    LocalMux I__2702 (
            .O(N__18589),
            .I(N__18584));
    Sp12to4 I__2701 (
            .O(N__18584),
            .I(N__18580));
    InMux I__2700 (
            .O(N__18583),
            .I(N__18577));
    Odrv12 I__2699 (
            .O(N__18580),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__2698 (
            .O(N__18577),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__2697 (
            .O(N__18572),
            .I(N__18568));
    InMux I__2696 (
            .O(N__18571),
            .I(N__18560));
    InMux I__2695 (
            .O(N__18568),
            .I(N__18560));
    InMux I__2694 (
            .O(N__18567),
            .I(N__18560));
    LocalMux I__2693 (
            .O(N__18560),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    IoInMux I__2692 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__2691 (
            .O(N__18554),
            .I(N__18551));
    Span4Mux_s1_h I__2690 (
            .O(N__18551),
            .I(N__18548));
    Span4Mux_h I__2689 (
            .O(N__18548),
            .I(N__18545));
    Odrv4 I__2688 (
            .O(N__18545),
            .I(vccst_en));
    IoInMux I__2687 (
            .O(N__18542),
            .I(N__18539));
    LocalMux I__2686 (
            .O(N__18539),
            .I(N__18536));
    Odrv12 I__2685 (
            .O(N__18536),
            .I(G_12));
    CascadeMux I__2684 (
            .O(N__18533),
            .I(N__18530));
    InMux I__2683 (
            .O(N__18530),
            .I(N__18527));
    LocalMux I__2682 (
            .O(N__18527),
            .I(\POWERLED.mult1_un68_sum_i_8 ));
    CascadeMux I__2681 (
            .O(N__18524),
            .I(N__18521));
    InMux I__2680 (
            .O(N__18521),
            .I(N__18518));
    LocalMux I__2679 (
            .O(N__18518),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    CascadeMux I__2678 (
            .O(N__18515),
            .I(N__18512));
    InMux I__2677 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__2676 (
            .O(N__18509),
            .I(N__18506));
    Span4Mux_h I__2675 (
            .O(N__18506),
            .I(N__18503));
    Odrv4 I__2674 (
            .O(N__18503),
            .I(\POWERLED.mult1_un89_sum_i ));
    CascadeMux I__2673 (
            .O(N__18500),
            .I(N__18497));
    InMux I__2672 (
            .O(N__18497),
            .I(N__18494));
    LocalMux I__2671 (
            .O(N__18494),
            .I(N__18491));
    Odrv4 I__2670 (
            .O(N__18491),
            .I(\POWERLED.mult1_un117_sum_i ));
    InMux I__2669 (
            .O(N__18488),
            .I(N__18484));
    InMux I__2668 (
            .O(N__18487),
            .I(N__18481));
    LocalMux I__2667 (
            .O(N__18484),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__2666 (
            .O(N__18481),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__2665 (
            .O(N__18476),
            .I(N__18472));
    InMux I__2664 (
            .O(N__18475),
            .I(N__18469));
    LocalMux I__2663 (
            .O(N__18472),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__2662 (
            .O(N__18469),
            .I(\COUNTER.counterZ0Z_20 ));
    CascadeMux I__2661 (
            .O(N__18464),
            .I(N__18460));
    InMux I__2660 (
            .O(N__18463),
            .I(N__18457));
    InMux I__2659 (
            .O(N__18460),
            .I(N__18454));
    LocalMux I__2658 (
            .O(N__18457),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__2657 (
            .O(N__18454),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__2656 (
            .O(N__18449),
            .I(N__18445));
    InMux I__2655 (
            .O(N__18448),
            .I(N__18442));
    LocalMux I__2654 (
            .O(N__18445),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__2653 (
            .O(N__18442),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__2652 (
            .O(N__18437),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    InMux I__2651 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__2650 (
            .O(N__18431),
            .I(N__18428));
    Span4Mux_v I__2649 (
            .O(N__18428),
            .I(N__18425));
    Odrv4 I__2648 (
            .O(N__18425),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__2647 (
            .O(N__18422),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__2646 (
            .O(N__18419),
            .I(N__18416));
    LocalMux I__2645 (
            .O(N__18416),
            .I(N__18413));
    Span4Mux_v I__2644 (
            .O(N__18413),
            .I(N__18410));
    Odrv4 I__2643 (
            .O(N__18410),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__2642 (
            .O(N__18407),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    CascadeMux I__2641 (
            .O(N__18404),
            .I(N__18401));
    InMux I__2640 (
            .O(N__18401),
            .I(N__18398));
    LocalMux I__2639 (
            .O(N__18398),
            .I(N__18395));
    Span4Mux_v I__2638 (
            .O(N__18395),
            .I(N__18392));
    Odrv4 I__2637 (
            .O(N__18392),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__2636 (
            .O(N__18389),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    CascadeMux I__2635 (
            .O(N__18386),
            .I(N__18383));
    InMux I__2634 (
            .O(N__18383),
            .I(N__18380));
    LocalMux I__2633 (
            .O(N__18380),
            .I(N__18377));
    Span4Mux_v I__2632 (
            .O(N__18377),
            .I(N__18374));
    Odrv4 I__2631 (
            .O(N__18374),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__2630 (
            .O(N__18371),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    InMux I__2629 (
            .O(N__18368),
            .I(N__18365));
    LocalMux I__2628 (
            .O(N__18365),
            .I(N__18362));
    Span4Mux_v I__2627 (
            .O(N__18362),
            .I(N__18359));
    Odrv4 I__2626 (
            .O(N__18359),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__2625 (
            .O(N__18356),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    InMux I__2624 (
            .O(N__18353),
            .I(N__18350));
    LocalMux I__2623 (
            .O(N__18350),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    CascadeMux I__2622 (
            .O(N__18347),
            .I(N__18342));
    InMux I__2621 (
            .O(N__18346),
            .I(N__18339));
    InMux I__2620 (
            .O(N__18345),
            .I(N__18336));
    InMux I__2619 (
            .O(N__18342),
            .I(N__18333));
    LocalMux I__2618 (
            .O(N__18339),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__2617 (
            .O(N__18336),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__2616 (
            .O(N__18333),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__2615 (
            .O(N__18326),
            .I(N__18322));
    InMux I__2614 (
            .O(N__18325),
            .I(N__18319));
    LocalMux I__2613 (
            .O(N__18322),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__2612 (
            .O(N__18319),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__2611 (
            .O(N__18314),
            .I(N__18310));
    InMux I__2610 (
            .O(N__18313),
            .I(N__18307));
    LocalMux I__2609 (
            .O(N__18310),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__2608 (
            .O(N__18307),
            .I(\COUNTER.counterZ0Z_11 ));
    CascadeMux I__2607 (
            .O(N__18302),
            .I(N__18298));
    InMux I__2606 (
            .O(N__18301),
            .I(N__18295));
    InMux I__2605 (
            .O(N__18298),
            .I(N__18292));
    LocalMux I__2604 (
            .O(N__18295),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__2603 (
            .O(N__18292),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__2602 (
            .O(N__18287),
            .I(N__18283));
    InMux I__2601 (
            .O(N__18286),
            .I(N__18280));
    LocalMux I__2600 (
            .O(N__18283),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__2599 (
            .O(N__18280),
            .I(\COUNTER.counterZ0Z_9 ));
    InMux I__2598 (
            .O(N__18275),
            .I(N__18271));
    InMux I__2597 (
            .O(N__18274),
            .I(N__18268));
    LocalMux I__2596 (
            .O(N__18271),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__2595 (
            .O(N__18268),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__2594 (
            .O(N__18263),
            .I(N__18259));
    InMux I__2593 (
            .O(N__18262),
            .I(N__18256));
    LocalMux I__2592 (
            .O(N__18259),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__2591 (
            .O(N__18256),
            .I(\COUNTER.counterZ0Z_15 ));
    CascadeMux I__2590 (
            .O(N__18251),
            .I(N__18247));
    InMux I__2589 (
            .O(N__18250),
            .I(N__18244));
    InMux I__2588 (
            .O(N__18247),
            .I(N__18241));
    LocalMux I__2587 (
            .O(N__18244),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__2586 (
            .O(N__18241),
            .I(\COUNTER.counterZ0Z_13 ));
    InMux I__2585 (
            .O(N__18236),
            .I(N__18232));
    InMux I__2584 (
            .O(N__18235),
            .I(N__18229));
    LocalMux I__2583 (
            .O(N__18232),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__2582 (
            .O(N__18229),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__2581 (
            .O(N__18224),
            .I(N__18220));
    InMux I__2580 (
            .O(N__18223),
            .I(N__18217));
    LocalMux I__2579 (
            .O(N__18220),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__2578 (
            .O(N__18217),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__2577 (
            .O(N__18212),
            .I(N__18208));
    InMux I__2576 (
            .O(N__18211),
            .I(N__18205));
    LocalMux I__2575 (
            .O(N__18208),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__2574 (
            .O(N__18205),
            .I(\COUNTER.counterZ0Z_18 ));
    CascadeMux I__2573 (
            .O(N__18200),
            .I(N__18196));
    InMux I__2572 (
            .O(N__18199),
            .I(N__18193));
    InMux I__2571 (
            .O(N__18196),
            .I(N__18190));
    LocalMux I__2570 (
            .O(N__18193),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__2569 (
            .O(N__18190),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__2568 (
            .O(N__18185),
            .I(N__18181));
    InMux I__2567 (
            .O(N__18184),
            .I(N__18178));
    LocalMux I__2566 (
            .O(N__18181),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__2565 (
            .O(N__18178),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__2564 (
            .O(N__18173),
            .I(N__18169));
    InMux I__2563 (
            .O(N__18172),
            .I(N__18166));
    InMux I__2562 (
            .O(N__18169),
            .I(N__18163));
    LocalMux I__2561 (
            .O(N__18166),
            .I(N__18156));
    LocalMux I__2560 (
            .O(N__18163),
            .I(N__18156));
    InMux I__2559 (
            .O(N__18162),
            .I(N__18151));
    InMux I__2558 (
            .O(N__18161),
            .I(N__18151));
    Odrv4 I__2557 (
            .O(N__18156),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__2556 (
            .O(N__18151),
            .I(\COUNTER.counterZ0Z_0 ));
    CascadeMux I__2555 (
            .O(N__18146),
            .I(N__18143));
    InMux I__2554 (
            .O(N__18143),
            .I(N__18140));
    LocalMux I__2553 (
            .O(N__18140),
            .I(N__18136));
    InMux I__2552 (
            .O(N__18139),
            .I(N__18133));
    Span4Mux_v I__2551 (
            .O(N__18136),
            .I(N__18130));
    LocalMux I__2550 (
            .O(N__18133),
            .I(\PCH_PWRGD.N_670 ));
    Odrv4 I__2549 (
            .O(N__18130),
            .I(\PCH_PWRGD.N_670 ));
    InMux I__2548 (
            .O(N__18125),
            .I(N__18121));
    InMux I__2547 (
            .O(N__18124),
            .I(N__18118));
    LocalMux I__2546 (
            .O(N__18121),
            .I(N__18115));
    LocalMux I__2545 (
            .O(N__18118),
            .I(N__18112));
    Span4Mux_h I__2544 (
            .O(N__18115),
            .I(N__18109));
    Odrv12 I__2543 (
            .O(N__18112),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2542 (
            .O(N__18109),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__2541 (
            .O(N__18104),
            .I(N__18100));
    InMux I__2540 (
            .O(N__18103),
            .I(N__18097));
    LocalMux I__2539 (
            .O(N__18100),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__2538 (
            .O(N__18097),
            .I(\COUNTER.counterZ0Z_27 ));
    InMux I__2537 (
            .O(N__18092),
            .I(N__18088));
    InMux I__2536 (
            .O(N__18091),
            .I(N__18085));
    LocalMux I__2535 (
            .O(N__18088),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__2534 (
            .O(N__18085),
            .I(\COUNTER.counterZ0Z_26 ));
    CascadeMux I__2533 (
            .O(N__18080),
            .I(N__18076));
    InMux I__2532 (
            .O(N__18079),
            .I(N__18073));
    InMux I__2531 (
            .O(N__18076),
            .I(N__18070));
    LocalMux I__2530 (
            .O(N__18073),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__2529 (
            .O(N__18070),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__2528 (
            .O(N__18065),
            .I(N__18061));
    InMux I__2527 (
            .O(N__18064),
            .I(N__18058));
    LocalMux I__2526 (
            .O(N__18061),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__2525 (
            .O(N__18058),
            .I(\COUNTER.counterZ0Z_25 ));
    CascadeMux I__2524 (
            .O(N__18053),
            .I(\VPP_VDDQ.count_2_1_0_cascade_ ));
    CascadeMux I__2523 (
            .O(N__18050),
            .I(\VPP_VDDQ.count_2Z0Z_0_cascade_ ));
    InMux I__2522 (
            .O(N__18047),
            .I(N__18044));
    LocalMux I__2521 (
            .O(N__18044),
            .I(\VPP_VDDQ.count_2_0_0 ));
    InMux I__2520 (
            .O(N__18041),
            .I(N__18038));
    LocalMux I__2519 (
            .O(N__18038),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__2518 (
            .O(N__18035),
            .I(N__18030));
    InMux I__2517 (
            .O(N__18034),
            .I(N__18027));
    InMux I__2516 (
            .O(N__18033),
            .I(N__18024));
    LocalMux I__2515 (
            .O(N__18030),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2514 (
            .O(N__18027),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2513 (
            .O(N__18024),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__2512 (
            .O(N__18017),
            .I(N__18014));
    LocalMux I__2511 (
            .O(N__18014),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__2510 (
            .O(N__18011),
            .I(N__18008));
    LocalMux I__2509 (
            .O(N__18008),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    CascadeMux I__2508 (
            .O(N__18005),
            .I(N__18000));
    CascadeMux I__2507 (
            .O(N__18004),
            .I(N__17997));
    InMux I__2506 (
            .O(N__18003),
            .I(N__17994));
    InMux I__2505 (
            .O(N__18000),
            .I(N__17989));
    InMux I__2504 (
            .O(N__17997),
            .I(N__17989));
    LocalMux I__2503 (
            .O(N__17994),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__2502 (
            .O(N__17989),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__2501 (
            .O(N__17984),
            .I(N__17981));
    LocalMux I__2500 (
            .O(N__17981),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    CascadeMux I__2499 (
            .O(N__17978),
            .I(N__17974));
    InMux I__2498 (
            .O(N__17977),
            .I(N__17970));
    InMux I__2497 (
            .O(N__17974),
            .I(N__17965));
    InMux I__2496 (
            .O(N__17973),
            .I(N__17965));
    LocalMux I__2495 (
            .O(N__17970),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__2494 (
            .O(N__17965),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__2493 (
            .O(N__17960),
            .I(N__17956));
    InMux I__2492 (
            .O(N__17959),
            .I(N__17953));
    LocalMux I__2491 (
            .O(N__17956),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__2490 (
            .O(N__17953),
            .I(\COUNTER.counterZ0Z_7 ));
    CascadeMux I__2489 (
            .O(N__17948),
            .I(N__17944));
    InMux I__2488 (
            .O(N__17947),
            .I(N__17940));
    InMux I__2487 (
            .O(N__17944),
            .I(N__17935));
    InMux I__2486 (
            .O(N__17943),
            .I(N__17935));
    LocalMux I__2485 (
            .O(N__17940),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__2484 (
            .O(N__17935),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__2483 (
            .O(N__17930),
            .I(N__17925));
    InMux I__2482 (
            .O(N__17929),
            .I(N__17920));
    InMux I__2481 (
            .O(N__17928),
            .I(N__17920));
    LocalMux I__2480 (
            .O(N__17925),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__2479 (
            .O(N__17920),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__2478 (
            .O(N__17915),
            .I(N__17912));
    LocalMux I__2477 (
            .O(N__17912),
            .I(N__17908));
    InMux I__2476 (
            .O(N__17911),
            .I(N__17905));
    Odrv4 I__2475 (
            .O(N__17908),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    LocalMux I__2474 (
            .O(N__17905),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    InMux I__2473 (
            .O(N__17900),
            .I(N__17896));
    InMux I__2472 (
            .O(N__17899),
            .I(N__17893));
    LocalMux I__2471 (
            .O(N__17896),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    LocalMux I__2470 (
            .O(N__17893),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    InMux I__2469 (
            .O(N__17888),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__2468 (
            .O(N__17885),
            .I(N__17881));
    InMux I__2467 (
            .O(N__17884),
            .I(N__17878));
    LocalMux I__2466 (
            .O(N__17881),
            .I(N__17873));
    LocalMux I__2465 (
            .O(N__17878),
            .I(N__17873));
    Odrv4 I__2464 (
            .O(N__17873),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    InMux I__2463 (
            .O(N__17870),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    InMux I__2462 (
            .O(N__17867),
            .I(N__17861));
    InMux I__2461 (
            .O(N__17866),
            .I(N__17861));
    LocalMux I__2460 (
            .O(N__17861),
            .I(N__17858));
    Odrv4 I__2459 (
            .O(N__17858),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ));
    CascadeMux I__2458 (
            .O(N__17855),
            .I(N__17852));
    InMux I__2457 (
            .O(N__17852),
            .I(N__17848));
    InMux I__2456 (
            .O(N__17851),
            .I(N__17845));
    LocalMux I__2455 (
            .O(N__17848),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    LocalMux I__2454 (
            .O(N__17845),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    InMux I__2453 (
            .O(N__17840),
            .I(N__17837));
    LocalMux I__2452 (
            .O(N__17837),
            .I(\VPP_VDDQ.count_2_1_13 ));
    InMux I__2451 (
            .O(N__17834),
            .I(N__17830));
    InMux I__2450 (
            .O(N__17833),
            .I(N__17827));
    LocalMux I__2449 (
            .O(N__17830),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    LocalMux I__2448 (
            .O(N__17827),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    CascadeMux I__2447 (
            .O(N__17822),
            .I(N__17819));
    InMux I__2446 (
            .O(N__17819),
            .I(N__17816));
    LocalMux I__2445 (
            .O(N__17816),
            .I(\VPP_VDDQ.un9_clk_100khz_10 ));
    InMux I__2444 (
            .O(N__17813),
            .I(N__17809));
    InMux I__2443 (
            .O(N__17812),
            .I(N__17806));
    LocalMux I__2442 (
            .O(N__17809),
            .I(N__17801));
    LocalMux I__2441 (
            .O(N__17806),
            .I(N__17801));
    Odrv4 I__2440 (
            .O(N__17801),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    InMux I__2439 (
            .O(N__17798),
            .I(N__17795));
    LocalMux I__2438 (
            .O(N__17795),
            .I(\VPP_VDDQ.un9_clk_100khz_7 ));
    InMux I__2437 (
            .O(N__17792),
            .I(N__17789));
    LocalMux I__2436 (
            .O(N__17789),
            .I(\VPP_VDDQ.count_2_1_7 ));
    CascadeMux I__2435 (
            .O(N__17786),
            .I(\VPP_VDDQ.count_2_1_7_cascade_ ));
    InMux I__2434 (
            .O(N__17783),
            .I(N__17780));
    LocalMux I__2433 (
            .O(N__17780),
            .I(N__17777));
    Odrv4 I__2432 (
            .O(N__17777),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    InMux I__2431 (
            .O(N__17774),
            .I(N__17768));
    InMux I__2430 (
            .O(N__17773),
            .I(N__17768));
    LocalMux I__2429 (
            .O(N__17768),
            .I(N__17765));
    Odrv4 I__2428 (
            .O(N__17765),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ));
    InMux I__2427 (
            .O(N__17762),
            .I(N__17756));
    InMux I__2426 (
            .O(N__17761),
            .I(N__17756));
    LocalMux I__2425 (
            .O(N__17756),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    InMux I__2424 (
            .O(N__17753),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    InMux I__2423 (
            .O(N__17750),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__2422 (
            .O(N__17747),
            .I(N__17743));
    InMux I__2421 (
            .O(N__17746),
            .I(N__17740));
    LocalMux I__2420 (
            .O(N__17743),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    LocalMux I__2419 (
            .O(N__17740),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    CascadeMux I__2418 (
            .O(N__17735),
            .I(N__17731));
    CascadeMux I__2417 (
            .O(N__17734),
            .I(N__17728));
    InMux I__2416 (
            .O(N__17731),
            .I(N__17723));
    InMux I__2415 (
            .O(N__17728),
            .I(N__17723));
    LocalMux I__2414 (
            .O(N__17723),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ));
    InMux I__2413 (
            .O(N__17720),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    InMux I__2412 (
            .O(N__17717),
            .I(N__17711));
    InMux I__2411 (
            .O(N__17716),
            .I(N__17711));
    LocalMux I__2410 (
            .O(N__17711),
            .I(N__17708));
    Odrv4 I__2409 (
            .O(N__17708),
            .I(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ));
    InMux I__2408 (
            .O(N__17705),
            .I(bfn_5_3_0_));
    CascadeMux I__2407 (
            .O(N__17702),
            .I(N__17699));
    InMux I__2406 (
            .O(N__17699),
            .I(N__17696));
    LocalMux I__2405 (
            .O(N__17696),
            .I(N__17692));
    InMux I__2404 (
            .O(N__17695),
            .I(N__17689));
    Odrv4 I__2403 (
            .O(N__17692),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ));
    LocalMux I__2402 (
            .O(N__17689),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ));
    InMux I__2401 (
            .O(N__17684),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__2400 (
            .O(N__17681),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__2399 (
            .O(N__17678),
            .I(N__17675));
    LocalMux I__2398 (
            .O(N__17675),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    InMux I__2397 (
            .O(N__17672),
            .I(N__17666));
    InMux I__2396 (
            .O(N__17671),
            .I(N__17666));
    LocalMux I__2395 (
            .O(N__17666),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ));
    InMux I__2394 (
            .O(N__17663),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    InMux I__2393 (
            .O(N__17660),
            .I(N__17656));
    InMux I__2392 (
            .O(N__17659),
            .I(N__17653));
    LocalMux I__2391 (
            .O(N__17656),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    LocalMux I__2390 (
            .O(N__17653),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    InMux I__2389 (
            .O(N__17648),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    CascadeMux I__2388 (
            .O(N__17645),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ));
    InMux I__2387 (
            .O(N__17642),
            .I(N__17639));
    LocalMux I__2386 (
            .O(N__17639),
            .I(\VPP_VDDQ.count_2_0_15 ));
    InMux I__2385 (
            .O(N__17636),
            .I(N__17633));
    LocalMux I__2384 (
            .O(N__17633),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    InMux I__2383 (
            .O(N__17630),
            .I(N__17624));
    InMux I__2382 (
            .O(N__17629),
            .I(N__17624));
    LocalMux I__2381 (
            .O(N__17624),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ));
    InMux I__2380 (
            .O(N__17621),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    InMux I__2379 (
            .O(N__17618),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__2378 (
            .O(N__17615),
            .I(N__17609));
    InMux I__2377 (
            .O(N__17614),
            .I(N__17609));
    LocalMux I__2376 (
            .O(N__17609),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ));
    InMux I__2375 (
            .O(N__17606),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    InMux I__2374 (
            .O(N__17603),
            .I(N__17600));
    LocalMux I__2373 (
            .O(N__17600),
            .I(N__17596));
    InMux I__2372 (
            .O(N__17599),
            .I(N__17593));
    Odrv4 I__2371 (
            .O(N__17596),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    LocalMux I__2370 (
            .O(N__17593),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    CascadeMux I__2369 (
            .O(N__17588),
            .I(N__17585));
    InMux I__2368 (
            .O(N__17585),
            .I(N__17579));
    InMux I__2367 (
            .O(N__17584),
            .I(N__17579));
    LocalMux I__2366 (
            .O(N__17579),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ));
    InMux I__2365 (
            .O(N__17576),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    InMux I__2364 (
            .O(N__17573),
            .I(N__17570));
    LocalMux I__2363 (
            .O(N__17570),
            .I(\POWERLED.count_0_14 ));
    CascadeMux I__2362 (
            .O(N__17567),
            .I(\POWERLED.countZ0Z_14_cascade_ ));
    InMux I__2361 (
            .O(N__17564),
            .I(N__17561));
    LocalMux I__2360 (
            .O(N__17561),
            .I(N__17558));
    Span4Mux_s3_h I__2359 (
            .O(N__17558),
            .I(N__17555));
    Odrv4 I__2358 (
            .O(N__17555),
            .I(\POWERLED.un79_clk_100khzlto15_5 ));
    InMux I__2357 (
            .O(N__17552),
            .I(N__17549));
    LocalMux I__2356 (
            .O(N__17549),
            .I(N__17546));
    Span4Mux_v I__2355 (
            .O(N__17546),
            .I(N__17543));
    Odrv4 I__2354 (
            .O(N__17543),
            .I(\POWERLED.g1_i_o4_4 ));
    InMux I__2353 (
            .O(N__17540),
            .I(N__17537));
    LocalMux I__2352 (
            .O(N__17537),
            .I(\POWERLED.count_0_15 ));
    InMux I__2351 (
            .O(N__17534),
            .I(N__17531));
    LocalMux I__2350 (
            .O(N__17531),
            .I(\VPP_VDDQ.count_2_0_2 ));
    CascadeMux I__2349 (
            .O(N__17528),
            .I(\VPP_VDDQ.count_2_1_2_cascade_ ));
    CascadeMux I__2348 (
            .O(N__17525),
            .I(\VPP_VDDQ.count_2Z0Z_2_cascade_ ));
    CascadeMux I__2347 (
            .O(N__17522),
            .I(\POWERLED.count_1_0_cascade_ ));
    CascadeMux I__2346 (
            .O(N__17519),
            .I(\POWERLED.countZ0Z_0_cascade_ ));
    InMux I__2345 (
            .O(N__17516),
            .I(N__17513));
    LocalMux I__2344 (
            .O(N__17513),
            .I(\POWERLED.count_1_1 ));
    CascadeMux I__2343 (
            .O(N__17510),
            .I(\POWERLED.count_1_1_cascade_ ));
    CascadeMux I__2342 (
            .O(N__17507),
            .I(\POWERLED.un1_count_axb_1_cascade_ ));
    InMux I__2341 (
            .O(N__17504),
            .I(N__17498));
    InMux I__2340 (
            .O(N__17503),
            .I(N__17498));
    LocalMux I__2339 (
            .O(N__17498),
            .I(\POWERLED.countZ0Z_1 ));
    InMux I__2338 (
            .O(N__17495),
            .I(N__17492));
    LocalMux I__2337 (
            .O(N__17492),
            .I(\POWERLED.count_0_0 ));
    InMux I__2336 (
            .O(N__17489),
            .I(N__17486));
    LocalMux I__2335 (
            .O(N__17486),
            .I(\POWERLED.count_0_11 ));
    CascadeMux I__2334 (
            .O(N__17483),
            .I(N__17479));
    InMux I__2333 (
            .O(N__17482),
            .I(N__17475));
    InMux I__2332 (
            .O(N__17479),
            .I(N__17470));
    InMux I__2331 (
            .O(N__17478),
            .I(N__17470));
    LocalMux I__2330 (
            .O(N__17475),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__2329 (
            .O(N__17470),
            .I(\POWERLED.countZ0Z_2 ));
    CascadeMux I__2328 (
            .O(N__17465),
            .I(\POWERLED.un79_clk_100khzlto4_0_cascade_ ));
    InMux I__2327 (
            .O(N__17462),
            .I(N__17458));
    InMux I__2326 (
            .O(N__17461),
            .I(N__17455));
    LocalMux I__2325 (
            .O(N__17458),
            .I(N__17452));
    LocalMux I__2324 (
            .O(N__17455),
            .I(N__17449));
    Odrv4 I__2323 (
            .O(N__17452),
            .I(\POWERLED.un79_clk_100khzlt6 ));
    Odrv4 I__2322 (
            .O(N__17449),
            .I(\POWERLED.un79_clk_100khzlt6 ));
    CascadeMux I__2321 (
            .O(N__17444),
            .I(N__17440));
    InMux I__2320 (
            .O(N__17443),
            .I(N__17437));
    InMux I__2319 (
            .O(N__17440),
            .I(N__17434));
    LocalMux I__2318 (
            .O(N__17437),
            .I(N__17431));
    LocalMux I__2317 (
            .O(N__17434),
            .I(N__17428));
    Odrv12 I__2316 (
            .O(N__17431),
            .I(\POWERLED.mult1_un138_sum_i_8 ));
    Odrv4 I__2315 (
            .O(N__17428),
            .I(\POWERLED.mult1_un138_sum_i_8 ));
    InMux I__2314 (
            .O(N__17423),
            .I(N__17414));
    InMux I__2313 (
            .O(N__17422),
            .I(N__17414));
    InMux I__2312 (
            .O(N__17421),
            .I(N__17414));
    LocalMux I__2311 (
            .O(N__17414),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__2310 (
            .O(N__17411),
            .I(N__17408));
    LocalMux I__2309 (
            .O(N__17408),
            .I(N__17405));
    Span4Mux_v I__2308 (
            .O(N__17405),
            .I(N__17402));
    Odrv4 I__2307 (
            .O(N__17402),
            .I(\POWERLED.count_RNIJEFE_0Z0Z_4 ));
    InMux I__2306 (
            .O(N__17399),
            .I(N__17396));
    LocalMux I__2305 (
            .O(N__17396),
            .I(N__17392));
    CascadeMux I__2304 (
            .O(N__17395),
            .I(N__17389));
    Span4Mux_v I__2303 (
            .O(N__17392),
            .I(N__17386));
    InMux I__2302 (
            .O(N__17389),
            .I(N__17383));
    Odrv4 I__2301 (
            .O(N__17386),
            .I(\POWERLED.mult1_un159_sum_i_8 ));
    LocalMux I__2300 (
            .O(N__17383),
            .I(\POWERLED.mult1_un159_sum_i_8 ));
    InMux I__2299 (
            .O(N__17378),
            .I(N__17375));
    LocalMux I__2298 (
            .O(N__17375),
            .I(N__17372));
    Span4Mux_v I__2297 (
            .O(N__17372),
            .I(N__17369));
    Odrv4 I__2296 (
            .O(N__17369),
            .I(\POWERLED.count_RNIUGSJ_0Z0Z_1 ));
    CascadeMux I__2295 (
            .O(N__17366),
            .I(N__17362));
    InMux I__2294 (
            .O(N__17365),
            .I(N__17351));
    InMux I__2293 (
            .O(N__17362),
            .I(N__17351));
    InMux I__2292 (
            .O(N__17361),
            .I(N__17351));
    InMux I__2291 (
            .O(N__17360),
            .I(N__17351));
    LocalMux I__2290 (
            .O(N__17351),
            .I(N__17347));
    InMux I__2289 (
            .O(N__17350),
            .I(N__17344));
    Span4Mux_h I__2288 (
            .O(N__17347),
            .I(N__17341));
    LocalMux I__2287 (
            .O(N__17344),
            .I(N__17338));
    Odrv4 I__2286 (
            .O(N__17341),
            .I(\POWERLED.N_660 ));
    Odrv12 I__2285 (
            .O(N__17338),
            .I(\POWERLED.N_660 ));
    CascadeMux I__2284 (
            .O(N__17333),
            .I(\POWERLED.count_0_sqmuxa_cascade_ ));
    CascadeMux I__2283 (
            .O(N__17330),
            .I(N__17327));
    InMux I__2282 (
            .O(N__17327),
            .I(N__17324));
    LocalMux I__2281 (
            .O(N__17324),
            .I(\POWERLED.mult1_un103_sum_i_8 ));
    InMux I__2280 (
            .O(N__17321),
            .I(N__17318));
    LocalMux I__2279 (
            .O(N__17318),
            .I(N__17314));
    CascadeMux I__2278 (
            .O(N__17317),
            .I(N__17310));
    Span4Mux_v I__2277 (
            .O(N__17314),
            .I(N__17305));
    InMux I__2276 (
            .O(N__17313),
            .I(N__17298));
    InMux I__2275 (
            .O(N__17310),
            .I(N__17298));
    InMux I__2274 (
            .O(N__17309),
            .I(N__17298));
    InMux I__2273 (
            .O(N__17308),
            .I(N__17295));
    Odrv4 I__2272 (
            .O(N__17305),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2271 (
            .O(N__17298),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2270 (
            .O(N__17295),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    InMux I__2269 (
            .O(N__17288),
            .I(N__17285));
    LocalMux I__2268 (
            .O(N__17285),
            .I(\POWERLED.mult1_un96_sum_i_8 ));
    CascadeMux I__2267 (
            .O(N__17282),
            .I(N__17279));
    InMux I__2266 (
            .O(N__17279),
            .I(N__17276));
    LocalMux I__2265 (
            .O(N__17276),
            .I(N__17273));
    Odrv12 I__2264 (
            .O(N__17273),
            .I(\POWERLED.mult1_un110_sum_i ));
    CascadeMux I__2263 (
            .O(N__17270),
            .I(\POWERLED.N_437_cascade_ ));
    InMux I__2262 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__2261 (
            .O(N__17264),
            .I(N__17260));
    InMux I__2260 (
            .O(N__17263),
            .I(N__17257));
    Span4Mux_s3_h I__2259 (
            .O(N__17260),
            .I(N__17254));
    LocalMux I__2258 (
            .O(N__17257),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__2257 (
            .O(N__17254),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    CascadeMux I__2256 (
            .O(N__17249),
            .I(N__17246));
    InMux I__2255 (
            .O(N__17246),
            .I(N__17240));
    InMux I__2254 (
            .O(N__17245),
            .I(N__17240));
    LocalMux I__2253 (
            .O(N__17240),
            .I(N__17237));
    Span4Mux_v I__2252 (
            .O(N__17237),
            .I(N__17234));
    Span4Mux_s1_h I__2251 (
            .O(N__17234),
            .I(N__17229));
    InMux I__2250 (
            .O(N__17233),
            .I(N__17224));
    InMux I__2249 (
            .O(N__17232),
            .I(N__17224));
    Odrv4 I__2248 (
            .O(N__17229),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    LocalMux I__2247 (
            .O(N__17224),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    CascadeMux I__2246 (
            .O(N__17219),
            .I(\POWERLED.curr_stateZ0Z_0_cascade_ ));
    InMux I__2245 (
            .O(N__17216),
            .I(N__17213));
    LocalMux I__2244 (
            .O(N__17213),
            .I(\POWERLED.curr_state_1_0 ));
    CascadeMux I__2243 (
            .O(N__17210),
            .I(N__17207));
    InMux I__2242 (
            .O(N__17207),
            .I(N__17204));
    LocalMux I__2241 (
            .O(N__17204),
            .I(\POWERLED.count_0_3 ));
    InMux I__2240 (
            .O(N__17201),
            .I(N__17197));
    CascadeMux I__2239 (
            .O(N__17200),
            .I(N__17194));
    LocalMux I__2238 (
            .O(N__17197),
            .I(N__17191));
    InMux I__2237 (
            .O(N__17194),
            .I(N__17188));
    Odrv12 I__2236 (
            .O(N__17191),
            .I(\POWERLED.mult1_un152_sum_i_8 ));
    LocalMux I__2235 (
            .O(N__17188),
            .I(\POWERLED.mult1_un152_sum_i_8 ));
    InMux I__2234 (
            .O(N__17183),
            .I(N__17180));
    LocalMux I__2233 (
            .O(N__17180),
            .I(N__17177));
    Span4Mux_v I__2232 (
            .O(N__17177),
            .I(N__17174));
    Odrv4 I__2231 (
            .O(N__17174),
            .I(\POWERLED.count_RNIAKSS_0Z0Z_2 ));
    InMux I__2230 (
            .O(N__17171),
            .I(N__17168));
    LocalMux I__2229 (
            .O(N__17168),
            .I(\POWERLED.N_4851_i ));
    InMux I__2228 (
            .O(N__17165),
            .I(N__17162));
    LocalMux I__2227 (
            .O(N__17162),
            .I(\POWERLED.N_4855_i ));
    InMux I__2226 (
            .O(N__17159),
            .I(N__17156));
    LocalMux I__2225 (
            .O(N__17156),
            .I(\POWERLED.N_4856_i ));
    InMux I__2224 (
            .O(N__17153),
            .I(bfn_4_11_0_));
    CascadeMux I__2223 (
            .O(N__17150),
            .I(N__17147));
    InMux I__2222 (
            .O(N__17147),
            .I(N__17144));
    LocalMux I__2221 (
            .O(N__17144),
            .I(N__17141));
    Odrv4 I__2220 (
            .O(N__17141),
            .I(\POWERLED.mult1_un117_sum_i_8 ));
    InMux I__2219 (
            .O(N__17138),
            .I(N__17134));
    CascadeMux I__2218 (
            .O(N__17137),
            .I(N__17130));
    LocalMux I__2217 (
            .O(N__17134),
            .I(N__17125));
    InMux I__2216 (
            .O(N__17133),
            .I(N__17118));
    InMux I__2215 (
            .O(N__17130),
            .I(N__17118));
    InMux I__2214 (
            .O(N__17129),
            .I(N__17118));
    InMux I__2213 (
            .O(N__17128),
            .I(N__17115));
    Odrv12 I__2212 (
            .O(N__17125),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2211 (
            .O(N__17118),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2210 (
            .O(N__17115),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__2209 (
            .O(N__17108),
            .I(N__17105));
    InMux I__2208 (
            .O(N__17105),
            .I(N__17102));
    LocalMux I__2207 (
            .O(N__17102),
            .I(\POWERLED.mult1_un110_sum_i_8 ));
    CascadeMux I__2206 (
            .O(N__17099),
            .I(N__17096));
    InMux I__2205 (
            .O(N__17096),
            .I(N__17093));
    LocalMux I__2204 (
            .O(N__17093),
            .I(\POWERLED.mult1_un89_sum_i_8 ));
    InMux I__2203 (
            .O(N__17090),
            .I(N__17087));
    LocalMux I__2202 (
            .O(N__17087),
            .I(N__17083));
    CascadeMux I__2201 (
            .O(N__17086),
            .I(N__17080));
    Span4Mux_h I__2200 (
            .O(N__17083),
            .I(N__17074));
    InMux I__2199 (
            .O(N__17080),
            .I(N__17067));
    InMux I__2198 (
            .O(N__17079),
            .I(N__17067));
    InMux I__2197 (
            .O(N__17078),
            .I(N__17067));
    InMux I__2196 (
            .O(N__17077),
            .I(N__17064));
    Odrv4 I__2195 (
            .O(N__17074),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__2194 (
            .O(N__17067),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__2193 (
            .O(N__17064),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    InMux I__2192 (
            .O(N__17057),
            .I(N__17054));
    LocalMux I__2191 (
            .O(N__17054),
            .I(N__17050));
    CascadeMux I__2190 (
            .O(N__17053),
            .I(N__17047));
    Span4Mux_h I__2189 (
            .O(N__17050),
            .I(N__17041));
    InMux I__2188 (
            .O(N__17047),
            .I(N__17034));
    InMux I__2187 (
            .O(N__17046),
            .I(N__17034));
    InMux I__2186 (
            .O(N__17045),
            .I(N__17034));
    InMux I__2185 (
            .O(N__17044),
            .I(N__17031));
    Odrv4 I__2184 (
            .O(N__17041),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2183 (
            .O(N__17034),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2182 (
            .O(N__17031),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    InMux I__2181 (
            .O(N__17024),
            .I(N__17021));
    LocalMux I__2180 (
            .O(N__17021),
            .I(N__17018));
    Span4Mux_h I__2179 (
            .O(N__17018),
            .I(N__17015));
    Odrv4 I__2178 (
            .O(N__17015),
            .I(\POWERLED.count_RNIGTVS_1Z0Z_5 ));
    InMux I__2177 (
            .O(N__17012),
            .I(N__17009));
    LocalMux I__2176 (
            .O(N__17009),
            .I(N__17005));
    CascadeMux I__2175 (
            .O(N__17008),
            .I(N__17002));
    Span4Mux_v I__2174 (
            .O(N__17005),
            .I(N__16999));
    InMux I__2173 (
            .O(N__17002),
            .I(N__16996));
    Odrv4 I__2172 (
            .O(N__16999),
            .I(\POWERLED.mult1_un131_sum_i_8 ));
    LocalMux I__2171 (
            .O(N__16996),
            .I(\POWERLED.mult1_un131_sum_i_8 ));
    CascadeMux I__2170 (
            .O(N__16991),
            .I(N__16988));
    InMux I__2169 (
            .O(N__16988),
            .I(N__16985));
    LocalMux I__2168 (
            .O(N__16985),
            .I(\POWERLED.count_i_6 ));
    InMux I__2167 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__2166 (
            .O(N__16979),
            .I(\POWERLED.N_4841_i ));
    InMux I__2165 (
            .O(N__16976),
            .I(N__16973));
    LocalMux I__2164 (
            .O(N__16973),
            .I(\POWERLED.count_i_8 ));
    InMux I__2163 (
            .O(N__16970),
            .I(N__16967));
    LocalMux I__2162 (
            .O(N__16967),
            .I(\POWERLED.N_4849_i ));
    CascadeMux I__2161 (
            .O(N__16964),
            .I(N__16961));
    InMux I__2160 (
            .O(N__16961),
            .I(N__16958));
    LocalMux I__2159 (
            .O(N__16958),
            .I(\POWERLED.count_i_10 ));
    InMux I__2158 (
            .O(N__16955),
            .I(N__16952));
    LocalMux I__2157 (
            .O(N__16952),
            .I(\POWERLED.count_i_11 ));
    InMux I__2156 (
            .O(N__16949),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__2155 (
            .O(N__16946),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__2154 (
            .O(N__16943),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__2153 (
            .O(N__16940),
            .I(\COUNTER.counter_1_cry_30 ));
    CascadeMux I__2152 (
            .O(N__16937),
            .I(N__16934));
    InMux I__2151 (
            .O(N__16934),
            .I(N__16928));
    InMux I__2150 (
            .O(N__16933),
            .I(N__16928));
    LocalMux I__2149 (
            .O(N__16928),
            .I(\COUNTER.counterZ0Z_30 ));
    InMux I__2148 (
            .O(N__16925),
            .I(N__16919));
    InMux I__2147 (
            .O(N__16924),
            .I(N__16919));
    LocalMux I__2146 (
            .O(N__16919),
            .I(\COUNTER.counterZ0Z_31 ));
    CascadeMux I__2145 (
            .O(N__16916),
            .I(N__16912));
    InMux I__2144 (
            .O(N__16915),
            .I(N__16907));
    InMux I__2143 (
            .O(N__16912),
            .I(N__16907));
    LocalMux I__2142 (
            .O(N__16907),
            .I(\COUNTER.counterZ0Z_29 ));
    InMux I__2141 (
            .O(N__16904),
            .I(N__16898));
    InMux I__2140 (
            .O(N__16903),
            .I(N__16898));
    LocalMux I__2139 (
            .O(N__16898),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__2138 (
            .O(N__16895),
            .I(N__16892));
    LocalMux I__2137 (
            .O(N__16892),
            .I(\POWERLED.N_4842_i ));
    CascadeMux I__2136 (
            .O(N__16889),
            .I(N__16886));
    InMux I__2135 (
            .O(N__16886),
            .I(N__16883));
    LocalMux I__2134 (
            .O(N__16883),
            .I(\POWERLED.count_i_3 ));
    InMux I__2133 (
            .O(N__16880),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__2132 (
            .O(N__16877),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__2131 (
            .O(N__16874),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__2130 (
            .O(N__16871),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__2129 (
            .O(N__16868),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__2128 (
            .O(N__16865),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__2127 (
            .O(N__16862),
            .I(bfn_4_8_0_));
    InMux I__2126 (
            .O(N__16859),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__2125 (
            .O(N__16856),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__2124 (
            .O(N__16853),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__2123 (
            .O(N__16850),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__2122 (
            .O(N__16847),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__2121 (
            .O(N__16844),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__2120 (
            .O(N__16841),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__2119 (
            .O(N__16838),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__2118 (
            .O(N__16835),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__2117 (
            .O(N__16832),
            .I(bfn_4_7_0_));
    InMux I__2116 (
            .O(N__16829),
            .I(\COUNTER.counter_1_cry_17 ));
    CascadeMux I__2115 (
            .O(N__16826),
            .I(\VPP_VDDQ.count_2_1_10_cascade_ ));
    InMux I__2114 (
            .O(N__16823),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__2113 (
            .O(N__16820),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__2112 (
            .O(N__16817),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__2111 (
            .O(N__16814),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__2110 (
            .O(N__16811),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__2109 (
            .O(N__16808),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__2108 (
            .O(N__16805),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__2107 (
            .O(N__16802),
            .I(bfn_4_6_0_));
    CascadeMux I__2106 (
            .O(N__16799),
            .I(\VPP_VDDQ.count_2Z0Z_12_cascade_ ));
    InMux I__2105 (
            .O(N__16796),
            .I(N__16793));
    LocalMux I__2104 (
            .O(N__16793),
            .I(\VPP_VDDQ.count_2_0_12 ));
    InMux I__2103 (
            .O(N__16790),
            .I(N__16787));
    LocalMux I__2102 (
            .O(N__16787),
            .I(\VPP_VDDQ.count_2_0_13 ));
    InMux I__2101 (
            .O(N__16784),
            .I(N__16781));
    LocalMux I__2100 (
            .O(N__16781),
            .I(\VPP_VDDQ.count_2_0_14 ));
    InMux I__2099 (
            .O(N__16778),
            .I(N__16775));
    LocalMux I__2098 (
            .O(N__16775),
            .I(N__16772));
    Span12Mux_s10_h I__2097 (
            .O(N__16772),
            .I(N__16765));
    InMux I__2096 (
            .O(N__16771),
            .I(N__16756));
    InMux I__2095 (
            .O(N__16770),
            .I(N__16756));
    InMux I__2094 (
            .O(N__16769),
            .I(N__16756));
    InMux I__2093 (
            .O(N__16768),
            .I(N__16756));
    Odrv12 I__2092 (
            .O(N__16765),
            .I(VPP_VDDQ_curr_state_0));
    LocalMux I__2091 (
            .O(N__16756),
            .I(VPP_VDDQ_curr_state_0));
    InMux I__2090 (
            .O(N__16751),
            .I(N__16745));
    InMux I__2089 (
            .O(N__16750),
            .I(N__16745));
    LocalMux I__2088 (
            .O(N__16745),
            .I(N__16742));
    Span4Mux_h I__2087 (
            .O(N__16742),
            .I(N__16738));
    CascadeMux I__2086 (
            .O(N__16741),
            .I(N__16735));
    Span4Mux_v I__2085 (
            .O(N__16738),
            .I(N__16728));
    InMux I__2084 (
            .O(N__16735),
            .I(N__16717));
    InMux I__2083 (
            .O(N__16734),
            .I(N__16717));
    InMux I__2082 (
            .O(N__16733),
            .I(N__16717));
    InMux I__2081 (
            .O(N__16732),
            .I(N__16717));
    InMux I__2080 (
            .O(N__16731),
            .I(N__16717));
    Odrv4 I__2079 (
            .O(N__16728),
            .I(VPP_VDDQ_curr_state_1));
    LocalMux I__2078 (
            .O(N__16717),
            .I(VPP_VDDQ_curr_state_1));
    CascadeMux I__2077 (
            .O(N__16712),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ));
    InMux I__2076 (
            .O(N__16709),
            .I(N__16706));
    LocalMux I__2075 (
            .O(N__16706),
            .I(N__16703));
    Span4Mux_h I__2074 (
            .O(N__16703),
            .I(N__16699));
    InMux I__2073 (
            .O(N__16702),
            .I(N__16694));
    Span4Mux_v I__2072 (
            .O(N__16699),
            .I(N__16691));
    InMux I__2071 (
            .O(N__16698),
            .I(N__16686));
    InMux I__2070 (
            .O(N__16697),
            .I(N__16686));
    LocalMux I__2069 (
            .O(N__16694),
            .I(N_626));
    Odrv4 I__2068 (
            .O(N__16691),
            .I(N_626));
    LocalMux I__2067 (
            .O(N__16686),
            .I(N_626));
    InMux I__2066 (
            .O(N__16679),
            .I(N__16673));
    InMux I__2065 (
            .O(N__16678),
            .I(N__16670));
    InMux I__2064 (
            .O(N__16677),
            .I(N__16667));
    CascadeMux I__2063 (
            .O(N__16676),
            .I(N__16664));
    LocalMux I__2062 (
            .O(N__16673),
            .I(N__16661));
    LocalMux I__2061 (
            .O(N__16670),
            .I(N__16658));
    LocalMux I__2060 (
            .O(N__16667),
            .I(N__16655));
    InMux I__2059 (
            .O(N__16664),
            .I(N__16652));
    Span4Mux_h I__2058 (
            .O(N__16661),
            .I(N__16649));
    Span12Mux_s1_h I__2057 (
            .O(N__16658),
            .I(N__16646));
    Odrv4 I__2056 (
            .O(N__16655),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    LocalMux I__2055 (
            .O(N__16652),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    Odrv4 I__2054 (
            .O(N__16649),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    Odrv12 I__2053 (
            .O(N__16646),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    InMux I__2052 (
            .O(N__16637),
            .I(N__16633));
    InMux I__2051 (
            .O(N__16636),
            .I(N__16630));
    LocalMux I__2050 (
            .O(N__16633),
            .I(N__16627));
    LocalMux I__2049 (
            .O(N__16630),
            .I(N__16624));
    Span4Mux_h I__2048 (
            .O(N__16627),
            .I(N__16621));
    Span12Mux_s1_v I__2047 (
            .O(N__16624),
            .I(N__16618));
    Odrv4 I__2046 (
            .O(N__16621),
            .I(\PCH_PWRGD.N_38_f0 ));
    Odrv12 I__2045 (
            .O(N__16618),
            .I(\PCH_PWRGD.N_38_f0 ));
    InMux I__2044 (
            .O(N__16613),
            .I(N__16610));
    LocalMux I__2043 (
            .O(N__16610),
            .I(N__16606));
    InMux I__2042 (
            .O(N__16609),
            .I(N__16603));
    Span4Mux_s3_v I__2041 (
            .O(N__16606),
            .I(N__16600));
    LocalMux I__2040 (
            .O(N__16603),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    Odrv4 I__2039 (
            .O(N__16600),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    InMux I__2038 (
            .O(N__16595),
            .I(N__16592));
    LocalMux I__2037 (
            .O(N__16592),
            .I(N__16589));
    Odrv4 I__2036 (
            .O(N__16589),
            .I(\VPP_VDDQ.count_2_0_10 ));
    CascadeMux I__2035 (
            .O(N__16586),
            .I(\VPP_VDDQ.count_2_1_14_cascade_ ));
    CascadeMux I__2034 (
            .O(N__16583),
            .I(\VPP_VDDQ.count_2_1_4_cascade_ ));
    InMux I__2033 (
            .O(N__16580),
            .I(N__16577));
    LocalMux I__2032 (
            .O(N__16577),
            .I(\VPP_VDDQ.count_2_0_4 ));
    InMux I__2031 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__2030 (
            .O(N__16571),
            .I(\VPP_VDDQ.count_2_0_5 ));
    CascadeMux I__2029 (
            .O(N__16568),
            .I(\VPP_VDDQ.count_2_1_5_cascade_ ));
    CascadeMux I__2028 (
            .O(N__16565),
            .I(\VPP_VDDQ.count_2_1_12_cascade_ ));
    InMux I__2027 (
            .O(N__16562),
            .I(bfn_2_16_0_));
    InMux I__2026 (
            .O(N__16559),
            .I(N__16555));
    InMux I__2025 (
            .O(N__16558),
            .I(N__16552));
    LocalMux I__2024 (
            .O(N__16555),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    LocalMux I__2023 (
            .O(N__16552),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    CEMux I__2022 (
            .O(N__16547),
            .I(N__16544));
    LocalMux I__2021 (
            .O(N__16544),
            .I(N__16541));
    Span4Mux_v I__2020 (
            .O(N__16541),
            .I(N__16538));
    Span4Mux_s1_h I__2019 (
            .O(N__16538),
            .I(N__16535));
    Odrv4 I__2018 (
            .O(N__16535),
            .I(\VPP_VDDQ.N_92_0 ));
    SRMux I__2017 (
            .O(N__16532),
            .I(N__16527));
    SRMux I__2016 (
            .O(N__16531),
            .I(N__16524));
    SRMux I__2015 (
            .O(N__16530),
            .I(N__16521));
    LocalMux I__2014 (
            .O(N__16527),
            .I(N__16518));
    LocalMux I__2013 (
            .O(N__16524),
            .I(N__16513));
    LocalMux I__2012 (
            .O(N__16521),
            .I(N__16513));
    Span4Mux_v I__2011 (
            .O(N__16518),
            .I(N__16508));
    Span4Mux_v I__2010 (
            .O(N__16513),
            .I(N__16508));
    Span4Mux_s1_h I__2009 (
            .O(N__16508),
            .I(N__16505));
    Odrv4 I__2008 (
            .O(N__16505),
            .I(G_30));
    CascadeMux I__2007 (
            .O(N__16502),
            .I(\VPP_VDDQ.count_2_1_8_cascade_ ));
    InMux I__2006 (
            .O(N__16499),
            .I(N__16496));
    LocalMux I__2005 (
            .O(N__16496),
            .I(\VPP_VDDQ.count_2_0_8 ));
    CascadeMux I__2004 (
            .O(N__16493),
            .I(\VPP_VDDQ.count_2_1_9_cascade_ ));
    InMux I__2003 (
            .O(N__16490),
            .I(N__16487));
    LocalMux I__2002 (
            .O(N__16487),
            .I(\VPP_VDDQ.count_2_0_9 ));
    InMux I__2001 (
            .O(N__16484),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__2000 (
            .O(N__16481),
            .I(N__16477));
    InMux I__1999 (
            .O(N__16480),
            .I(N__16474));
    LocalMux I__1998 (
            .O(N__16477),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    LocalMux I__1997 (
            .O(N__16474),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__1996 (
            .O(N__16469),
            .I(bfn_2_15_0_));
    InMux I__1995 (
            .O(N__16466),
            .I(N__16462));
    InMux I__1994 (
            .O(N__16465),
            .I(N__16459));
    LocalMux I__1993 (
            .O(N__16462),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__1992 (
            .O(N__16459),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__1991 (
            .O(N__16454),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    InMux I__1990 (
            .O(N__16451),
            .I(N__16447));
    InMux I__1989 (
            .O(N__16450),
            .I(N__16444));
    LocalMux I__1988 (
            .O(N__16447),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__1987 (
            .O(N__16444),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__1986 (
            .O(N__16439),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    CascadeMux I__1985 (
            .O(N__16436),
            .I(N__16432));
    InMux I__1984 (
            .O(N__16435),
            .I(N__16429));
    InMux I__1983 (
            .O(N__16432),
            .I(N__16426));
    LocalMux I__1982 (
            .O(N__16429),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__1981 (
            .O(N__16426),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__1980 (
            .O(N__16421),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    CascadeMux I__1979 (
            .O(N__16418),
            .I(N__16414));
    InMux I__1978 (
            .O(N__16417),
            .I(N__16411));
    InMux I__1977 (
            .O(N__16414),
            .I(N__16408));
    LocalMux I__1976 (
            .O(N__16411),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    LocalMux I__1975 (
            .O(N__16408),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__1974 (
            .O(N__16403),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    InMux I__1973 (
            .O(N__16400),
            .I(N__16396));
    InMux I__1972 (
            .O(N__16399),
            .I(N__16393));
    LocalMux I__1971 (
            .O(N__16396),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__1970 (
            .O(N__16393),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__1969 (
            .O(N__16388),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__1968 (
            .O(N__16385),
            .I(N__16381));
    InMux I__1967 (
            .O(N__16384),
            .I(N__16378));
    LocalMux I__1966 (
            .O(N__16381),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__1965 (
            .O(N__16378),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__1964 (
            .O(N__16373),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    CascadeMux I__1963 (
            .O(N__16370),
            .I(\POWERLED.un79_clk_100khz_cascade_ ));
    InMux I__1962 (
            .O(N__16367),
            .I(N__16352));
    InMux I__1961 (
            .O(N__16366),
            .I(N__16352));
    InMux I__1960 (
            .O(N__16365),
            .I(N__16352));
    InMux I__1959 (
            .O(N__16364),
            .I(N__16352));
    InMux I__1958 (
            .O(N__16363),
            .I(N__16349));
    InMux I__1957 (
            .O(N__16362),
            .I(N__16344));
    InMux I__1956 (
            .O(N__16361),
            .I(N__16344));
    LocalMux I__1955 (
            .O(N__16352),
            .I(\POWERLED.N_2360_i ));
    LocalMux I__1954 (
            .O(N__16349),
            .I(\POWERLED.N_2360_i ));
    LocalMux I__1953 (
            .O(N__16344),
            .I(\POWERLED.N_2360_i ));
    SRMux I__1952 (
            .O(N__16337),
            .I(N__16334));
    LocalMux I__1951 (
            .O(N__16334),
            .I(N__16331));
    Span4Mux_s1_h I__1950 (
            .O(N__16331),
            .I(N__16328));
    Odrv4 I__1949 (
            .O(N__16328),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    CascadeMux I__1948 (
            .O(N__16325),
            .I(N__16321));
    InMux I__1947 (
            .O(N__16324),
            .I(N__16318));
    InMux I__1946 (
            .O(N__16321),
            .I(N__16315));
    LocalMux I__1945 (
            .O(N__16318),
            .I(N__16310));
    LocalMux I__1944 (
            .O(N__16315),
            .I(N__16310));
    Odrv12 I__1943 (
            .O(N__16310),
            .I(\VPP_VDDQ.N_64_i ));
    InMux I__1942 (
            .O(N__16307),
            .I(N__16303));
    InMux I__1941 (
            .O(N__16306),
            .I(N__16300));
    LocalMux I__1940 (
            .O(N__16303),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__1939 (
            .O(N__16300),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    CascadeMux I__1938 (
            .O(N__16295),
            .I(N__16291));
    InMux I__1937 (
            .O(N__16294),
            .I(N__16288));
    InMux I__1936 (
            .O(N__16291),
            .I(N__16285));
    LocalMux I__1935 (
            .O(N__16288),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__1934 (
            .O(N__16285),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__1933 (
            .O(N__16280),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__1932 (
            .O(N__16277),
            .I(N__16273));
    InMux I__1931 (
            .O(N__16276),
            .I(N__16270));
    LocalMux I__1930 (
            .O(N__16273),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__1929 (
            .O(N__16270),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__1928 (
            .O(N__16265),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__1927 (
            .O(N__16262),
            .I(N__16258));
    InMux I__1926 (
            .O(N__16261),
            .I(N__16255));
    LocalMux I__1925 (
            .O(N__16258),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__1924 (
            .O(N__16255),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__1923 (
            .O(N__16250),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__1922 (
            .O(N__16247),
            .I(N__16243));
    InMux I__1921 (
            .O(N__16246),
            .I(N__16240));
    LocalMux I__1920 (
            .O(N__16243),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__1919 (
            .O(N__16240),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__1918 (
            .O(N__16235),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__1917 (
            .O(N__16232),
            .I(N__16228));
    InMux I__1916 (
            .O(N__16231),
            .I(N__16225));
    LocalMux I__1915 (
            .O(N__16228),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__1914 (
            .O(N__16225),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__1913 (
            .O(N__16220),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__1912 (
            .O(N__16217),
            .I(N__16213));
    InMux I__1911 (
            .O(N__16216),
            .I(N__16210));
    LocalMux I__1910 (
            .O(N__16213),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__1909 (
            .O(N__16210),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__1908 (
            .O(N__16205),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    CascadeMux I__1907 (
            .O(N__16202),
            .I(N__16198));
    InMux I__1906 (
            .O(N__16201),
            .I(N__16195));
    InMux I__1905 (
            .O(N__16198),
            .I(N__16192));
    LocalMux I__1904 (
            .O(N__16195),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__1903 (
            .O(N__16192),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__1902 (
            .O(N__16187),
            .I(N__16184));
    LocalMux I__1901 (
            .O(N__16184),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__1900 (
            .O(N__16181),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    InMux I__1899 (
            .O(N__16178),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__1898 (
            .O(N__16175),
            .I(N__16172));
    InMux I__1897 (
            .O(N__16172),
            .I(N__16163));
    InMux I__1896 (
            .O(N__16171),
            .I(N__16163));
    InMux I__1895 (
            .O(N__16170),
            .I(N__16163));
    LocalMux I__1894 (
            .O(N__16163),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    CascadeMux I__1893 (
            .O(N__16160),
            .I(\POWERLED.count_1_5_cascade_ ));
    InMux I__1892 (
            .O(N__16157),
            .I(N__16150));
    InMux I__1891 (
            .O(N__16156),
            .I(N__16150));
    InMux I__1890 (
            .O(N__16155),
            .I(N__16147));
    LocalMux I__1889 (
            .O(N__16150),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__1888 (
            .O(N__16147),
            .I(\POWERLED.countZ0Z_5 ));
    CascadeMux I__1887 (
            .O(N__16142),
            .I(N__16139));
    InMux I__1886 (
            .O(N__16139),
            .I(N__16133));
    InMux I__1885 (
            .O(N__16138),
            .I(N__16133));
    LocalMux I__1884 (
            .O(N__16133),
            .I(\POWERLED.count_1_5 ));
    CascadeMux I__1883 (
            .O(N__16130),
            .I(\POWERLED.un79_clk_100khzlto6_0_cascade_ ));
    InMux I__1882 (
            .O(N__16127),
            .I(N__16123));
    InMux I__1881 (
            .O(N__16126),
            .I(N__16120));
    LocalMux I__1880 (
            .O(N__16123),
            .I(\POWERLED.un79_clk_100khz ));
    LocalMux I__1879 (
            .O(N__16120),
            .I(\POWERLED.un79_clk_100khz ));
    InMux I__1878 (
            .O(N__16115),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    CascadeMux I__1877 (
            .O(N__16112),
            .I(N__16109));
    InMux I__1876 (
            .O(N__16109),
            .I(N__16106));
    LocalMux I__1875 (
            .O(N__16106),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__1874 (
            .O(N__16103),
            .I(N__16100));
    LocalMux I__1873 (
            .O(N__16100),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__1872 (
            .O(N__16097),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__1871 (
            .O(N__16094),
            .I(N__16091));
    LocalMux I__1870 (
            .O(N__16091),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__1869 (
            .O(N__16088),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__1868 (
            .O(N__16085),
            .I(N__16081));
    InMux I__1867 (
            .O(N__16084),
            .I(N__16073));
    InMux I__1866 (
            .O(N__16081),
            .I(N__16073));
    InMux I__1865 (
            .O(N__16080),
            .I(N__16073));
    LocalMux I__1864 (
            .O(N__16073),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    InMux I__1863 (
            .O(N__16070),
            .I(N__16067));
    LocalMux I__1862 (
            .O(N__16067),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__1861 (
            .O(N__16064),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    CascadeMux I__1860 (
            .O(N__16061),
            .I(N__16058));
    InMux I__1859 (
            .O(N__16058),
            .I(N__16055));
    LocalMux I__1858 (
            .O(N__16055),
            .I(N__16052));
    Odrv4 I__1857 (
            .O(N__16052),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__1856 (
            .O(N__16049),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    InMux I__1855 (
            .O(N__16046),
            .I(N__16043));
    LocalMux I__1854 (
            .O(N__16043),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__1853 (
            .O(N__16040),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    CascadeMux I__1852 (
            .O(N__16037),
            .I(N__16034));
    InMux I__1851 (
            .O(N__16034),
            .I(N__16031));
    LocalMux I__1850 (
            .O(N__16031),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    InMux I__1849 (
            .O(N__16028),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    CascadeMux I__1848 (
            .O(N__16025),
            .I(N__16022));
    InMux I__1847 (
            .O(N__16022),
            .I(N__16019));
    LocalMux I__1846 (
            .O(N__16019),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__1845 (
            .O(N__16016),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    InMux I__1844 (
            .O(N__16013),
            .I(N__16010));
    LocalMux I__1843 (
            .O(N__16010),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__1842 (
            .O(N__16007),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__1841 (
            .O(N__16004),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    CascadeMux I__1840 (
            .O(N__16001),
            .I(N__15998));
    InMux I__1839 (
            .O(N__15998),
            .I(N__15995));
    LocalMux I__1838 (
            .O(N__15995),
            .I(\POWERLED.mult1_un124_sum_axb_4_l_fx ));
    InMux I__1837 (
            .O(N__15992),
            .I(N__15986));
    InMux I__1836 (
            .O(N__15991),
            .I(N__15986));
    LocalMux I__1835 (
            .O(N__15986),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__1834 (
            .O(N__15983),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__1833 (
            .O(N__15980),
            .I(N__15977));
    LocalMux I__1832 (
            .O(N__15977),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    CascadeMux I__1831 (
            .O(N__15974),
            .I(N__15971));
    InMux I__1830 (
            .O(N__15971),
            .I(N__15968));
    LocalMux I__1829 (
            .O(N__15968),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__1828 (
            .O(N__15965),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__1827 (
            .O(N__15962),
            .I(N__15959));
    LocalMux I__1826 (
            .O(N__15959),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__1825 (
            .O(N__15956),
            .I(N__15953));
    LocalMux I__1824 (
            .O(N__15953),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__1823 (
            .O(N__15950),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    CascadeMux I__1822 (
            .O(N__15947),
            .I(N__15944));
    InMux I__1821 (
            .O(N__15944),
            .I(N__15941));
    LocalMux I__1820 (
            .O(N__15941),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    CascadeMux I__1819 (
            .O(N__15938),
            .I(N_626_cascade_));
    CascadeMux I__1818 (
            .O(N__15935),
            .I(\POWERLED.G_30Z0Z_0_cascade_ ));
    InMux I__1817 (
            .O(N__15932),
            .I(N__15926));
    InMux I__1816 (
            .O(N__15931),
            .I(N__15926));
    LocalMux I__1815 (
            .O(N__15926),
            .I(N__15923));
    Span4Mux_v I__1814 (
            .O(N__15923),
            .I(N__15920));
    Odrv4 I__1813 (
            .O(N__15920),
            .I(VPP_VDDQ_un6_count));
    CascadeMux I__1812 (
            .O(N__15917),
            .I(G_30_cascade_));
    InMux I__1811 (
            .O(N__15914),
            .I(N__15911));
    LocalMux I__1810 (
            .O(N__15911),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__1809 (
            .O(N__15908),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    CascadeMux I__1808 (
            .O(N__15905),
            .I(N__15902));
    InMux I__1807 (
            .O(N__15902),
            .I(N__15899));
    LocalMux I__1806 (
            .O(N__15899),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__1805 (
            .O(N__15896),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__1804 (
            .O(N__15893),
            .I(N__15890));
    LocalMux I__1803 (
            .O(N__15890),
            .I(N__15887));
    Odrv4 I__1802 (
            .O(N__15887),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__1801 (
            .O(N__15884),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__1800 (
            .O(N__15881),
            .I(N__15878));
    LocalMux I__1799 (
            .O(N__15878),
            .I(N__15875));
    Odrv12 I__1798 (
            .O(N__15875),
            .I(\PCH_PWRGD.curr_state_0_0 ));
    InMux I__1797 (
            .O(N__15872),
            .I(N__15869));
    LocalMux I__1796 (
            .O(N__15869),
            .I(\PCH_PWRGD.N_2244_i ));
    InMux I__1795 (
            .O(N__15866),
            .I(N__15860));
    InMux I__1794 (
            .O(N__15865),
            .I(N__15860));
    LocalMux I__1793 (
            .O(N__15860),
            .I(N__15857));
    Span4Mux_v I__1792 (
            .O(N__15857),
            .I(N__15854));
    Odrv4 I__1791 (
            .O(N__15854),
            .I(vr_ready_vccin));
    CascadeMux I__1790 (
            .O(N__15851),
            .I(\PCH_PWRGD.N_2244_i_cascade_ ));
    CascadeMux I__1789 (
            .O(N__15848),
            .I(\PCH_PWRGD.N_655_cascade_ ));
    InMux I__1788 (
            .O(N__15845),
            .I(N__15842));
    LocalMux I__1787 (
            .O(N__15842),
            .I(\PCH_PWRGD.m6_i_i_a2 ));
    InMux I__1786 (
            .O(N__15839),
            .I(N__15835));
    CascadeMux I__1785 (
            .O(N__15838),
            .I(N__15832));
    LocalMux I__1784 (
            .O(N__15835),
            .I(N__15827));
    InMux I__1783 (
            .O(N__15832),
            .I(N__15824));
    InMux I__1782 (
            .O(N__15831),
            .I(N__15819));
    InMux I__1781 (
            .O(N__15830),
            .I(N__15819));
    Odrv12 I__1780 (
            .O(N__15827),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__1779 (
            .O(N__15824),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__1778 (
            .O(N__15819),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    InMux I__1777 (
            .O(N__15812),
            .I(N__15806));
    InMux I__1776 (
            .O(N__15811),
            .I(N__15806));
    LocalMux I__1775 (
            .O(N__15806),
            .I(N__15789));
    InMux I__1774 (
            .O(N__15805),
            .I(N__15784));
    InMux I__1773 (
            .O(N__15804),
            .I(N__15784));
    InMux I__1772 (
            .O(N__15803),
            .I(N__15781));
    InMux I__1771 (
            .O(N__15802),
            .I(N__15777));
    InMux I__1770 (
            .O(N__15801),
            .I(N__15770));
    InMux I__1769 (
            .O(N__15800),
            .I(N__15770));
    InMux I__1768 (
            .O(N__15799),
            .I(N__15770));
    InMux I__1767 (
            .O(N__15798),
            .I(N__15763));
    InMux I__1766 (
            .O(N__15797),
            .I(N__15763));
    InMux I__1765 (
            .O(N__15796),
            .I(N__15763));
    InMux I__1764 (
            .O(N__15795),
            .I(N__15754));
    InMux I__1763 (
            .O(N__15794),
            .I(N__15754));
    InMux I__1762 (
            .O(N__15793),
            .I(N__15754));
    InMux I__1761 (
            .O(N__15792),
            .I(N__15754));
    Span4Mux_s1_h I__1760 (
            .O(N__15789),
            .I(N__15747));
    LocalMux I__1759 (
            .O(N__15784),
            .I(N__15747));
    LocalMux I__1758 (
            .O(N__15781),
            .I(N__15747));
    InMux I__1757 (
            .O(N__15780),
            .I(N__15744));
    LocalMux I__1756 (
            .O(N__15777),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1755 (
            .O(N__15770),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1754 (
            .O(N__15763),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1753 (
            .O(N__15754),
            .I(\PCH_PWRGD.N_386 ));
    Odrv4 I__1752 (
            .O(N__15747),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1751 (
            .O(N__15744),
            .I(\PCH_PWRGD.N_386 ));
    InMux I__1750 (
            .O(N__15731),
            .I(N__15724));
    InMux I__1749 (
            .O(N__15730),
            .I(N__15721));
    InMux I__1748 (
            .O(N__15729),
            .I(N__15718));
    InMux I__1747 (
            .O(N__15728),
            .I(N__15715));
    InMux I__1746 (
            .O(N__15727),
            .I(N__15712));
    LocalMux I__1745 (
            .O(N__15724),
            .I(N__15707));
    LocalMux I__1744 (
            .O(N__15721),
            .I(N__15707));
    LocalMux I__1743 (
            .O(N__15718),
            .I(N__15702));
    LocalMux I__1742 (
            .O(N__15715),
            .I(N__15702));
    LocalMux I__1741 (
            .O(N__15712),
            .I(N__15699));
    Span4Mux_v I__1740 (
            .O(N__15707),
            .I(N__15696));
    Odrv12 I__1739 (
            .O(N__15702),
            .I(\PCH_PWRGD.N_2226_i ));
    Odrv4 I__1738 (
            .O(N__15699),
            .I(\PCH_PWRGD.N_2226_i ));
    Odrv4 I__1737 (
            .O(N__15696),
            .I(\PCH_PWRGD.N_2226_i ));
    CascadeMux I__1736 (
            .O(N__15689),
            .I(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ));
    InMux I__1735 (
            .O(N__15686),
            .I(N__15681));
    InMux I__1734 (
            .O(N__15685),
            .I(N__15678));
    InMux I__1733 (
            .O(N__15684),
            .I(N__15675));
    LocalMux I__1732 (
            .O(N__15681),
            .I(\PCH_PWRGD.N_655 ));
    LocalMux I__1731 (
            .O(N__15678),
            .I(\PCH_PWRGD.N_655 ));
    LocalMux I__1730 (
            .O(N__15675),
            .I(\PCH_PWRGD.N_655 ));
    InMux I__1729 (
            .O(N__15668),
            .I(N__15665));
    LocalMux I__1728 (
            .O(N__15665),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    InMux I__1727 (
            .O(N__15662),
            .I(N__15659));
    LocalMux I__1726 (
            .O(N__15659),
            .I(\PCH_PWRGD.count_rst_14 ));
    InMux I__1725 (
            .O(N__15656),
            .I(N__15653));
    LocalMux I__1724 (
            .O(N__15653),
            .I(\PCH_PWRGD.count_0_0 ));
    CascadeMux I__1723 (
            .O(N__15650),
            .I(\PCH_PWRGD.count_0_sqmuxa_cascade_ ));
    InMux I__1722 (
            .O(N__15647),
            .I(N__15644));
    LocalMux I__1721 (
            .O(N__15644),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    CascadeMux I__1720 (
            .O(N__15641),
            .I(\PCH_PWRGD.countZ0Z_6_cascade_ ));
    InMux I__1719 (
            .O(N__15638),
            .I(N__15635));
    LocalMux I__1718 (
            .O(N__15635),
            .I(\PCH_PWRGD.count_1_i_a2_0_0 ));
    CascadeMux I__1717 (
            .O(N__15632),
            .I(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ));
    InMux I__1716 (
            .O(N__15629),
            .I(N__15626));
    LocalMux I__1715 (
            .O(N__15626),
            .I(N__15622));
    InMux I__1714 (
            .O(N__15625),
            .I(N__15619));
    Odrv12 I__1713 (
            .O(N__15622),
            .I(\PCH_PWRGD.count_rst_13 ));
    LocalMux I__1712 (
            .O(N__15619),
            .I(\PCH_PWRGD.count_rst_13 ));
    InMux I__1711 (
            .O(N__15614),
            .I(N__15608));
    InMux I__1710 (
            .O(N__15613),
            .I(N__15608));
    LocalMux I__1709 (
            .O(N__15608),
            .I(\PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ));
    InMux I__1708 (
            .O(N__15605),
            .I(N__15602));
    LocalMux I__1707 (
            .O(N__15602),
            .I(\PCH_PWRGD.count_0_6 ));
    InMux I__1706 (
            .O(N__15599),
            .I(N__15596));
    LocalMux I__1705 (
            .O(N__15596),
            .I(\PCH_PWRGD.un2_count_1_axb_10 ));
    InMux I__1704 (
            .O(N__15593),
            .I(N__15584));
    InMux I__1703 (
            .O(N__15592),
            .I(N__15584));
    InMux I__1702 (
            .O(N__15591),
            .I(N__15584));
    LocalMux I__1701 (
            .O(N__15584),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__1700 (
            .O(N__15581),
            .I(N__15575));
    InMux I__1699 (
            .O(N__15580),
            .I(N__15575));
    LocalMux I__1698 (
            .O(N__15575),
            .I(\PCH_PWRGD.count_0_10 ));
    InMux I__1697 (
            .O(N__15572),
            .I(N__15566));
    InMux I__1696 (
            .O(N__15571),
            .I(N__15566));
    LocalMux I__1695 (
            .O(N__15566),
            .I(N__15563));
    Odrv4 I__1694 (
            .O(N__15563),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    CascadeMux I__1693 (
            .O(N__15560),
            .I(\PCH_PWRGD.countZ0Z_3_cascade_ ));
    InMux I__1692 (
            .O(N__15557),
            .I(N__15554));
    LocalMux I__1691 (
            .O(N__15554),
            .I(\PCH_PWRGD.count_0_3 ));
    InMux I__1690 (
            .O(N__15551),
            .I(N__15548));
    LocalMux I__1689 (
            .O(N__15548),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    CascadeMux I__1688 (
            .O(N__15545),
            .I(\PCH_PWRGD.countZ0Z_14_cascade_ ));
    InMux I__1687 (
            .O(N__15542),
            .I(N__15538));
    InMux I__1686 (
            .O(N__15541),
            .I(N__15535));
    LocalMux I__1685 (
            .O(N__15538),
            .I(N__15532));
    LocalMux I__1684 (
            .O(N__15535),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    Odrv4 I__1683 (
            .O(N__15532),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    CascadeMux I__1682 (
            .O(N__15527),
            .I(\PCH_PWRGD.count_1_i_a2_1_0_cascade_ ));
    InMux I__1681 (
            .O(N__15524),
            .I(N__15521));
    LocalMux I__1680 (
            .O(N__15521),
            .I(N__15518));
    Odrv4 I__1679 (
            .O(N__15518),
            .I(\PCH_PWRGD.count_1_i_a2_2_0 ));
    CascadeMux I__1678 (
            .O(N__15515),
            .I(N__15512));
    InMux I__1677 (
            .O(N__15512),
            .I(N__15506));
    InMux I__1676 (
            .O(N__15511),
            .I(N__15506));
    LocalMux I__1675 (
            .O(N__15506),
            .I(\PCH_PWRGD.count_1_i_a2_11_0 ));
    CascadeMux I__1674 (
            .O(N__15503),
            .I(\PCH_PWRGD.count_1_i_a2_11_0_cascade_ ));
    InMux I__1673 (
            .O(N__15500),
            .I(N__15497));
    LocalMux I__1672 (
            .O(N__15497),
            .I(N__15492));
    InMux I__1671 (
            .O(N__15496),
            .I(N__15487));
    InMux I__1670 (
            .O(N__15495),
            .I(N__15487));
    Odrv4 I__1669 (
            .O(N__15492),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    LocalMux I__1668 (
            .O(N__15487),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    InMux I__1667 (
            .O(N__15482),
            .I(N__15476));
    InMux I__1666 (
            .O(N__15481),
            .I(N__15476));
    LocalMux I__1665 (
            .O(N__15476),
            .I(\PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ));
    CascadeMux I__1664 (
            .O(N__15473),
            .I(N__15470));
    InMux I__1663 (
            .O(N__15470),
            .I(N__15467));
    LocalMux I__1662 (
            .O(N__15467),
            .I(\PCH_PWRGD.count_0_14 ));
    InMux I__1661 (
            .O(N__15464),
            .I(N__15455));
    InMux I__1660 (
            .O(N__15463),
            .I(N__15455));
    InMux I__1659 (
            .O(N__15462),
            .I(N__15455));
    LocalMux I__1658 (
            .O(N__15455),
            .I(\PCH_PWRGD.count_rst_12 ));
    InMux I__1657 (
            .O(N__15452),
            .I(N__15446));
    InMux I__1656 (
            .O(N__15451),
            .I(N__15446));
    LocalMux I__1655 (
            .O(N__15446),
            .I(\PCH_PWRGD.count_0_2 ));
    InMux I__1654 (
            .O(N__15443),
            .I(N__15440));
    LocalMux I__1653 (
            .O(N__15440),
            .I(\PCH_PWRGD.un2_count_1_axb_2 ));
    CascadeMux I__1652 (
            .O(N__15437),
            .I(\PCH_PWRGD.countZ0Z_11_cascade_ ));
    InMux I__1651 (
            .O(N__15434),
            .I(N__15431));
    LocalMux I__1650 (
            .O(N__15431),
            .I(\PCH_PWRGD.count_1_i_a2_4_0 ));
    InMux I__1649 (
            .O(N__15428),
            .I(N__15425));
    LocalMux I__1648 (
            .O(N__15425),
            .I(\PCH_PWRGD.count_1_i_a2_5_0 ));
    CascadeMux I__1647 (
            .O(N__15422),
            .I(\PCH_PWRGD.count_1_i_a2_3_0_cascade_ ));
    InMux I__1646 (
            .O(N__15419),
            .I(N__15416));
    LocalMux I__1645 (
            .O(N__15416),
            .I(\PCH_PWRGD.count_1_i_a2_6_0 ));
    CascadeMux I__1644 (
            .O(N__15413),
            .I(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__1643 (
            .O(N__15410),
            .I(\PCH_PWRGD.N_2226_i_cascade_ ));
    InMux I__1642 (
            .O(N__15407),
            .I(N__15404));
    LocalMux I__1641 (
            .O(N__15404),
            .I(\PCH_PWRGD.curr_state_7_0 ));
    CascadeMux I__1640 (
            .O(N__15401),
            .I(\PCH_PWRGD.N_386_cascade_ ));
    CascadeMux I__1639 (
            .O(N__15398),
            .I(\PCH_PWRGD.count_rst_11_cascade_ ));
    InMux I__1638 (
            .O(N__15395),
            .I(N__15390));
    InMux I__1637 (
            .O(N__15394),
            .I(N__15387));
    InMux I__1636 (
            .O(N__15393),
            .I(N__15384));
    LocalMux I__1635 (
            .O(N__15390),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__1634 (
            .O(N__15387),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__1633 (
            .O(N__15384),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    InMux I__1632 (
            .O(N__15377),
            .I(N__15373));
    InMux I__1631 (
            .O(N__15376),
            .I(N__15370));
    LocalMux I__1630 (
            .O(N__15373),
            .I(\HDA_STRAP.countZ0Z_15 ));
    LocalMux I__1629 (
            .O(N__15370),
            .I(\HDA_STRAP.countZ0Z_15 ));
    InMux I__1628 (
            .O(N__15365),
            .I(\HDA_STRAP.un1_count_1_cry_14 ));
    InMux I__1627 (
            .O(N__15362),
            .I(N__15357));
    InMux I__1626 (
            .O(N__15361),
            .I(N__15352));
    InMux I__1625 (
            .O(N__15360),
            .I(N__15352));
    LocalMux I__1624 (
            .O(N__15357),
            .I(\HDA_STRAP.countZ0Z_16 ));
    LocalMux I__1623 (
            .O(N__15352),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__1622 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__1621 (
            .O(N__15344),
            .I(\HDA_STRAP.un1_count_1_cry_15_THRU_CO ));
    InMux I__1620 (
            .O(N__15341),
            .I(bfn_2_3_0_));
    CascadeMux I__1619 (
            .O(N__15338),
            .I(N__15330));
    CascadeMux I__1618 (
            .O(N__15337),
            .I(N__15326));
    InMux I__1617 (
            .O(N__15336),
            .I(N__15321));
    InMux I__1616 (
            .O(N__15335),
            .I(N__15321));
    CascadeMux I__1615 (
            .O(N__15334),
            .I(N__15316));
    CascadeMux I__1614 (
            .O(N__15333),
            .I(N__15313));
    InMux I__1613 (
            .O(N__15330),
            .I(N__15309));
    InMux I__1612 (
            .O(N__15329),
            .I(N__15306));
    InMux I__1611 (
            .O(N__15326),
            .I(N__15303));
    LocalMux I__1610 (
            .O(N__15321),
            .I(N__15300));
    InMux I__1609 (
            .O(N__15320),
            .I(N__15289));
    InMux I__1608 (
            .O(N__15319),
            .I(N__15289));
    InMux I__1607 (
            .O(N__15316),
            .I(N__15289));
    InMux I__1606 (
            .O(N__15313),
            .I(N__15289));
    InMux I__1605 (
            .O(N__15312),
            .I(N__15289));
    LocalMux I__1604 (
            .O(N__15309),
            .I(N__15284));
    LocalMux I__1603 (
            .O(N__15306),
            .I(N__15284));
    LocalMux I__1602 (
            .O(N__15303),
            .I(N__15281));
    Odrv4 I__1601 (
            .O(N__15300),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    LocalMux I__1600 (
            .O(N__15289),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    Odrv4 I__1599 (
            .O(N__15284),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    Odrv4 I__1598 (
            .O(N__15281),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    CascadeMux I__1597 (
            .O(N__15272),
            .I(N__15267));
    CascadeMux I__1596 (
            .O(N__15271),
            .I(N__15263));
    InMux I__1595 (
            .O(N__15270),
            .I(N__15253));
    InMux I__1594 (
            .O(N__15267),
            .I(N__15253));
    InMux I__1593 (
            .O(N__15266),
            .I(N__15250));
    InMux I__1592 (
            .O(N__15263),
            .I(N__15247));
    InMux I__1591 (
            .O(N__15262),
            .I(N__15236));
    InMux I__1590 (
            .O(N__15261),
            .I(N__15236));
    InMux I__1589 (
            .O(N__15260),
            .I(N__15236));
    InMux I__1588 (
            .O(N__15259),
            .I(N__15236));
    InMux I__1587 (
            .O(N__15258),
            .I(N__15236));
    LocalMux I__1586 (
            .O(N__15253),
            .I(N__15233));
    LocalMux I__1585 (
            .O(N__15250),
            .I(\HDA_STRAP.un4_count ));
    LocalMux I__1584 (
            .O(N__15247),
            .I(\HDA_STRAP.un4_count ));
    LocalMux I__1583 (
            .O(N__15236),
            .I(\HDA_STRAP.un4_count ));
    Odrv4 I__1582 (
            .O(N__15233),
            .I(\HDA_STRAP.un4_count ));
    InMux I__1581 (
            .O(N__15224),
            .I(\HDA_STRAP.un1_count_1_cry_16 ));
    InMux I__1580 (
            .O(N__15221),
            .I(N__15217));
    InMux I__1579 (
            .O(N__15220),
            .I(N__15214));
    LocalMux I__1578 (
            .O(N__15217),
            .I(\HDA_STRAP.countZ0Z_17 ));
    LocalMux I__1577 (
            .O(N__15214),
            .I(\HDA_STRAP.countZ0Z_17 ));
    CascadeMux I__1576 (
            .O(N__15209),
            .I(N__15205));
    InMux I__1575 (
            .O(N__15208),
            .I(N__15202));
    InMux I__1574 (
            .O(N__15205),
            .I(N__15199));
    LocalMux I__1573 (
            .O(N__15202),
            .I(N__15194));
    LocalMux I__1572 (
            .O(N__15199),
            .I(N__15194));
    Span4Mux_s3_v I__1571 (
            .O(N__15194),
            .I(N__15191));
    Odrv4 I__1570 (
            .O(N__15191),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    InMux I__1569 (
            .O(N__15188),
            .I(N__15183));
    InMux I__1568 (
            .O(N__15187),
            .I(N__15180));
    InMux I__1567 (
            .O(N__15186),
            .I(N__15177));
    LocalMux I__1566 (
            .O(N__15183),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1565 (
            .O(N__15180),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1564 (
            .O(N__15177),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    CascadeMux I__1563 (
            .O(N__15170),
            .I(\PCH_PWRGD.count_rst_7_cascade_ ));
    InMux I__1562 (
            .O(N__15167),
            .I(N__15161));
    InMux I__1561 (
            .O(N__15166),
            .I(N__15161));
    LocalMux I__1560 (
            .O(N__15161),
            .I(N__15158));
    Span4Mux_h I__1559 (
            .O(N__15158),
            .I(N__15155));
    Odrv4 I__1558 (
            .O(N__15155),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    InMux I__1557 (
            .O(N__15152),
            .I(N__15149));
    LocalMux I__1556 (
            .O(N__15149),
            .I(\PCH_PWRGD.count_rst_7 ));
    InMux I__1555 (
            .O(N__15146),
            .I(N__15140));
    InMux I__1554 (
            .O(N__15145),
            .I(N__15140));
    LocalMux I__1553 (
            .O(N__15140),
            .I(\PCH_PWRGD.count_0_7 ));
    InMux I__1552 (
            .O(N__15137),
            .I(N__15134));
    LocalMux I__1551 (
            .O(N__15134),
            .I(N__15129));
    InMux I__1550 (
            .O(N__15133),
            .I(N__15124));
    InMux I__1549 (
            .O(N__15132),
            .I(N__15124));
    Odrv4 I__1548 (
            .O(N__15129),
            .I(\PCH_PWRGD.un2_count_1_axb_7 ));
    LocalMux I__1547 (
            .O(N__15124),
            .I(\PCH_PWRGD.un2_count_1_axb_7 ));
    InMux I__1546 (
            .O(N__15119),
            .I(N__15116));
    LocalMux I__1545 (
            .O(N__15116),
            .I(\PCH_PWRGD.count_rst_3 ));
    InMux I__1544 (
            .O(N__15113),
            .I(N__15110));
    LocalMux I__1543 (
            .O(N__15110),
            .I(\PCH_PWRGD.count_0_11 ));
    InMux I__1542 (
            .O(N__15107),
            .I(N__15104));
    LocalMux I__1541 (
            .O(N__15104),
            .I(N__15100));
    CascadeMux I__1540 (
            .O(N__15103),
            .I(N__15097));
    Span12Mux_v I__1539 (
            .O(N__15100),
            .I(N__15093));
    InMux I__1538 (
            .O(N__15097),
            .I(N__15090));
    InMux I__1537 (
            .O(N__15096),
            .I(N__15087));
    Odrv12 I__1536 (
            .O(N__15093),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    LocalMux I__1535 (
            .O(N__15090),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    LocalMux I__1534 (
            .O(N__15087),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    CascadeMux I__1533 (
            .O(N__15080),
            .I(N__15077));
    InMux I__1532 (
            .O(N__15077),
            .I(N__15073));
    InMux I__1531 (
            .O(N__15076),
            .I(N__15070));
    LocalMux I__1530 (
            .O(N__15073),
            .I(\HDA_STRAP.countZ0Z_7 ));
    LocalMux I__1529 (
            .O(N__15070),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__1528 (
            .O(N__15065),
            .I(\HDA_STRAP.un1_count_1_cry_6 ));
    InMux I__1527 (
            .O(N__15062),
            .I(N__15057));
    InMux I__1526 (
            .O(N__15061),
            .I(N__15052));
    InMux I__1525 (
            .O(N__15060),
            .I(N__15052));
    LocalMux I__1524 (
            .O(N__15057),
            .I(\HDA_STRAP.countZ0Z_8 ));
    LocalMux I__1523 (
            .O(N__15052),
            .I(\HDA_STRAP.countZ0Z_8 ));
    CascadeMux I__1522 (
            .O(N__15047),
            .I(N__15044));
    InMux I__1521 (
            .O(N__15044),
            .I(N__15041));
    LocalMux I__1520 (
            .O(N__15041),
            .I(\HDA_STRAP.un1_count_1_cry_7_THRU_CO ));
    InMux I__1519 (
            .O(N__15038),
            .I(bfn_2_2_0_));
    InMux I__1518 (
            .O(N__15035),
            .I(N__15031));
    InMux I__1517 (
            .O(N__15034),
            .I(N__15028));
    LocalMux I__1516 (
            .O(N__15031),
            .I(\HDA_STRAP.countZ0Z_9 ));
    LocalMux I__1515 (
            .O(N__15028),
            .I(\HDA_STRAP.countZ0Z_9 ));
    InMux I__1514 (
            .O(N__15023),
            .I(\HDA_STRAP.un1_count_1_cry_8 ));
    InMux I__1513 (
            .O(N__15020),
            .I(N__15015));
    InMux I__1512 (
            .O(N__15019),
            .I(N__15012));
    InMux I__1511 (
            .O(N__15018),
            .I(N__15009));
    LocalMux I__1510 (
            .O(N__15015),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__1509 (
            .O(N__15012),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__1508 (
            .O(N__15009),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__1507 (
            .O(N__15002),
            .I(N__14999));
    LocalMux I__1506 (
            .O(N__14999),
            .I(\HDA_STRAP.un1_count_1_cry_9_THRU_CO ));
    InMux I__1505 (
            .O(N__14996),
            .I(\HDA_STRAP.un1_count_1_cry_9 ));
    InMux I__1504 (
            .O(N__14993),
            .I(N__14988));
    InMux I__1503 (
            .O(N__14992),
            .I(N__14985));
    InMux I__1502 (
            .O(N__14991),
            .I(N__14982));
    LocalMux I__1501 (
            .O(N__14988),
            .I(\HDA_STRAP.countZ0Z_11 ));
    LocalMux I__1500 (
            .O(N__14985),
            .I(\HDA_STRAP.countZ0Z_11 ));
    LocalMux I__1499 (
            .O(N__14982),
            .I(\HDA_STRAP.countZ0Z_11 ));
    CascadeMux I__1498 (
            .O(N__14975),
            .I(N__14972));
    InMux I__1497 (
            .O(N__14972),
            .I(N__14969));
    LocalMux I__1496 (
            .O(N__14969),
            .I(\HDA_STRAP.un1_count_1_cry_10_THRU_CO ));
    InMux I__1495 (
            .O(N__14966),
            .I(\HDA_STRAP.un1_count_1_cry_10 ));
    InMux I__1494 (
            .O(N__14963),
            .I(N__14959));
    InMux I__1493 (
            .O(N__14962),
            .I(N__14956));
    LocalMux I__1492 (
            .O(N__14959),
            .I(\HDA_STRAP.countZ0Z_12 ));
    LocalMux I__1491 (
            .O(N__14956),
            .I(\HDA_STRAP.countZ0Z_12 ));
    InMux I__1490 (
            .O(N__14951),
            .I(\HDA_STRAP.un1_count_1_cry_11 ));
    InMux I__1489 (
            .O(N__14948),
            .I(N__14944));
    InMux I__1488 (
            .O(N__14947),
            .I(N__14941));
    LocalMux I__1487 (
            .O(N__14944),
            .I(\HDA_STRAP.countZ0Z_13 ));
    LocalMux I__1486 (
            .O(N__14941),
            .I(\HDA_STRAP.countZ0Z_13 ));
    InMux I__1485 (
            .O(N__14936),
            .I(\HDA_STRAP.un1_count_1_cry_12 ));
    InMux I__1484 (
            .O(N__14933),
            .I(N__14929));
    InMux I__1483 (
            .O(N__14932),
            .I(N__14926));
    LocalMux I__1482 (
            .O(N__14929),
            .I(\HDA_STRAP.countZ0Z_14 ));
    LocalMux I__1481 (
            .O(N__14926),
            .I(\HDA_STRAP.countZ0Z_14 ));
    InMux I__1480 (
            .O(N__14921),
            .I(\HDA_STRAP.un1_count_1_cry_13 ));
    InMux I__1479 (
            .O(N__14918),
            .I(N__14915));
    LocalMux I__1478 (
            .O(N__14915),
            .I(N__14912));
    Span4Mux_s3_v I__1477 (
            .O(N__14912),
            .I(N__14909));
    Odrv4 I__1476 (
            .O(N__14909),
            .I(vpp_ok));
    IoInMux I__1475 (
            .O(N__14906),
            .I(N__14903));
    LocalMux I__1474 (
            .O(N__14903),
            .I(vddq_en));
    CascadeMux I__1473 (
            .O(N__14900),
            .I(N__14897));
    InMux I__1472 (
            .O(N__14897),
            .I(N__14892));
    InMux I__1471 (
            .O(N__14896),
            .I(N__14889));
    InMux I__1470 (
            .O(N__14895),
            .I(N__14886));
    LocalMux I__1469 (
            .O(N__14892),
            .I(N__14883));
    LocalMux I__1468 (
            .O(N__14889),
            .I(N__14878));
    LocalMux I__1467 (
            .O(N__14886),
            .I(N__14878));
    Odrv4 I__1466 (
            .O(N__14883),
            .I(\HDA_STRAP.countZ0Z_0 ));
    Odrv4 I__1465 (
            .O(N__14878),
            .I(\HDA_STRAP.countZ0Z_0 ));
    InMux I__1464 (
            .O(N__14873),
            .I(N__14870));
    LocalMux I__1463 (
            .O(N__14870),
            .I(N__14866));
    InMux I__1462 (
            .O(N__14869),
            .I(N__14863));
    Odrv4 I__1461 (
            .O(N__14866),
            .I(\HDA_STRAP.countZ0Z_1 ));
    LocalMux I__1460 (
            .O(N__14863),
            .I(\HDA_STRAP.countZ0Z_1 ));
    InMux I__1459 (
            .O(N__14858),
            .I(\HDA_STRAP.un1_count_1_cry_0 ));
    InMux I__1458 (
            .O(N__14855),
            .I(N__14851));
    InMux I__1457 (
            .O(N__14854),
            .I(N__14848));
    LocalMux I__1456 (
            .O(N__14851),
            .I(N__14845));
    LocalMux I__1455 (
            .O(N__14848),
            .I(\HDA_STRAP.countZ0Z_2 ));
    Odrv4 I__1454 (
            .O(N__14845),
            .I(\HDA_STRAP.countZ0Z_2 ));
    InMux I__1453 (
            .O(N__14840),
            .I(\HDA_STRAP.un1_count_1_cry_1 ));
    InMux I__1452 (
            .O(N__14837),
            .I(N__14833));
    InMux I__1451 (
            .O(N__14836),
            .I(N__14830));
    LocalMux I__1450 (
            .O(N__14833),
            .I(N__14827));
    LocalMux I__1449 (
            .O(N__14830),
            .I(\HDA_STRAP.countZ0Z_3 ));
    Odrv4 I__1448 (
            .O(N__14827),
            .I(\HDA_STRAP.countZ0Z_3 ));
    InMux I__1447 (
            .O(N__14822),
            .I(\HDA_STRAP.un1_count_1_cry_2 ));
    CascadeMux I__1446 (
            .O(N__14819),
            .I(N__14816));
    InMux I__1445 (
            .O(N__14816),
            .I(N__14813));
    LocalMux I__1444 (
            .O(N__14813),
            .I(N__14809));
    InMux I__1443 (
            .O(N__14812),
            .I(N__14806));
    Odrv4 I__1442 (
            .O(N__14809),
            .I(\HDA_STRAP.countZ0Z_4 ));
    LocalMux I__1441 (
            .O(N__14806),
            .I(\HDA_STRAP.countZ0Z_4 ));
    InMux I__1440 (
            .O(N__14801),
            .I(\HDA_STRAP.un1_count_1_cry_3 ));
    InMux I__1439 (
            .O(N__14798),
            .I(N__14794));
    InMux I__1438 (
            .O(N__14797),
            .I(N__14791));
    LocalMux I__1437 (
            .O(N__14794),
            .I(N__14788));
    LocalMux I__1436 (
            .O(N__14791),
            .I(\HDA_STRAP.countZ0Z_5 ));
    Odrv4 I__1435 (
            .O(N__14788),
            .I(\HDA_STRAP.countZ0Z_5 ));
    InMux I__1434 (
            .O(N__14783),
            .I(\HDA_STRAP.un1_count_1_cry_4 ));
    CascadeMux I__1433 (
            .O(N__14780),
            .I(N__14776));
    InMux I__1432 (
            .O(N__14779),
            .I(N__14770));
    InMux I__1431 (
            .O(N__14776),
            .I(N__14770));
    InMux I__1430 (
            .O(N__14775),
            .I(N__14767));
    LocalMux I__1429 (
            .O(N__14770),
            .I(\HDA_STRAP.countZ0Z_6 ));
    LocalMux I__1428 (
            .O(N__14767),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__1427 (
            .O(N__14762),
            .I(N__14759));
    LocalMux I__1426 (
            .O(N__14759),
            .I(N__14756));
    Odrv4 I__1425 (
            .O(N__14756),
            .I(\HDA_STRAP.un1_count_1_cry_5_THRU_CO ));
    InMux I__1424 (
            .O(N__14753),
            .I(\HDA_STRAP.un1_count_1_cry_5 ));
    InMux I__1423 (
            .O(N__14750),
            .I(N__14747));
    LocalMux I__1422 (
            .O(N__14747),
            .I(\POWERLED.N_11 ));
    CascadeMux I__1421 (
            .O(N__14744),
            .I(N__14741));
    InMux I__1420 (
            .O(N__14741),
            .I(N__14738));
    LocalMux I__1419 (
            .O(N__14738),
            .I(\POWERLED.g0_2_1 ));
    InMux I__1418 (
            .O(N__14735),
            .I(N__14729));
    InMux I__1417 (
            .O(N__14734),
            .I(N__14729));
    LocalMux I__1416 (
            .O(N__14729),
            .I(\POWERLED.pwm_outZ0 ));
    CascadeMux I__1415 (
            .O(N__14726),
            .I(\POWERLED.N_2360_i_cascade_ ));
    CascadeMux I__1414 (
            .O(N__14723),
            .I(\VPP_VDDQ.un6_count_11_cascade_ ));
    InMux I__1413 (
            .O(N__14720),
            .I(N__14717));
    LocalMux I__1412 (
            .O(N__14717),
            .I(\VPP_VDDQ.un6_count_9 ));
    InMux I__1411 (
            .O(N__14714),
            .I(N__14711));
    LocalMux I__1410 (
            .O(N__14711),
            .I(\VPP_VDDQ.un6_count_10 ));
    InMux I__1409 (
            .O(N__14708),
            .I(N__14705));
    LocalMux I__1408 (
            .O(N__14705),
            .I(\VPP_VDDQ.un6_count_8 ));
    CascadeMux I__1407 (
            .O(N__14702),
            .I(N__14698));
    InMux I__1406 (
            .O(N__14701),
            .I(N__14690));
    InMux I__1405 (
            .O(N__14698),
            .I(N__14690));
    InMux I__1404 (
            .O(N__14697),
            .I(N__14690));
    LocalMux I__1403 (
            .O(N__14690),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    CascadeMux I__1402 (
            .O(N__14687),
            .I(N__14684));
    InMux I__1401 (
            .O(N__14684),
            .I(N__14681));
    LocalMux I__1400 (
            .O(N__14681),
            .I(N__14678));
    Odrv4 I__1399 (
            .O(N__14678),
            .I(\POWERLED.mult1_un96_sum_i ));
    CascadeMux I__1398 (
            .O(N__14675),
            .I(N__14672));
    InMux I__1397 (
            .O(N__14672),
            .I(N__14669));
    LocalMux I__1396 (
            .O(N__14669),
            .I(N__14666));
    Odrv4 I__1395 (
            .O(N__14666),
            .I(\POWERLED.mult1_un103_sum_i ));
    CascadeMux I__1394 (
            .O(N__14663),
            .I(N__14659));
    InMux I__1393 (
            .O(N__14662),
            .I(N__14651));
    InMux I__1392 (
            .O(N__14659),
            .I(N__14651));
    InMux I__1391 (
            .O(N__14658),
            .I(N__14651));
    LocalMux I__1390 (
            .O(N__14651),
            .I(N__14648));
    Odrv4 I__1389 (
            .O(N__14648),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    CascadeMux I__1388 (
            .O(N__14645),
            .I(\POWERLED.g1_i_a4_0_1_cascade_ ));
    InMux I__1387 (
            .O(N__14642),
            .I(N__14639));
    LocalMux I__1386 (
            .O(N__14639),
            .I(\POWERLED.N_12 ));
    CascadeMux I__1385 (
            .O(N__14636),
            .I(\POWERLED.N_5_cascade_ ));
    CascadeMux I__1384 (
            .O(N__14633),
            .I(\POWERLED.pwm_out_en_cascade_ ));
    IoInMux I__1383 (
            .O(N__14630),
            .I(N__14627));
    LocalMux I__1382 (
            .O(N__14627),
            .I(N__14624));
    Odrv4 I__1381 (
            .O(N__14624),
            .I(pwrbtn_led));
    CascadeMux I__1380 (
            .O(N__14621),
            .I(N__14617));
    InMux I__1379 (
            .O(N__14620),
            .I(N__14609));
    InMux I__1378 (
            .O(N__14617),
            .I(N__14609));
    InMux I__1377 (
            .O(N__14616),
            .I(N__14609));
    LocalMux I__1376 (
            .O(N__14609),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    InMux I__1375 (
            .O(N__14606),
            .I(N__14603));
    LocalMux I__1374 (
            .O(N__14603),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__1373 (
            .O(N__14600),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    CascadeMux I__1372 (
            .O(N__14597),
            .I(N__14594));
    InMux I__1371 (
            .O(N__14594),
            .I(N__14591));
    LocalMux I__1370 (
            .O(N__14591),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__1369 (
            .O(N__14588),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__1368 (
            .O(N__14585),
            .I(N__14582));
    LocalMux I__1367 (
            .O(N__14582),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__1366 (
            .O(N__14579),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    CascadeMux I__1365 (
            .O(N__14576),
            .I(N__14573));
    InMux I__1364 (
            .O(N__14573),
            .I(N__14570));
    LocalMux I__1363 (
            .O(N__14570),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__1362 (
            .O(N__14567),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__1361 (
            .O(N__14564),
            .I(N__14561));
    LocalMux I__1360 (
            .O(N__14561),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__1359 (
            .O(N__14558),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    InMux I__1358 (
            .O(N__14555),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    InMux I__1357 (
            .O(N__14552),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__1356 (
            .O(N__14549),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__1355 (
            .O(N__14546),
            .I(N__14543));
    InMux I__1354 (
            .O(N__14543),
            .I(N__14540));
    LocalMux I__1353 (
            .O(N__14540),
            .I(\POWERLED.mult1_un124_sum_i ));
    InMux I__1352 (
            .O(N__14537),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    InMux I__1351 (
            .O(N__14534),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    InMux I__1350 (
            .O(N__14531),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__1349 (
            .O(N__14528),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    InMux I__1348 (
            .O(N__14525),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__1347 (
            .O(N__14522),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    InMux I__1346 (
            .O(N__14519),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__1345 (
            .O(N__14516),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CascadeMux I__1344 (
            .O(N__14513),
            .I(N__14509));
    InMux I__1343 (
            .O(N__14512),
            .I(N__14501));
    InMux I__1342 (
            .O(N__14509),
            .I(N__14501));
    InMux I__1341 (
            .O(N__14508),
            .I(N__14501));
    LocalMux I__1340 (
            .O(N__14501),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    InMux I__1339 (
            .O(N__14498),
            .I(N__14495));
    LocalMux I__1338 (
            .O(N__14495),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__1337 (
            .O(N__14492),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    CascadeMux I__1336 (
            .O(N__14489),
            .I(N__14486));
    InMux I__1335 (
            .O(N__14486),
            .I(N__14483));
    LocalMux I__1334 (
            .O(N__14483),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__1333 (
            .O(N__14480),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__1332 (
            .O(N__14477),
            .I(N__14474));
    LocalMux I__1331 (
            .O(N__14474),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__1330 (
            .O(N__14471),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    CascadeMux I__1329 (
            .O(N__14468),
            .I(N__14465));
    InMux I__1328 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__1327 (
            .O(N__14462),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__1326 (
            .O(N__14459),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__1325 (
            .O(N__14456),
            .I(N__14453));
    LocalMux I__1324 (
            .O(N__14453),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__1323 (
            .O(N__14450),
            .I(N__14444));
    InMux I__1322 (
            .O(N__14449),
            .I(N__14444));
    LocalMux I__1321 (
            .O(N__14444),
            .I(\PCH_PWRGD.count_0_13 ));
    CascadeMux I__1320 (
            .O(N__14441),
            .I(\PCH_PWRGD.countZ0Z_15_cascade_ ));
    InMux I__1319 (
            .O(N__14438),
            .I(N__14433));
    InMux I__1318 (
            .O(N__14437),
            .I(N__14428));
    InMux I__1317 (
            .O(N__14436),
            .I(N__14428));
    LocalMux I__1316 (
            .O(N__14433),
            .I(\PCH_PWRGD.count_rst_1 ));
    LocalMux I__1315 (
            .O(N__14428),
            .I(\PCH_PWRGD.count_rst_1 ));
    InMux I__1314 (
            .O(N__14423),
            .I(N__14417));
    InMux I__1313 (
            .O(N__14422),
            .I(N__14417));
    LocalMux I__1312 (
            .O(N__14417),
            .I(\PCH_PWRGD.count_rst_2 ));
    InMux I__1311 (
            .O(N__14414),
            .I(N__14411));
    LocalMux I__1310 (
            .O(N__14411),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__1309 (
            .O(N__14408),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    InMux I__1308 (
            .O(N__14405),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    InMux I__1307 (
            .O(N__14402),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    InMux I__1306 (
            .O(N__14399),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__1305 (
            .O(N__14396),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__1304 (
            .O(N__14393),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__1303 (
            .O(N__14390),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    InMux I__1302 (
            .O(N__14387),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__1301 (
            .O(N__14384),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__1300 (
            .O(N__14381),
            .I(N__14378));
    LocalMux I__1299 (
            .O(N__14378),
            .I(\PCH_PWRGD.un2_count_1_axb_13 ));
    InMux I__1298 (
            .O(N__14375),
            .I(N__14372));
    LocalMux I__1297 (
            .O(N__14372),
            .I(\PCH_PWRGD.count_0_15 ));
    InMux I__1296 (
            .O(N__14369),
            .I(N__14363));
    InMux I__1295 (
            .O(N__14368),
            .I(N__14363));
    LocalMux I__1294 (
            .O(N__14363),
            .I(\PCH_PWRGD.count_rst ));
    InMux I__1293 (
            .O(N__14360),
            .I(N__14357));
    LocalMux I__1292 (
            .O(N__14357),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    InMux I__1291 (
            .O(N__14354),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    InMux I__1290 (
            .O(N__14351),
            .I(N__14347));
    InMux I__1289 (
            .O(N__14350),
            .I(N__14344));
    LocalMux I__1288 (
            .O(N__14347),
            .I(\PCH_PWRGD.un2_count_1_axb_4 ));
    LocalMux I__1287 (
            .O(N__14344),
            .I(\PCH_PWRGD.un2_count_1_axb_4 ));
    CascadeMux I__1286 (
            .O(N__14339),
            .I(N__14335));
    InMux I__1285 (
            .O(N__14338),
            .I(N__14330));
    InMux I__1284 (
            .O(N__14335),
            .I(N__14330));
    LocalMux I__1283 (
            .O(N__14330),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1282 (
            .O(N__14327),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    InMux I__1281 (
            .O(N__14324),
            .I(N__14318));
    InMux I__1280 (
            .O(N__14323),
            .I(N__14318));
    LocalMux I__1279 (
            .O(N__14318),
            .I(N__14315));
    Odrv4 I__1278 (
            .O(N__14315),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    InMux I__1277 (
            .O(N__14312),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    InMux I__1276 (
            .O(N__14309),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    InMux I__1275 (
            .O(N__14306),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    InMux I__1274 (
            .O(N__14303),
            .I(N__14300));
    LocalMux I__1273 (
            .O(N__14300),
            .I(N__14295));
    InMux I__1272 (
            .O(N__14299),
            .I(N__14290));
    InMux I__1271 (
            .O(N__14298),
            .I(N__14290));
    Odrv4 I__1270 (
            .O(N__14295),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__1269 (
            .O(N__14290),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    CascadeMux I__1268 (
            .O(N__14285),
            .I(N__14281));
    InMux I__1267 (
            .O(N__14284),
            .I(N__14276));
    InMux I__1266 (
            .O(N__14281),
            .I(N__14276));
    LocalMux I__1265 (
            .O(N__14276),
            .I(N__14273));
    Odrv4 I__1264 (
            .O(N__14273),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__1263 (
            .O(N__14270),
            .I(\PCH_PWRGD.un2_count_1_cry_7 ));
    InMux I__1262 (
            .O(N__14267),
            .I(N__14264));
    LocalMux I__1261 (
            .O(N__14264),
            .I(N__14260));
    InMux I__1260 (
            .O(N__14263),
            .I(N__14257));
    Odrv12 I__1259 (
            .O(N__14260),
            .I(\PCH_PWRGD.un2_count_1_axb_9 ));
    LocalMux I__1258 (
            .O(N__14257),
            .I(\PCH_PWRGD.un2_count_1_axb_9 ));
    InMux I__1257 (
            .O(N__14252),
            .I(N__14246));
    InMux I__1256 (
            .O(N__14251),
            .I(N__14246));
    LocalMux I__1255 (
            .O(N__14246),
            .I(N__14243));
    Odrv12 I__1254 (
            .O(N__14243),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    InMux I__1253 (
            .O(N__14240),
            .I(bfn_1_7_0_));
    InMux I__1252 (
            .O(N__14237),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    CascadeMux I__1251 (
            .O(N__14234),
            .I(\PCH_PWRGD.count_rst_9_cascade_ ));
    CascadeMux I__1250 (
            .O(N__14231),
            .I(\PCH_PWRGD.countZ0Z_5_cascade_ ));
    InMux I__1249 (
            .O(N__14228),
            .I(N__14225));
    LocalMux I__1248 (
            .O(N__14225),
            .I(\PCH_PWRGD.count_0_5 ));
    CascadeMux I__1247 (
            .O(N__14222),
            .I(\PCH_PWRGD.count_rst_10_cascade_ ));
    CascadeMux I__1246 (
            .O(N__14219),
            .I(\PCH_PWRGD.un2_count_1_axb_4_cascade_ ));
    InMux I__1245 (
            .O(N__14216),
            .I(N__14213));
    LocalMux I__1244 (
            .O(N__14213),
            .I(\PCH_PWRGD.count_rst_10 ));
    InMux I__1243 (
            .O(N__14210),
            .I(N__14204));
    InMux I__1242 (
            .O(N__14209),
            .I(N__14204));
    LocalMux I__1241 (
            .O(N__14204),
            .I(\PCH_PWRGD.count_0_4 ));
    InMux I__1240 (
            .O(N__14201),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    InMux I__1239 (
            .O(N__14198),
            .I(N__14195));
    LocalMux I__1238 (
            .O(N__14195),
            .I(N__14192));
    Odrv4 I__1237 (
            .O(N__14192),
            .I(\HDA_STRAP.un4_count_10 ));
    CascadeMux I__1236 (
            .O(N__14189),
            .I(\HDA_STRAP.un4_count_cascade_ ));
    InMux I__1235 (
            .O(N__14186),
            .I(N__14183));
    LocalMux I__1234 (
            .O(N__14183),
            .I(\PCH_PWRGD.count_rst_5 ));
    CascadeMux I__1233 (
            .O(N__14180),
            .I(\PCH_PWRGD.count_rst_5_cascade_ ));
    CascadeMux I__1232 (
            .O(N__14177),
            .I(\PCH_PWRGD.un2_count_1_axb_9_cascade_ ));
    InMux I__1231 (
            .O(N__14174),
            .I(N__14168));
    InMux I__1230 (
            .O(N__14173),
            .I(N__14168));
    LocalMux I__1229 (
            .O(N__14168),
            .I(\PCH_PWRGD.count_0_9 ));
    CascadeMux I__1228 (
            .O(N__14165),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__1227 (
            .O(N__14162),
            .I(\PCH_PWRGD.countZ0Z_8_cascade_ ));
    InMux I__1226 (
            .O(N__14159),
            .I(N__14156));
    LocalMux I__1225 (
            .O(N__14156),
            .I(\PCH_PWRGD.count_0_8 ));
    CascadeMux I__1224 (
            .O(N__14153),
            .I(\HDA_STRAP.N_16_cascade_ ));
    InMux I__1223 (
            .O(N__14150),
            .I(N__14147));
    LocalMux I__1222 (
            .O(N__14147),
            .I(\HDA_STRAP.HDA_SDO_ATP_3_0 ));
    InMux I__1221 (
            .O(N__14144),
            .I(N__14140));
    InMux I__1220 (
            .O(N__14143),
            .I(N__14137));
    LocalMux I__1219 (
            .O(N__14140),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    LocalMux I__1218 (
            .O(N__14137),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    CascadeMux I__1217 (
            .O(N__14132),
            .I(\HDA_STRAP.un4_count_9_cascade_ ));
    InMux I__1216 (
            .O(N__14129),
            .I(N__14126));
    LocalMux I__1215 (
            .O(N__14126),
            .I(\HDA_STRAP.un4_count_12 ));
    InMux I__1214 (
            .O(N__14123),
            .I(N__14120));
    LocalMux I__1213 (
            .O(N__14120),
            .I(\HDA_STRAP.un4_count_11 ));
    CascadeMux I__1212 (
            .O(N__14117),
            .I(\HDA_STRAP.un4_count_13_cascade_ ));
    InMux I__1211 (
            .O(N__14114),
            .I(N__14111));
    LocalMux I__1210 (
            .O(N__14111),
            .I(\PCH_PWRGD.delayed_vccin_okZ0 ));
    InMux I__1209 (
            .O(N__14108),
            .I(N__14105));
    LocalMux I__1208 (
            .O(N__14105),
            .I(N__14102));
    Span4Mux_h I__1207 (
            .O(N__14102),
            .I(N__14099));
    Span4Mux_h I__1206 (
            .O(N__14099),
            .I(N__14096));
    Odrv4 I__1205 (
            .O(N__14096),
            .I(gpio_fpga_soc_1));
    InMux I__1204 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__1203 (
            .O(N__14090),
            .I(\HDA_STRAP.m14_i_0 ));
    CascadeMux I__1202 (
            .O(N__14087),
            .I(N__14084));
    InMux I__1201 (
            .O(N__14084),
            .I(N__14069));
    InMux I__1200 (
            .O(N__14083),
            .I(N__14069));
    InMux I__1199 (
            .O(N__14082),
            .I(N__14069));
    InMux I__1198 (
            .O(N__14081),
            .I(N__14069));
    InMux I__1197 (
            .O(N__14080),
            .I(N__14069));
    LocalMux I__1196 (
            .O(N__14069),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    CascadeMux I__1195 (
            .O(N__14066),
            .I(N__14060));
    InMux I__1194 (
            .O(N__14065),
            .I(N__14056));
    InMux I__1193 (
            .O(N__14064),
            .I(N__14047));
    InMux I__1192 (
            .O(N__14063),
            .I(N__14047));
    InMux I__1191 (
            .O(N__14060),
            .I(N__14047));
    InMux I__1190 (
            .O(N__14059),
            .I(N__14047));
    LocalMux I__1189 (
            .O(N__14056),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__1188 (
            .O(N__14047),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    CascadeMux I__1187 (
            .O(N__14042),
            .I(\HDA_STRAP.HDA_SDO_ATP_3_0_cascade_ ));
    IoInMux I__1186 (
            .O(N__14039),
            .I(N__14036));
    LocalMux I__1185 (
            .O(N__14036),
            .I(N__14033));
    Span12Mux_s0_h I__1184 (
            .O(N__14033),
            .I(N__14030));
    Odrv12 I__1183 (
            .O(N__14030),
            .I(hda_sdo_atp));
    CascadeMux I__1182 (
            .O(N__14027),
            .I(N_428_cascade_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_2_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_1_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_7 ),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_15 ),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(COUNTER_un4_counter_7),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    ICE_GB N_92_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18542),
            .GLOBALBUFFEROUTPUT(N_92_g));
    ICE_GB N_557_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__33621),
            .GLOBALBUFFEROUTPUT(N_557_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_LC_1_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_LC_1_1_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(N__14114),
            .in2(_gnd_net_),
            .in3(N__30799),
            .lcout(N_428),
            .ltout(N_428_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_1_1_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_1_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_1_1_1 .LUT_INIT=16'b1111111100001001;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_1_1_1  (
            .in0(N__14065),
            .in1(N__14083),
            .in2(N__14027),
            .in3(N__14093),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34403),
            .ce(N__24047),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIJRUK1_LC_1_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIJRUK1_LC_1_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIJRUK1_LC_1_1_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIJRUK1_LC_1_1_2  (
            .in0(N__16636),
            .in1(N__16678),
            .in2(N__21247),
            .in3(N__16613),
            .lcout(\PCH_PWRGD.delayed_vccin_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_1_1_3 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_1_1_3 .LUT_INIT=16'b0001000100001100;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_0_LC_1_1_3  (
            .in0(N__14108),
            .in1(N__14063),
            .in2(N__15272),
            .in3(N__14082),
            .lcout(\HDA_STRAP.m14_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_1_1_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_1_1_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_1_1_4 .LUT_INIT=16'b0101100011111000;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_1_1_4  (
            .in0(N__14064),
            .in1(N__15270),
            .in2(N__14087),
            .in3(N__25106),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34403),
            .ce(N__24047),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_1_1_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_1_1_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_0_LC_1_1_5  (
            .in0(_gnd_net_),
            .in1(N__14080),
            .in2(_gnd_net_),
            .in3(N__14059),
            .lcout(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIRV1F_2_LC_1_1_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIRV1F_2_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIRV1F_2_LC_1_1_6 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \HDA_STRAP.curr_state_RNIRV1F_2_LC_1_1_6  (
            .in0(N__14081),
            .in1(_gnd_net_),
            .in2(N__14066),
            .in3(N__14143),
            .lcout(\HDA_STRAP.HDA_SDO_ATP_3_0 ),
            .ltout(\HDA_STRAP.HDA_SDO_ATP_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_1_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_1_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_1_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_1_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14042),
            .in3(_gnd_net_),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34403),
            .ce(N__24047),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_1_2_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_1_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNIBJB61_7_LC_1_2_0  (
            .in0(N__14962),
            .in1(N__15034),
            .in2(N__15080),
            .in3(N__14947),
            .lcout(\HDA_STRAP.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_1_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_1_2_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \HDA_STRAP.count_RNIDLB61_6_LC_1_2_1  (
            .in0(N__14932),
            .in1(N__15060),
            .in2(N__14780),
            .in3(N__15376),
            .lcout(\HDA_STRAP.un4_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_1_2_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_1_2_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_1_2_2 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \HDA_STRAP.count_6_LC_1_2_2  (
            .in0(N__14762),
            .in1(N__15262),
            .in2(N__15334),
            .in3(N__14779),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34405),
            .ce(N__24035),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_1_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_1_2_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_1_2_3 .LUT_INIT=16'b0000011101110000;
    LogicCell40 \HDA_STRAP.count_8_LC_1_2_3  (
            .in0(N__15260),
            .in1(N__15320),
            .in2(N__15047),
            .in3(N__15061),
            .lcout(\HDA_STRAP.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34405),
            .ce(N__24035),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_1_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_1_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_1_2_4 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_10_LC_1_2_4  (
            .in0(N__15020),
            .in1(N__15002),
            .in2(N__15333),
            .in3(N__15261),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34405),
            .ce(N__24035),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_1_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_1_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_1_2_5 .LUT_INIT=16'b0000011101110000;
    LogicCell40 \HDA_STRAP.count_11_LC_1_2_5  (
            .in0(N__15259),
            .in1(N__15319),
            .in2(N__14975),
            .in3(N__14993),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34405),
            .ce(N__24035),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_1_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_1_2_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_2_LC_1_2_6  (
            .in0(N__15312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15258),
            .lcout(),
            .ltout(\HDA_STRAP.N_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_1_2_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_1_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_1_2_7 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_1_2_7  (
            .in0(N__14144),
            .in1(N__25107),
            .in2(N__14153),
            .in3(N__14150),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34405),
            .ce(N__24035),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI2L821_2_LC_1_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_1_3_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNI2L821_2_LC_1_3_1  (
            .in0(N__14798),
            .in1(N__14837),
            .in2(N__14819),
            .in3(N__14855),
            .lcout(\HDA_STRAP.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_1_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_1_3_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_1_3_2 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_0_LC_1_3_2  (
            .in0(N__14896),
            .in1(N__15335),
            .in2(N__15338),
            .in3(N__15266),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(N__24039),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_1_3_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_1_3_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \HDA_STRAP.count_RNI4CB61_17_LC_1_3_3  (
            .in0(N__15360),
            .in1(N__14873),
            .in2(N__14900),
            .in3(N__15220),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_1_3_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_1_3_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \HDA_STRAP.count_RNIH7IR1_10_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__14991),
            .in2(N__14132),
            .in3(N__15018),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_1_3_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_1_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIB5IA5_2_LC_1_3_5  (
            .in0(N__14129),
            .in1(N__14123),
            .in2(N__14117),
            .in3(N__14198),
            .lcout(\HDA_STRAP.un4_count ),
            .ltout(\HDA_STRAP.un4_count_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_1_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_1_3_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_1_3_6 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \HDA_STRAP.count_16_LC_1_3_6  (
            .in0(N__15347),
            .in1(N__15336),
            .in2(N__14189),
            .in3(N__15361),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(N__24039),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOV3T1_0_9_LC_1_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOV3T1_0_9_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOV3T1_0_9_LC_1_4_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \PCH_PWRGD.count_RNIOV3T1_0_9_LC_1_4_0  (
            .in0(N__14299),
            .in1(N__14186),
            .in2(N__25572),
            .in3(N__14174),
            .lcout(\PCH_PWRGD.count_1_i_a2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIGD4H1_LC_1_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIGD4H1_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIGD4H1_LC_1_4_1 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNIGD4H1_LC_1_4_1  (
            .in0(N__15796),
            .in1(N__14251),
            .in2(N__25409),
            .in3(N__14263),
            .lcout(\PCH_PWRGD.count_rst_5 ),
            .ltout(\PCH_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOV3T1_9_LC_1_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOV3T1_9_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOV3T1_9_LC_1_4_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIOV3T1_9_LC_1_4_2  (
            .in0(N__25544),
            .in1(_gnd_net_),
            .in2(N__14180),
            .in3(N__14173),
            .lcout(\PCH_PWRGD.un2_count_1_axb_9 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_9_LC_1_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_1_4_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_1_4_3 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.count_9_LC_1_4_3  (
            .in0(N__25385),
            .in1(N__15811),
            .in2(N__14177),
            .in3(N__14252),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34727),
            .ce(N__25566),
            .sr(N__25405));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIFB3H1_LC_1_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIFB3H1_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIFB3H1_LC_1_4_4 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNIFB3H1_LC_1_4_4  (
            .in0(N__14298),
            .in1(N__25380),
            .in2(N__14285),
            .in3(N__15797),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI6A7E3_8_LC_1_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI6A7E3_8_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI6A7E3_8_LC_1_4_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNI6A7E3_8_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(N__14159),
            .in2(N__14165),
            .in3(N__25543),
            .lcout(\PCH_PWRGD.countZ0Z_8 ),
            .ltout(\PCH_PWRGD.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_8_LC_1_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_1_4_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_1_4_6 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.count_8_LC_1_4_6  (
            .in0(N__14284),
            .in1(N__25384),
            .in2(N__14162),
            .in3(N__15798),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34727),
            .ce(N__25566),
            .sr(N__25405));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIPMNB1_LC_1_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIPMNB1_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIPMNB1_LC_1_4_7 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNIPMNB1_LC_1_4_7  (
            .in0(N__15208),
            .in1(N__15812),
            .in2(N__15103),
            .in3(N__25406),
            .lcout(\PCH_PWRGD.count_rst_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIC50H1_LC_1_5_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIC50H1_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIC50H1_LC_1_5_0 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNIC50H1_LC_1_5_0  (
            .in0(N__15792),
            .in1(N__14323),
            .in2(N__25410),
            .in3(N__15186),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI014E3_5_LC_1_5_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI014E3_5_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI014E3_5_LC_1_5_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \PCH_PWRGD.count_RNI014E3_5_LC_1_5_1  (
            .in0(N__25539),
            .in1(N__14228),
            .in2(N__14234),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(\PCH_PWRGD.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_5_LC_1_5_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_1_5_2 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \PCH_PWRGD.count_5_LC_1_5_2  (
            .in0(N__15794),
            .in1(N__25367),
            .in2(N__14231),
            .in3(N__14324),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34700),
            .ce(N__25573),
            .sr(N__25391));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIB3VG1_LC_1_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIB3VG1_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIB3VG1_LC_1_5_3 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNIB3VG1_LC_1_5_3  (
            .in0(N__14350),
            .in1(N__25386),
            .in2(N__14339),
            .in3(N__15793),
            .lcout(\PCH_PWRGD.count_rst_10 ),
            .ltout(\PCH_PWRGD.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIJQ3T1_4_LC_1_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIJQ3T1_4_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIJQ3T1_4_LC_1_5_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PCH_PWRGD.count_RNIJQ3T1_4_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__25538),
            .in2(N__14222),
            .in3(N__14210),
            .lcout(\PCH_PWRGD.un2_count_1_axb_4 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_1_5_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_1_5_5 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_1_5_5 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.count_4_LC_1_5_5  (
            .in0(N__14338),
            .in1(N__25390),
            .in2(N__14219),
            .in3(N__15795),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34700),
            .ce(N__25573),
            .sr(N__25391));
    defparam \PCH_PWRGD.count_RNIJQ3T1_0_4_LC_1_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIJQ3T1_0_4_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIJQ3T1_0_4_LC_1_5_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \PCH_PWRGD.count_RNIJQ3T1_0_4_LC_1_5_6  (
            .in0(N__14216),
            .in1(N__14209),
            .in2(N__25584),
            .in3(N__15393),
            .lcout(\PCH_PWRGD.count_1_i_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_6_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__25621),
            .in2(N__25672),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_1_6_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_1_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_1_6_1  (
            .in0(N__25300),
            .in1(N__15443),
            .in2(_gnd_net_),
            .in3(N__14201),
            .lcout(\PCH_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_6_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__15395),
            .in2(_gnd_net_),
            .in3(N__14354),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_6_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__14351),
            .in2(_gnd_net_),
            .in3(N__14327),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_6_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__15187),
            .in2(_gnd_net_),
            .in3(N__14312),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_6_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__15647),
            .in2(_gnd_net_),
            .in3(N__14309),
            .lcout(\PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_6_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__15137),
            .in2(_gnd_net_),
            .in3(N__14306),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_6_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__14303),
            .in2(_gnd_net_),
            .in3(N__14270),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_7_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__14267),
            .in2(_gnd_net_),
            .in3(N__14240),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIHF5H1_LC_1_7_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIHF5H1_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIHF5H1_LC_1_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNIHF5H1_LC_1_7_1  (
            .in0(N__25298),
            .in1(N__15599),
            .in2(_gnd_net_),
            .in3(N__14237),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_7_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__15107),
            .in2(_gnd_net_),
            .in3(N__14396),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIQOOB1_LC_1_7_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIQOOB1_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIQOOB1_LC_1_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNIQOOB1_LC_1_7_3  (
            .in0(N__25299),
            .in1(N__15541),
            .in2(_gnd_net_),
            .in3(N__14393),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIRQPB1_LC_1_7_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIRQPB1_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIRQPB1_LC_1_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNIRQPB1_LC_1_7_4  (
            .in0(N__25310),
            .in1(N__14381),
            .in2(_gnd_net_),
            .in3(N__14390),
            .lcout(\PCH_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_7_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__15551),
            .in2(_gnd_net_),
            .in3(N__14387),
            .lcout(\PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNITURB1_LC_1_7_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNITURB1_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNITURB1_LC_1_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNITURB1_LC_1_7_6  (
            .in0(N__25311),
            .in1(N__14360),
            .in2(_gnd_net_),
            .in3(N__14384),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_1_7_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_1_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_0_LC_1_7_7  (
            .in0(N__18139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15731),
            .lcout(\PCH_PWRGD.N_38_f0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_15_LC_1_8_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_1_8_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_1_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_15_LC_1_8_0  (
            .in0(N__14369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34740),
            .ce(N__25582),
            .sr(N__25373));
    defparam \PCH_PWRGD.count_RNIU7DH3_13_LC_1_8_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIU7DH3_13_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIU7DH3_13_LC_1_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIU7DH3_13_LC_1_8_1  (
            .in0(N__14450),
            .in1(N__14438),
            .in2(_gnd_net_),
            .in3(N__25549),
            .lcout(\PCH_PWRGD.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_13_LC_1_8_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_13_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14436),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34740),
            .ce(N__25582),
            .sr(N__25373));
    defparam \PCH_PWRGD.count_RNI2EFH3_15_LC_1_8_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI2EFH3_15_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI2EFH3_15_LC_1_8_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNI2EFH3_15_LC_1_8_3  (
            .in0(N__14375),
            .in1(N__25550),
            .in2(_gnd_net_),
            .in3(N__14368),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(\PCH_PWRGD.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIU7DH3_0_13_LC_1_8_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIU7DH3_0_13_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIU7DH3_0_13_LC_1_8_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \PCH_PWRGD.count_RNIU7DH3_0_13_LC_1_8_4  (
            .in0(N__25551),
            .in1(N__14449),
            .in2(N__14441),
            .in3(N__14437),
            .lcout(\PCH_PWRGD.count_1_i_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIS4CH3_12_LC_1_8_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIS4CH3_12_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIS4CH3_12_LC_1_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIS4CH3_12_LC_1_8_5  (
            .in0(N__14423),
            .in1(N__14414),
            .in2(_gnd_net_),
            .in3(N__25548),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_12_LC_1_8_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_1_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_12_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14422),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34740),
            .ce(N__25582),
            .sr(N__25373));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_1_8_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_1_8_7 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_1_8_7  (
            .in0(N__15686),
            .in1(N__15730),
            .in2(N__15838),
            .in3(N__15803),
            .lcout(\PCH_PWRGD.m6_i_i_a2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__22316),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__14508),
            .in2(N__20213),
            .in3(N__14408),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__14498),
            .in2(N__14513),
            .in3(N__14405),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__17046),
            .in2(N__14489),
            .in3(N__14402),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__14477),
            .in2(N__17053),
            .in3(N__14399),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_9_5  (
            .in0(N__18583),
            .in1(N__14512),
            .in2(N__14468),
            .in3(N__14519),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_9_6  (
            .in0(N__14456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14516),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17045),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__22625),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__14658),
            .in2(N__14546),
            .in3(N__14492),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__15914),
            .in2(N__14663),
            .in3(N__14480),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18683),
            .in2(N__15905),
            .in3(N__14471),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__15893),
            .in2(N__18693),
            .in3(N__14459),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5  (
            .in0(N__17044),
            .in1(N__14662),
            .in2(N__16025),
            .in3(N__14552),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__16013),
            .in2(_gnd_net_),
            .in3(N__14549),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_1_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22586),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__22508),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__14616),
            .in2(N__14675),
            .in3(N__14537),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__14606),
            .in2(N__14621),
            .in3(N__14534),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__17079),
            .in2(N__14597),
            .in3(N__14531),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__14585),
            .in2(N__17086),
            .in3(N__14528),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_11_5  (
            .in0(N__17128),
            .in1(N__14620),
            .in2(N__14576),
            .in3(N__14525),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_11_6  (
            .in0(N__14564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14522),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17078),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__22486),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__14697),
            .in2(N__14687),
            .in3(N__14600),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__16070),
            .in2(N__14702),
            .in3(N__14588),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__17309),
            .in2(N__16061),
            .in3(N__14579),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__16046),
            .in2(N__17317),
            .in3(N__14567),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_12_5  (
            .in0(N__17077),
            .in1(N__14701),
            .in2(N__16037),
            .in3(N__14558),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_12_6  (
            .in0(N__16187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14555),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17313),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_1_LC_1_13_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_1_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_1_LC_1_13_0 .LUT_INIT=16'b0011101110111011;
    LogicCell40 \POWERLED.pwm_out_RNO_1_LC_1_13_0  (
            .in0(N__16361),
            .in1(N__21245),
            .in2(N__24696),
            .in3(N__16126),
            .lcout(\POWERLED.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_13_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__22463),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_1_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_1_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_1_13_2  (
            .in0(N__22487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18695),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNIBLUJ_LC_1_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_5_c_RNIBLUJ_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNIBLUJ_LC_1_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNIBLUJ_LC_1_13_6  (
            .in0(N__19181),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(),
            .ltout(\POWERLED.g1_i_a4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIM0E82_4_LC_1_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIM0E82_4_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIM0E82_4_LC_1_13_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_RNIM0E82_4_LC_1_13_7  (
            .in0(N__18917),
            .in1(N__16362),
            .in2(N__14645),
            .in3(N__17462),
            .lcout(\POWERLED.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI9JIT_LC_1_14_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI9JIT_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI9JIT_LC_1_14_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI9JIT_LC_1_14_0  (
            .in0(N__16367),
            .in1(_gnd_net_),
            .in2(N__17249),
            .in3(N__19352),
            .lcout(),
            .ltout(\POWERLED.N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI4GUQ5_LC_1_14_1 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI4GUQ5_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI4GUQ5_LC_1_14_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI4GUQ5_LC_1_14_1  (
            .in0(N__21246),
            .in1(N__14642),
            .in2(N__14636),
            .in3(N__14750),
            .lcout(),
            .ltout(\POWERLED.pwm_out_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNIV9LA6_LC_1_14_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIV9LA6_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIV9LA6_LC_1_14_2 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \POWERLED.pwm_out_RNIV9LA6_LC_1_14_2  (
            .in0(N__16365),
            .in1(_gnd_net_),
            .in2(N__14633),
            .in3(N__14735),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNI48JU1_LC_1_14_4 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_10_c_RNI48JU1_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNI48JU1_LC_1_14_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNI48JU1_LC_1_14_4  (
            .in0(N__16366),
            .in1(N__20777),
            .in2(_gnd_net_),
            .in3(N__17552),
            .lcout(\POWERLED.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_1_14_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_1_14_5 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_1_14_5 .LUT_INIT=16'b1010001110100010;
    LogicCell40 \POWERLED.pwm_out_LC_1_14_5  (
            .in0(N__14734),
            .in1(N__16364),
            .in2(N__14744),
            .in3(N__17245),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34717),
            .ce(),
            .sr(N__16337));
    defparam \POWERLED.curr_state_RNI_0_LC_1_14_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI_0_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI_0_LC_1_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.curr_state_RNI_0_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17267),
            .lcout(\POWERLED.N_2360_i ),
            .ltout(\POWERLED.N_2360_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIPOU53_0_5_LC_1_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIPOU53_0_5_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIPOU53_0_5_LC_1_14_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.count_RNIPOU53_0_5_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14726),
            .in3(N__16127),
            .lcout(\POWERLED.N_660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_1_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_1_15_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_1_15_0  (
            .in0(N__16465),
            .in1(N__16480),
            .in2(N__16436),
            .in3(N__16306),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_1_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_1_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_1_15_1  (
            .in0(N__14714),
            .in1(N__14720),
            .in2(N__14723),
            .in3(N__14708),
            .lcout(VPP_VDDQ_un6_count),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_1_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_1_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_1_15_2  (
            .in0(N__16558),
            .in1(N__16399),
            .in2(N__16418),
            .in3(N__16384),
            .lcout(\VPP_VDDQ.un6_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_1_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_1_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_1_15_3  (
            .in0(N__16231),
            .in1(N__16246),
            .in2(N__16202),
            .in3(N__16261),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_1_15_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_1_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_1_15_6  (
            .in0(N__16216),
            .in1(N__16450),
            .in2(N__16295),
            .in3(N__16276),
            .lcout(\VPP_VDDQ.un6_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_16_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_16_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_1_16_4  (
            .in0(N__32030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14918),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_2_1_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_2_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_0_c_LC_2_1_0  (
            .in0(_gnd_net_),
            .in1(N__14895),
            .in2(N__15337),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_1_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_2_1_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_1_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_2_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_1_LC_2_1_1  (
            .in0(_gnd_net_),
            .in1(N__14869),
            .in2(_gnd_net_),
            .in3(N__14858),
            .lcout(\HDA_STRAP.countZ0Z_1 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_0 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_1 ),
            .clk(N__34463),
            .ce(N__24038),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_2_1_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_2_LC_2_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_2_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_2_LC_2_1_2  (
            .in0(_gnd_net_),
            .in1(N__14854),
            .in2(_gnd_net_),
            .in3(N__14840),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_2 ),
            .clk(N__34463),
            .ce(N__24038),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_2_1_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_3_LC_2_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_2_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_3_LC_2_1_3  (
            .in0(_gnd_net_),
            .in1(N__14836),
            .in2(_gnd_net_),
            .in3(N__14822),
            .lcout(\HDA_STRAP.countZ0Z_3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_3 ),
            .clk(N__34463),
            .ce(N__24038),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_2_1_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_4_LC_2_1_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_2_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_4_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(N__14812),
            .in2(_gnd_net_),
            .in3(N__14801),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_4 ),
            .clk(N__34463),
            .ce(N__24038),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_2_1_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_5_LC_2_1_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_2_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_5_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(N__14797),
            .in2(_gnd_net_),
            .in3(N__14783),
            .lcout(\HDA_STRAP.countZ0Z_5 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_5 ),
            .clk(N__34463),
            .ce(N__24038),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_2_1_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_2_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_2_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_2_1_6  (
            .in0(_gnd_net_),
            .in1(N__14775),
            .in2(_gnd_net_),
            .in3(N__14753),
            .lcout(\HDA_STRAP.un1_count_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_5 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_2_1_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_7_LC_2_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_2_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_7_LC_2_1_7  (
            .in0(_gnd_net_),
            .in1(N__15076),
            .in2(_gnd_net_),
            .in3(N__15065),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_7 ),
            .clk(N__34463),
            .ce(N__24038),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_2_2_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_2_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__15062),
            .in2(_gnd_net_),
            .in3(N__15038),
            .lcout(\HDA_STRAP.un1_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_2_2_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_9_LC_2_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_2_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_9_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__15035),
            .in2(_gnd_net_),
            .in3(N__15023),
            .lcout(\HDA_STRAP.countZ0Z_9 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_8 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_9 ),
            .clk(N__34404),
            .ce(N__24036),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_2_2_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_2_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_2_2_2  (
            .in0(_gnd_net_),
            .in1(N__15019),
            .in2(_gnd_net_),
            .in3(N__14996),
            .lcout(\HDA_STRAP.un1_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_2_2_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_2_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_2_2_3  (
            .in0(_gnd_net_),
            .in1(N__14992),
            .in2(_gnd_net_),
            .in3(N__14966),
            .lcout(\HDA_STRAP.un1_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_2_2_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_12_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_2_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_12_LC_2_2_4  (
            .in0(_gnd_net_),
            .in1(N__14963),
            .in2(_gnd_net_),
            .in3(N__14951),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_12 ),
            .clk(N__34404),
            .ce(N__24036),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_2_2_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_13_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_2_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_13_LC_2_2_5  (
            .in0(_gnd_net_),
            .in1(N__14948),
            .in2(_gnd_net_),
            .in3(N__14936),
            .lcout(\HDA_STRAP.countZ0Z_13 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_13 ),
            .clk(N__34404),
            .ce(N__24036),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_2_2_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_14_LC_2_2_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_2_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_14_LC_2_2_6  (
            .in0(_gnd_net_),
            .in1(N__14933),
            .in2(_gnd_net_),
            .in3(N__14921),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_14 ),
            .clk(N__34404),
            .ce(N__24036),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_2_2_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_15_LC_2_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_2_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_15_LC_2_2_7  (
            .in0(_gnd_net_),
            .in1(N__15377),
            .in2(_gnd_net_),
            .in3(N__15365),
            .lcout(\HDA_STRAP.countZ0Z_15 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_15 ),
            .clk(N__34404),
            .ce(N__24036),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_2_3_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_2_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(N__15362),
            .in2(_gnd_net_),
            .in3(N__15341),
            .lcout(\HDA_STRAP.un1_count_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_2_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_2_3_1 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \HDA_STRAP.count_17_LC_2_3_1  (
            .in0(N__15329),
            .in1(N__15221),
            .in2(N__15271),
            .in3(N__15224),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34464),
            .ce(N__24037),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_11_LC_2_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_2_4_0 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \PCH_PWRGD.count_11_LC_2_4_0  (
            .in0(N__15096),
            .in1(N__25392),
            .in2(N__15209),
            .in3(N__15800),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__25560),
            .sr(N__25365));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIE92H1_LC_2_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIE92H1_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIE92H1_LC_2_4_1 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNIE92H1_LC_2_4_1  (
            .in0(N__15801),
            .in1(N__15167),
            .in2(N__25412),
            .in3(N__15133),
            .lcout(\PCH_PWRGD.count_rst_7 ),
            .ltout(\PCH_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIMT3T1_0_7_LC_2_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMT3T1_0_7_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMT3T1_0_7_LC_2_4_2 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \PCH_PWRGD.count_RNIMT3T1_0_7_LC_2_4_2  (
            .in0(N__25561),
            .in1(N__15188),
            .in2(N__15170),
            .in3(N__15146),
            .lcout(\PCH_PWRGD.count_1_i_a2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_7_LC_2_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_2_4_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_2_4_3 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \PCH_PWRGD.count_7_LC_2_4_3  (
            .in0(N__15799),
            .in1(N__15166),
            .in2(N__25411),
            .in3(N__15132),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__25560),
            .sr(N__25365));
    defparam \PCH_PWRGD.count_RNIMT3T1_7_LC_2_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMT3T1_7_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMT3T1_7_LC_2_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIMT3T1_7_LC_2_4_4  (
            .in0(N__15152),
            .in1(N__15145),
            .in2(_gnd_net_),
            .in3(N__25541),
            .lcout(\PCH_PWRGD.un2_count_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQ1BH3_11_LC_2_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQ1BH3_11_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQ1BH3_11_LC_2_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PCH_PWRGD.count_RNIQ1BH3_11_LC_2_4_5  (
            .in0(N__25540),
            .in1(N__15119),
            .in2(_gnd_net_),
            .in3(N__15113),
            .lcout(\PCH_PWRGD.countZ0Z_11 ),
            .ltout(\PCH_PWRGD.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIGN3T1_0_1_LC_2_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIGN3T1_0_1_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIGN3T1_0_1_LC_2_4_6 .LUT_INIT=16'b0011000001010000;
    LogicCell40 \PCH_PWRGD.count_RNIGN3T1_0_1_LC_2_4_6  (
            .in0(N__25610),
            .in1(N__15629),
            .in2(N__15437),
            .in3(N__25542),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIHFFK7_1_LC_2_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHFFK7_1_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHFFK7_1_LC_2_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIHFFK7_1_LC_2_4_7  (
            .in0(N__15434),
            .in1(N__15428),
            .in2(N__15422),
            .in3(N__15419),
            .lcout(\PCH_PWRGD.count_1_i_a2_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI1TUH1_0_LC_2_5_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI1TUH1_0_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI1TUH1_0_LC_2_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNI1TUH1_0_LC_2_5_0  (
            .in0(N__15881),
            .in1(N__15407),
            .in2(_gnd_net_),
            .in3(N__24668),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_5_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_5_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15413),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2226_i ),
            .ltout(\PCH_PWRGD.N_2226_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_5_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_5_2 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_5_2  (
            .in0(N__15839),
            .in1(N__16677),
            .in2(N__15410),
            .in3(N__15780),
            .lcout(\PCH_PWRGD.curr_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI22GO8_1_LC_2_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI22GO8_1_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI22GO8_1_LC_2_5_3 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \PCH_PWRGD.count_RNI22GO8_1_LC_2_5_3  (
            .in0(N__15496),
            .in1(N__25663),
            .in2(N__15515),
            .in3(N__25401),
            .lcout(\PCH_PWRGD.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIHFFK7_0_1_LC_2_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHFFK7_0_1_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHFFK7_0_1_LC_2_5_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \PCH_PWRGD.count_RNIHFFK7_0_1_LC_2_5_4  (
            .in0(N__25664),
            .in1(N__15511),
            .in2(_gnd_net_),
            .in3(N__15495),
            .lcout(\PCH_PWRGD.N_386 ),
            .ltout(\PCH_PWRGD.N_386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIA1UG1_LC_2_5_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIA1UG1_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIA1UG1_LC_2_5_5 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNIA1UG1_LC_2_5_5  (
            .in0(N__15571),
            .in1(N__25402),
            .in2(N__15401),
            .in3(N__15394),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISQ1E3_3_LC_2_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISQ1E3_3_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISQ1E3_3_LC_2_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNISQ1E3_3_LC_2_5_6  (
            .in0(N__25571),
            .in1(_gnd_net_),
            .in2(N__15398),
            .in3(N__15557),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(\PCH_PWRGD.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_3_LC_2_5_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_2_5_7 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \PCH_PWRGD.count_3_LC_2_5_7  (
            .in0(N__15572),
            .in1(N__15802),
            .in2(N__15560),
            .in3(N__25399),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34699),
            .ce(N__25570),
            .sr(N__25400));
    defparam \PCH_PWRGD.count_2_LC_2_6_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_2_6_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \PCH_PWRGD.count_2_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__15463),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34540),
            .ce(N__25562),
            .sr(N__25366));
    defparam \PCH_PWRGD.count_RNI0BEH3_14_LC_2_6_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI0BEH3_14_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI0BEH3_14_LC_2_6_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \PCH_PWRGD.count_RNI0BEH3_14_LC_2_6_1  (
            .in0(N__15481),
            .in1(N__25295),
            .in2(N__15473),
            .in3(N__25534),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(\PCH_PWRGD.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQN0E3_0_2_LC_2_6_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQN0E3_0_2_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQN0E3_0_2_LC_2_6_2 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \PCH_PWRGD.count_RNIQN0E3_0_2_LC_2_6_2  (
            .in0(N__25537),
            .in1(N__15462),
            .in2(N__15545),
            .in3(N__15452),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI9P6MA_2_LC_2_6_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI9P6MA_2_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI9P6MA_2_LC_2_6_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI9P6MA_2_LC_2_6_3  (
            .in0(N__15542),
            .in1(N__15638),
            .in2(N__15527),
            .in3(N__15524),
            .lcout(\PCH_PWRGD.count_1_i_a2_11_0 ),
            .ltout(\PCH_PWRGD.count_1_i_a2_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_2_6_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_2_6_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \PCH_PWRGD.count_0_LC_2_6_4  (
            .in0(N__25296),
            .in1(N__25662),
            .in2(N__15503),
            .in3(N__15500),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34540),
            .ce(N__25562),
            .sr(N__25366));
    defparam \PCH_PWRGD.count_14_LC_2_6_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_2_6_5 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_2_6_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \PCH_PWRGD.count_14_LC_2_6_5  (
            .in0(N__15482),
            .in1(N__25297),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34540),
            .ce(N__25562),
            .sr(N__25366));
    defparam \PCH_PWRGD.count_RNIQN0E3_2_LC_2_6_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQN0E3_2_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQN0E3_2_LC_2_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PCH_PWRGD.count_RNIQN0E3_2_LC_2_6_6  (
            .in0(N__25535),
            .in1(N__15464),
            .in2(_gnd_net_),
            .in3(N__15451),
            .lcout(\PCH_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIHOJLA_0_LC_2_6_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHOJLA_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHOJLA_0_LC_2_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIHOJLA_0_LC_2_6_7  (
            .in0(N__15662),
            .in1(N__15656),
            .in2(_gnd_net_),
            .in3(N__25536),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIHI041_0_LC_2_7_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIHI041_0_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIHI041_0_LC_2_7_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIHI041_0_LC_2_7_0  (
            .in0(N__15727),
            .in1(N__15684),
            .in2(_gnd_net_),
            .in3(N__24620),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(\PCH_PWRGD.count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI245E3_6_LC_2_7_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI245E3_6_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI245E3_6_LC_2_7_1 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \PCH_PWRGD.count_RNI245E3_6_LC_2_7_1  (
            .in0(N__15605),
            .in1(N__25467),
            .in2(N__15650),
            .in3(N__15613),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(\PCH_PWRGD.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIHPOM3_0_10_LC_2_7_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHPOM3_0_10_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHPOM3_0_10_LC_2_7_2 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \PCH_PWRGD.count_RNIHPOM3_0_10_LC_2_7_2  (
            .in0(N__25469),
            .in1(N__15591),
            .in2(N__15641),
            .in3(N__15581),
            .lcout(\PCH_PWRGD.count_1_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIGN3T1_1_LC_2_7_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIGN3T1_1_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIGN3T1_1_LC_2_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIGN3T1_1_LC_2_7_3  (
            .in0(N__15625),
            .in1(N__25606),
            .in2(_gnd_net_),
            .in3(N__25586),
            .lcout(\PCH_PWRGD.un2_count_1_axb_1 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIHI041_1_LC_2_7_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHI041_1_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHI041_1_LC_2_7_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \PCH_PWRGD.count_RNIHI041_1_LC_2_7_4  (
            .in0(N__25404),
            .in1(_gnd_net_),
            .in2(N__15632),
            .in3(N__25665),
            .lcout(\PCH_PWRGD.count_rst_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_6_LC_2_7_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_2_7_5 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_2_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PCH_PWRGD.count_6_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__15614),
            .in2(_gnd_net_),
            .in3(N__25312),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(N__25585),
            .sr(N__25403));
    defparam \PCH_PWRGD.count_RNIHPOM3_10_LC_2_7_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHPOM3_10_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHPOM3_10_LC_2_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PCH_PWRGD.count_RNIHPOM3_10_LC_2_7_6  (
            .in0(N__25468),
            .in1(N__15593),
            .in2(_gnd_net_),
            .in3(N__15580),
            .lcout(\PCH_PWRGD.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_10_LC_2_7_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_2_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_10_LC_2_7_7  (
            .in0(N__15592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(N__25585),
            .sr(N__25403));
    defparam \PCH_PWRGD.curr_state_0_LC_2_8_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_2_8_0 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_2_8_0  (
            .in0(N__15831),
            .in1(N__15728),
            .in2(N__16676),
            .in3(N__15805),
            .lcout(\PCH_PWRGD.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34551),
            .ce(N__21206),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_8_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_8_1 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_8_1  (
            .in0(N__15866),
            .in1(_gnd_net_),
            .in2(N__30810),
            .in3(N__15872),
            .lcout(\PCH_PWRGD.N_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_8_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15830),
            .lcout(\PCH_PWRGD.N_2244_i ),
            .ltout(\PCH_PWRGD.N_2244_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_1_LC_2_8_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_1_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI3DJU_0_1_LC_2_8_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI3DJU_0_1_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__15865),
            .in2(N__15851),
            .in3(N__30800),
            .lcout(\PCH_PWRGD.N_655 ),
            .ltout(\PCH_PWRGD.N_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_8_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_8_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15848),
            .in3(N__18124),
            .lcout(\PCH_PWRGD.curr_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_2_8_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_2_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_2_8_6  (
            .in0(N__15668),
            .in1(N__15845),
            .in2(_gnd_net_),
            .in3(N__24667),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_2_8_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_2_8_7 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_2_8_7  (
            .in0(N__15804),
            .in1(N__15729),
            .in2(N__15689),
            .in3(N__15685),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34551),
            .ce(N__21206),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_2_9_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_2_9_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_2_9_1  (
            .in0(N__16768),
            .in1(N__16732),
            .in2(_gnd_net_),
            .in3(N__16697),
            .lcout(\VPP_VDDQ.N_64_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_2_9_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_2_9_2 .LUT_INIT=16'b0101001101010000;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_2_9_2  (
            .in0(N__15932),
            .in1(N__16702),
            .in2(N__16741),
            .in3(N__16771),
            .lcout(VPP_VDDQ_curr_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34651),
            .ce(N__24048),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_2_9_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_2_9_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__21313),
            .in2(_gnd_net_),
            .in3(N__32021),
            .lcout(N_626),
            .ltout(N_626_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_30_0_LC_2_9_4 .C_ON=1'b0;
    defparam \POWERLED.G_30_0_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_30_0_LC_2_9_4 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \POWERLED.G_30_0_LC_2_9_4  (
            .in0(N__16731),
            .in1(N__16769),
            .in2(N__15938),
            .in3(N__24132),
            .lcout(),
            .ltout(\POWERLED.G_30Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_30_LC_2_9_5 .C_ON=1'b0;
    defparam \POWERLED.G_30_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_30_LC_2_9_5 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \POWERLED.G_30_LC_2_9_5  (
            .in0(N__16770),
            .in1(N__16733),
            .in2(N__15935),
            .in3(N__15931),
            .lcout(G_30),
            .ltout(G_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_2_9_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_2_9_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15917),
            .in3(N__24133),
            .lcout(\VPP_VDDQ.N_92_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_2_9_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_2_9_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__16734),
            .in2(_gnd_net_),
            .in3(N__16698),
            .lcout(VPP_VDDQ_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34651),
            .ce(N__24048),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__22585),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__25130),
            .in2(N__18500),
            .in3(N__15908),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__15992),
            .in2(N__16001),
            .in3(N__15896),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__25154),
            .in2(N__15974),
            .in3(N__15884),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__15956),
            .in2(N__25164),
            .in3(N__16016),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_10_5  (
            .in0(N__18682),
            .in1(N__25190),
            .in2(N__25207),
            .in3(N__16007),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_10_6  (
            .in0(N__16103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16004),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_2_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_2_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_2_10_7  (
            .in0(N__15991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25153),
            .lcout(\POWERLED.mult1_un124_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__22532),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__16080),
            .in2(N__17282),
            .in3(N__15983),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__15980),
            .in2(N__16085),
            .in3(N__15965),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__15962),
            .in2(N__17137),
            .in3(N__15950),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__17133),
            .in2(N__15947),
            .in3(N__16115),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_11_5  (
            .in0(N__25152),
            .in1(N__16084),
            .in2(N__16112),
            .in3(N__16097),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_11_6  (
            .in0(N__16094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16088),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_11_7  (
            .in0(N__17129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__22462),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__16171),
            .in2(N__18515),
            .in3(N__16064),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__18872),
            .in2(N__16175),
            .in3(N__16049),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__18854),
            .in2(N__18767),
            .in3(N__16040),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__18766),
            .in2(N__18833),
            .in3(N__16028),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_12_5  (
            .in0(N__17308),
            .in1(N__16170),
            .in2(N__18812),
            .in3(N__16181),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_12_6  (
            .in0(N__18788),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16178),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_12_7  (
            .in0(N__18762),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNISDGE_LC_2_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_4_c_RNISDGE_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNISDGE_LC_2_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNISDGE_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__19179),
            .in2(_gnd_net_),
            .in3(N__18915),
            .lcout(\POWERLED.count_1_5 ),
            .ltout(\POWERLED.count_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGTVS_5_LC_2_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGTVS_5_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGTVS_5_LC_2_13_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIGTVS_5_LC_2_13_1  (
            .in0(N__24611),
            .in1(_gnd_net_),
            .in2(N__16160),
            .in3(N__16155),
            .lcout(\POWERLED.un1_count_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGTVS_1_5_LC_2_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGTVS_1_5_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGTVS_1_5_LC_2_13_2 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \POWERLED.count_RNIGTVS_1_5_LC_2_13_2  (
            .in0(N__17012),
            .in1(N__16157),
            .in2(N__16142),
            .in3(N__24616),
            .lcout(\POWERLED.count_RNIGTVS_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_2_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_2_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_5_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__19180),
            .in2(_gnd_net_),
            .in3(N__18916),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34715),
            .ce(N__21214),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGTVS_0_5_LC_2_13_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGTVS_0_5_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGTVS_0_5_LC_2_13_5 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \POWERLED.count_RNIGTVS_0_5_LC_2_13_5  (
            .in0(N__16156),
            .in1(N__16138),
            .in2(N__24676),
            .in3(N__19412),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIPOU53_5_LC_2_13_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIPOU53_5_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIPOU53_5_LC_2_13_6 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \POWERLED.count_RNIPOU53_5_LC_2_13_6  (
            .in0(N__20447),
            .in1(N__17461),
            .in2(N__16130),
            .in3(N__17564),
            .lcout(\POWERLED.un79_clk_100khz ),
            .ltout(\POWERLED.un79_clk_100khz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_2_13_7 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_2_13_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_2_13_7  (
            .in0(N__24615),
            .in1(_gnd_net_),
            .in2(N__16370),
            .in3(N__16363),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_2_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_2_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_2_14_0  (
            .in0(N__24156),
            .in1(N__16307),
            .in2(N__16325),
            .in3(N__16324),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_1_LC_2_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_2_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_2_14_1  (
            .in0(N__24152),
            .in1(N__16294),
            .in2(_gnd_net_),
            .in3(N__16280),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_2_LC_2_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_2_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_2_14_2  (
            .in0(N__24157),
            .in1(N__16277),
            .in2(_gnd_net_),
            .in3(N__16265),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_3_LC_2_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_2_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_2_14_3  (
            .in0(N__24153),
            .in1(N__16262),
            .in2(_gnd_net_),
            .in3(N__16250),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_4_LC_2_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_2_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_2_14_4  (
            .in0(N__24158),
            .in1(N__16247),
            .in2(_gnd_net_),
            .in3(N__16235),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_5_LC_2_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_2_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_2_14_5  (
            .in0(N__24154),
            .in1(N__16232),
            .in2(_gnd_net_),
            .in3(N__16220),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_6_LC_2_14_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_2_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_2_14_6  (
            .in0(N__24159),
            .in1(N__16217),
            .in2(_gnd_net_),
            .in3(N__16205),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_7_LC_2_14_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_2_14_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_2_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_2_14_7  (
            .in0(N__24155),
            .in1(N__16201),
            .in2(_gnd_net_),
            .in3(N__16484),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__34660),
            .ce(),
            .sr(N__16530));
    defparam \VPP_VDDQ.count_8_LC_2_15_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_2_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_2_15_0  (
            .in0(N__24166),
            .in1(N__16481),
            .in2(_gnd_net_),
            .in3(N__16469),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.count_9_LC_2_15_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_2_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_2_15_1  (
            .in0(N__24162),
            .in1(N__16466),
            .in2(_gnd_net_),
            .in3(N__16454),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.count_10_LC_2_15_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_2_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_2_15_2  (
            .in0(N__24163),
            .in1(N__16451),
            .in2(_gnd_net_),
            .in3(N__16439),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.count_11_LC_2_15_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_2_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_2_15_3  (
            .in0(N__24160),
            .in1(N__16435),
            .in2(_gnd_net_),
            .in3(N__16421),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.count_12_LC_2_15_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_2_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_2_15_4  (
            .in0(N__24164),
            .in1(N__16417),
            .in2(_gnd_net_),
            .in3(N__16403),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.count_13_LC_2_15_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_2_15_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_2_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_2_15_5  (
            .in0(N__24161),
            .in1(N__16400),
            .in2(_gnd_net_),
            .in3(N__16388),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.count_14_LC_2_15_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_2_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_2_15_6  (
            .in0(N__24165),
            .in1(N__16385),
            .in2(_gnd_net_),
            .in3(N__16373),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__34726),
            .ce(),
            .sr(N__16532));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__23167),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_2_16_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_2_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__16559),
            .in2(_gnd_net_),
            .in3(N__16562),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34718),
            .ce(N__16547),
            .sr(N__16531));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_4_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_4_1_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_4_1_0  (
            .in0(N__21482),
            .in1(N__20997),
            .in2(N__17734),
            .in3(N__21703),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_4_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_4_1_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIPM861_8_LC_4_1_1  (
            .in0(_gnd_net_),
            .in1(N__19979),
            .in2(N__16502),
            .in3(N__16499),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_8_LC_4_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_8_LC_4_1_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_4_1_2  (
            .in0(N__21485),
            .in1(N__21698),
            .in2(N__17735),
            .in3(N__21000),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34539),
            .ce(N__20046),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_4_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_9_LC_4_1_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_4_1_3  (
            .in0(N__17717),
            .in1(N__21057),
            .in2(N__21719),
            .in3(N__21486),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34539),
            .ce(N__20046),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_4_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_4_1_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_4_1_4  (
            .in0(N__21483),
            .in1(N__17716),
            .in2(N__21718),
            .in3(N__20998),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_4_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_4_1_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIRP961_9_LC_4_1_5  (
            .in0(_gnd_net_),
            .in1(N__19980),
            .in2(N__16493),
            .in3(N__16490),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_10_LC_4_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_4_1_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_10_LC_4_1_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_4_1_6  (
            .in0(N__21484),
            .in1(N__20999),
            .in2(N__17702),
            .in3(N__21702),
            .lcout(\VPP_VDDQ.count_2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34539),
            .ce(N__20046),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_4_2_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_4_2_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_4_2_0  (
            .in0(N__21538),
            .in1(N__21714),
            .in2(N__21063),
            .in3(N__17899),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_4_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_4_2_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJ48C1_14_LC_4_2_1  (
            .in0(_gnd_net_),
            .in1(N__16784),
            .in2(N__16586),
            .in3(N__20029),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_4_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_4_2_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_4_2_2  (
            .in0(N__17614),
            .in1(N__21536),
            .in2(N__21062),
            .in3(N__21713),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_4_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_4_2_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIHA461_4_LC_4_2_3  (
            .in0(_gnd_net_),
            .in1(N__16580),
            .in2(N__16583),
            .in3(N__20028),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_4_LC_4_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_4_LC_4_2_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_4_2_4  (
            .in0(N__17615),
            .in1(N__21537),
            .in2(N__21065),
            .in3(N__21717),
            .lcout(\VPP_VDDQ.count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34265),
            .ce(N__20035),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_5_LC_4_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_5_LC_4_2_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_4_2_5  (
            .in0(N__21716),
            .in1(N__21540),
            .in2(N__17588),
            .in3(N__21047),
            .lcout(\VPP_VDDQ.count_2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34265),
            .ce(N__20035),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_4_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_4_2_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_4_2_6  (
            .in0(N__21539),
            .in1(N__17584),
            .in2(N__21064),
            .in3(N__21715),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_4_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_4_2_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJD561_5_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(N__16574),
            .in2(N__16568),
            .in3(N__20030),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_4_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_4_3_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIH17C1_13_LC_4_3_0  (
            .in0(N__16790),
            .in1(N__20027),
            .in2(_gnd_net_),
            .in3(N__17840),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_4_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_4_3_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_4_3_1  (
            .in0(N__21709),
            .in1(N__21547),
            .in2(N__21059),
            .in3(N__17671),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_4_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_4_3_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIFU5C1_12_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__16796),
            .in2(N__16565),
            .in3(N__20026),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_15_LC_4_3_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_4_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_15_LC_4_3_3  (
            .in0(N__17885),
            .in1(N__17660),
            .in2(N__16799),
            .in3(N__17915),
            .lcout(\VPP_VDDQ.un9_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_12_LC_4_3_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_12_LC_4_3_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_4_3_5  (
            .in0(N__21710),
            .in1(N__21549),
            .in2(N__21060),
            .in3(N__17672),
            .lcout(\VPP_VDDQ.count_2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34354),
            .ce(N__20034),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_13_LC_4_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_13_LC_4_3_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_4_3_6  (
            .in0(N__21548),
            .in1(N__21028),
            .in2(N__17855),
            .in3(N__21712),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34354),
            .ce(N__20034),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_14_LC_4_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_14_LC_4_3_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_4_3_7  (
            .in0(N__21711),
            .in1(N__21550),
            .in2(N__21061),
            .in3(N__17900),
            .lcout(\VPP_VDDQ.count_2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34354),
            .ce(N__20034),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_0 .LUT_INIT=16'b0000100111101001;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_0  (
            .in0(N__16750),
            .in1(N__32880),
            .in2(N__24167),
            .in3(N__16778),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_1 .LUT_INIT=16'b1110001111000010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_1  (
            .in0(N__32881),
            .in1(N__16751),
            .in2(N__16712),
            .in3(N__16709),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_4_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_4_4_4  (
            .in0(N__16679),
            .in1(N__16637),
            .in2(N__21248),
            .in3(N__16609),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_4_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_4_4_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_4_4_6  (
            .in0(N__21545),
            .in1(N__17695),
            .in2(N__21058),
            .in3(N__21708),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_4_4_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_4_4_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI4TU51_10_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__16595),
            .in2(N__16826),
            .in3(N__20025),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_4_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_4_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__17947),
            .in2(N__18173),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__18003),
            .in2(_gnd_net_),
            .in3(N__16823),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__18034),
            .in2(_gnd_net_),
            .in3(N__16820),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__17977),
            .in2(_gnd_net_),
            .in3(N__16817),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__17930),
            .in2(_gnd_net_),
            .in3(N__16814),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__18345),
            .in2(_gnd_net_),
            .in3(N__16811),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_4_5_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_4_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__17960),
            .in2(_gnd_net_),
            .in3(N__16808),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__34491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_4_5_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_4_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(N__18326),
            .in2(_gnd_net_),
            .in3(N__16805),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__34491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_4_6_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_4_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__18287),
            .in2(_gnd_net_),
            .in3(N__16802),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_4_6_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_4_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__18301),
            .in2(_gnd_net_),
            .in3(N__16853),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_4_6_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_4_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__18314),
            .in2(_gnd_net_),
            .in3(N__16850),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_4_6_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_4_6_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_4_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__18275),
            .in2(_gnd_net_),
            .in3(N__16847),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_4_6_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_4_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(N__18250),
            .in2(_gnd_net_),
            .in3(N__16844),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_4_6_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_4_6_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_4_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__18236),
            .in2(_gnd_net_),
            .in3(N__16841),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_4_6_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_4_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__18263),
            .in2(_gnd_net_),
            .in3(N__16838),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_4_6_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_4_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(N__18224),
            .in2(_gnd_net_),
            .in3(N__16835),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__34550),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_4_7_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_4_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__18185),
            .in2(_gnd_net_),
            .in3(N__16832),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_4_7_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_4_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__18212),
            .in2(_gnd_net_),
            .in3(N__16829),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_4_7_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_4_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__18199),
            .in2(_gnd_net_),
            .in3(N__16880),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_4_7_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_4_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__18476),
            .in2(_gnd_net_),
            .in3(N__16877),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_4_7_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_4_7_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_4_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__18463),
            .in2(_gnd_net_),
            .in3(N__16874),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_4_7_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_4_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(N__18488),
            .in2(_gnd_net_),
            .in3(N__16871),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_4_7_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_4_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__18449),
            .in2(_gnd_net_),
            .in3(N__16868),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_4_7_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_4_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(N__18079),
            .in2(_gnd_net_),
            .in3(N__16865),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__34495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_4_8_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_4_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(N__18065),
            .in2(_gnd_net_),
            .in3(N__16862),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_4_8_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_4_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(N__18092),
            .in2(_gnd_net_),
            .in3(N__16859),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_4_8_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_4_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__18104),
            .in2(_gnd_net_),
            .in3(N__16856),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_4_8_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_4_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__16904),
            .in2(_gnd_net_),
            .in3(N__16949),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_4_8_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_4_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__16915),
            .in2(_gnd_net_),
            .in3(N__16946),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_4_8_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_4_8_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_30_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16937),
            .in3(N__16943),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_4_8_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_4_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.counter_31_LC_4_8_6  (
            .in0(N__16925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16940),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34600),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_4_8_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_4_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_4_8_7  (
            .in0(N__16933),
            .in1(N__16924),
            .in2(N__16916),
            .in3(N__16903),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_9_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__16895),
            .in2(N__20135),
            .in3(N__19064),
            .lcout(\POWERLED.N_4842_i ),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_9_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__17378),
            .in2(N__17395),
            .in3(N__22133),
            .lcout(\POWERLED.mult1_un159_sum_i_8 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_9_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__17183),
            .in2(N__17200),
            .in3(N__22241),
            .lcout(\POWERLED.mult1_un152_sum_i_8 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_9_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__20120),
            .in2(N__16889),
            .in3(N__18995),
            .lcout(\POWERLED.count_i_3 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_9_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__17411),
            .in2(N__17444),
            .in3(N__18595),
            .lcout(\POWERLED.mult1_un138_sum_i_8 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_9_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_9_5  (
            .in0(N__17057),
            .in1(N__17024),
            .in2(N__17008),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_8 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_9_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_9_6  (
            .in0(N__19411),
            .in1(N__18659),
            .in2(N__16991),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_6 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_9_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__16982),
            .in2(N__17150),
            .in3(N__20762),
            .lcout(\POWERLED.N_4841_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_10_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_10_0  (
            .in0(N__20519),
            .in1(N__16976),
            .in2(N__17108),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_8 ),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_10_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__16970),
            .in2(N__17330),
            .in3(N__20489),
            .lcout(\POWERLED.N_4849_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_10_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__17288),
            .in2(N__16964),
            .in3(N__19280),
            .lcout(\POWERLED.count_i_10 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_10_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_10_3  (
            .in0(N__19250),
            .in1(N__16955),
            .in2(N__17099),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_11 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_10_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_10_4  (
            .in0(N__18736),
            .in1(N__20612),
            .in2(N__20629),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_10_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_10_5  (
            .in0(N__20582),
            .in1(N__17171),
            .in2(N__20276),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4851_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_10_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_10_6  (
            .in0(N__20806),
            .in1(N__17165),
            .in2(N__18533),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4855_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_10_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_10_7  (
            .in0(N__20843),
            .in1(N__17159),
            .in2(N__18524),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4856_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_11_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17153),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_11_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25165),
            .lcout(\POWERLED.mult1_un117_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_11_2  (
            .in0(N__17138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18754),
            .lcout(\POWERLED.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17090),
            .lcout(\POWERLED.mult1_un103_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_11_5  (
            .in0(N__17321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22507),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_4_12_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_4_12_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_4_12_0  (
            .in0(N__17263),
            .in1(N__17365),
            .in2(_gnd_net_),
            .in3(N__17232),
            .lcout(),
            .ltout(\POWERLED.N_437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNICO541_0_LC_4_12_1 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNICO541_0_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNICO541_0_LC_4_12_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.curr_state_RNICO541_0_LC_4_12_1  (
            .in0(N__24555),
            .in1(_gnd_net_),
            .in2(N__17270),
            .in3(N__17216),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(\POWERLED.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_4_12_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_4_12_2 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \POWERLED.curr_state_0_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__17233),
            .in2(N__17219),
            .in3(N__17361),
            .lcout(\POWERLED.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34680),
            .ce(N__21211),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_4_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_4_12_3 .LUT_INIT=16'b0000101010101010;
    LogicCell40 \POWERLED.count_3_LC_4_12_3  (
            .in0(N__18971),
            .in1(_gnd_net_),
            .in2(N__17366),
            .in3(N__24693),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34680),
            .ce(N__21211),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUHGN_3_LC_4_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUHGN_3_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUHGN_3_LC_4_12_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \POWERLED.count_RNIUHGN_3_LC_4_12_4  (
            .in0(N__24692),
            .in1(N__17360),
            .in2(N__17210),
            .in3(N__18970),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIAKSS_0_2_LC_4_13_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIAKSS_0_2_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIAKSS_0_2_LC_4_13_0 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \POWERLED.count_RNIAKSS_0_2_LC_4_13_0  (
            .in0(N__19013),
            .in1(N__17201),
            .in2(N__17483),
            .in3(N__24654),
            .lcout(\POWERLED.count_RNIAKSS_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIAKSS_2_LC_4_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIAKSS_2_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIAKSS_2_LC_4_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNIAKSS_2_LC_4_13_1  (
            .in0(N__24648),
            .in1(N__17478),
            .in2(_gnd_net_),
            .in3(N__19010),
            .lcout(\POWERLED.un1_count_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_4_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_4_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_2_LC_4_13_2  (
            .in0(N__19012),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34685),
            .ce(N__21210),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIAKSS_1_2_LC_4_13_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNIAKSS_1_2_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIAKSS_1_2_LC_4_13_3 .LUT_INIT=16'b0000000000110101;
    LogicCell40 \POWERLED.count_RNIAKSS_1_2_LC_4_13_3  (
            .in0(N__17482),
            .in1(N__19011),
            .in2(N__24691),
            .in3(N__18990),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIT2CB1_4_LC_4_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIT2CB1_4_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIT2CB1_4_LC_4_13_4 .LUT_INIT=16'b0001000011010000;
    LogicCell40 \POWERLED.count_RNIT2CB1_4_LC_4_13_4  (
            .in0(N__17422),
            .in1(N__24653),
            .in2(N__17465),
            .in3(N__18945),
            .lcout(\POWERLED.un79_clk_100khzlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_4_LC_4_13_5 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_4_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_4_LC_4_13_5  (
            .in0(N__18946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34685),
            .ce(N__21210),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIJEFE_4_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIJEFE_4_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIJEFE_4_LC_4_13_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIJEFE_4_LC_4_13_6  (
            .in0(N__17421),
            .in1(N__24649),
            .in2(_gnd_net_),
            .in3(N__18944),
            .lcout(\POWERLED.un1_count_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIJEFE_0_4_LC_4_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIJEFE_0_4_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIJEFE_0_4_LC_4_13_7 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \POWERLED.count_RNIJEFE_0_4_LC_4_13_7  (
            .in0(N__24655),
            .in1(N__17443),
            .in2(N__18950),
            .in3(N__17423),
            .lcout(\POWERLED.count_RNIJEFE_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUGSJ_0_1_LC_4_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUGSJ_0_1_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUGSJ_0_1_LC_4_14_0 .LUT_INIT=16'b0011010100110101;
    LogicCell40 \POWERLED.count_RNIUGSJ_0_1_LC_4_14_0  (
            .in0(N__17504),
            .in1(N__17516),
            .in2(N__24690),
            .in3(N__17399),
            .lcout(\POWERLED.count_RNIUGSJ_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIE5D5_5_LC_4_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIE5D5_5_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIE5D5_5_LC_4_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_RNIE5D5_5_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__24642),
            .in2(_gnd_net_),
            .in3(N__17350),
            .lcout(\POWERLED.count_0_sqmuxa ),
            .ltout(\POWERLED.count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIE5D5_0_LC_4_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIE5D5_0_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIE5D5_0_LC_4_14_2 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \POWERLED.count_RNIE5D5_0_LC_4_14_2  (
            .in0(N__19060),
            .in1(_gnd_net_),
            .in2(N__17333),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNITFSJ_0_LC_4_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNITFSJ_0_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNITFSJ_0_LC_4_14_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNITFSJ_0_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__17495),
            .in2(N__17522),
            .in3(N__24643),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(\POWERLED.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIE5D5_1_LC_4_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIE5D5_1_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIE5D5_1_LC_4_14_4 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \POWERLED.count_RNIE5D5_1_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__19036),
            .in2(N__17519),
            .in3(N__19141),
            .lcout(\POWERLED.count_1_1 ),
            .ltout(\POWERLED.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUGSJ_1_LC_4_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUGSJ_1_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUGSJ_1_LC_4_14_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNIUGSJ_1_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__17503),
            .in2(N__17510),
            .in3(N__24644),
            .lcout(\POWERLED.un1_count_axb_1 ),
            .ltout(\POWERLED.un1_count_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_4_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_4_14_6 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \POWERLED.count_1_LC_4_14_6  (
            .in0(N__19059),
            .in1(_gnd_net_),
            .in2(N__17507),
            .in3(N__19143),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34681),
            .ce(N__21209),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_4_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_4_14_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \POWERLED.count_0_LC_4_14_7  (
            .in0(N__19142),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19058),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34681),
            .ce(N__21209),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_4_15_0 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_4_15_0 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_14_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19196),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34725),
            .ce(N__21215),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIALHT_11_LC_4_15_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIALHT_11_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIALHT_11_LC_4_15_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIALHT_11_LC_4_15_1  (
            .in0(N__17489),
            .in1(N__24688),
            .in2(_gnd_net_),
            .in3(N__19218),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_4_15_2 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_4_15_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_4_15_2 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_11_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19225),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34725),
            .ce(N__21215),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_4_15_4 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_4_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_15_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19087),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34725),
            .ce(N__21215),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGUKT_14_LC_4_15_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGUKT_14_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGUKT_14_LC_4_15_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIGUKT_14_LC_4_15_5  (
            .in0(N__17573),
            .in1(N__24689),
            .in2(_gnd_net_),
            .in3(N__19192),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(\POWERLED.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_4_15_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_4_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_10_LC_4_15_6  (
            .in0(N__19245),
            .in1(N__19272),
            .in2(N__17567),
            .in3(N__20823),
            .lcout(\POWERLED.un79_clk_100khzlto15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI1Q9V_10_LC_4_15_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI1Q9V_10_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI1Q9V_10_LC_4_15_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI1Q9V_10_LC_4_15_7  (
            .in0(N__19418),
            .in1(N__24687),
            .in2(_gnd_net_),
            .in3(N__19434),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNIOF011_LC_4_16_3 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_10_c_RNIOF011_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNIOF011_LC_4_16_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNIOF011_LC_4_16_3  (
            .in0(N__24666),
            .in1(N__19439),
            .in2(N__20485),
            .in3(N__19226),
            .lcout(\POWERLED.g1_i_o4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNII1MT_15_LC_4_16_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNII1MT_15_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNII1MT_15_LC_4_16_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNII1MT_15_LC_4_16_5  (
            .in0(N__24665),
            .in1(_gnd_net_),
            .in2(N__19091),
            .in3(N__17540),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_5_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_2_LC_5_1_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_5_1_0  (
            .in0(N__21490),
            .in1(N__17630),
            .in2(N__21694),
            .in3(N__21008),
            .lcout(\VPP_VDDQ.count_2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34254),
            .ce(N__20040),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_5_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_5_1_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_5_1_1  (
            .in0(N__17629),
            .in1(N__21487),
            .in2(N__21052),
            .in3(N__21636),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_5_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_5_1_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNID4261_2_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(N__17534),
            .in2(N__17528),
            .in3(N__19952),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_2_LC_5_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_5_1_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_2_LC_5_1_3  (
            .in0(N__19295),
            .in1(N__17603),
            .in2(N__17525),
            .in3(N__17747),
            .lcout(\VPP_VDDQ.un9_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_5_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_15_LC_5_1_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_5_1_4  (
            .in0(N__21489),
            .in1(N__21004),
            .in2(N__21693),
            .in3(N__17866),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34254),
            .ce(N__20040),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_5_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_5_1_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_5_1_5  (
            .in0(N__17867),
            .in1(N__21491),
            .in2(N__21054),
            .in3(N__21644),
            .lcout(),
            .ltout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_5_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_5_1_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIL79C1_15_LC_5_1_6  (
            .in0(N__20041),
            .in1(_gnd_net_),
            .in2(N__17645),
            .in3(N__17642),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_5_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_3_LC_5_1_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_5_1_7  (
            .in0(N__19316),
            .in1(N__21488),
            .in2(N__21053),
            .in3(N__21643),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34254),
            .ce(N__20040),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_2_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__19621),
            .in2(N__19604),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_2_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__17636),
            .in2(_gnd_net_),
            .in3(N__17621),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_2_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__19294),
            .in2(_gnd_net_),
            .in3(N__17618),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_2_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__19522),
            .in2(_gnd_net_),
            .in3(N__17606),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_2_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__17599),
            .in2(_gnd_net_),
            .in3(N__17576),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_5_2_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_5_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__19463),
            .in2(_gnd_net_),
            .in3(N__17753),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_2_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__17783),
            .in2(_gnd_net_),
            .in3(N__17750),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_2_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__17746),
            .in2(_gnd_net_),
            .in3(N__17720),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_3_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__17812),
            .in2(_gnd_net_),
            .in3(N__17705),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_3_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__17833),
            .in2(_gnd_net_),
            .in3(N__17684),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_3_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__19871),
            .in2(_gnd_net_),
            .in3(N__17681),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_3_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__17678),
            .in2(_gnd_net_),
            .in3(N__17663),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_3_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(N__17659),
            .in2(_gnd_net_),
            .in3(N__17648),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_3_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__17911),
            .in2(_gnd_net_),
            .in3(N__17888),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_3_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(N__17884),
            .in2(_gnd_net_),
            .in3(N__17870),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_5_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_5_3_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_5_3_7  (
            .in0(N__21551),
            .in1(N__21646),
            .in2(N__21051),
            .in3(N__17851),
            .lcout(\VPP_VDDQ.count_2_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_5_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_5_4_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_1_7_LC_5_4_0  (
            .in0(N__17834),
            .in1(N__17798),
            .in2(N__17822),
            .in3(N__19870),
            .lcout(\VPP_VDDQ.un9_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_5_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_5_4_1 .LUT_INIT=16'b0001000000010011;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_0_7_LC_5_4_1  (
            .in0(N__17792),
            .in1(N__17813),
            .in2(N__20039),
            .in3(N__17762),
            .lcout(\VPP_VDDQ.un9_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_5_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_5_4_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_5_4_2  (
            .in0(N__21705),
            .in1(N__21542),
            .in2(N__21055),
            .in3(N__17774),
            .lcout(\VPP_VDDQ.count_2_1_7 ),
            .ltout(\VPP_VDDQ.count_2_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_5_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_5_4_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_7_LC_5_4_3  (
            .in0(N__20009),
            .in1(_gnd_net_),
            .in2(N__17786),
            .in3(N__17761),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_5_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_7_LC_5_4_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_5_4_4  (
            .in0(N__21706),
            .in1(N__21544),
            .in2(N__21056),
            .in3(N__17773),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34489),
            .ce(N__20047),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_0_LC_5_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_5_4_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_0_LC_5_4_5  (
            .in0(N__21541),
            .in1(N__19599),
            .in2(N__21048),
            .in3(N__21704),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_5_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_5_4_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIT1QU_0_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__18047),
            .in2(N__18053),
            .in3(N__20008),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_0_LC_5_4_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_0_LC_5_4_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_5_4_7  (
            .in0(N__21543),
            .in1(N__21015),
            .in2(N__18050),
            .in3(N__21707),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34489),
            .ce(N__20047),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_5_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_5_5_0  (
            .in0(N__18033),
            .in1(N__17973),
            .in2(N__18004),
            .in3(N__18161),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_5_5_1 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_5_5_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_3_LC_5_5_1  (
            .in0(N__18035),
            .in1(N__29841),
            .in2(_gnd_net_),
            .in3(N__18041),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_5_5_2 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_5_5_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_5_LC_5_5_2  (
            .in0(N__18017),
            .in1(N__17929),
            .in2(_gnd_net_),
            .in3(N__29846),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_5_5_3 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_5_5_3 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \COUNTER.counter_1_LC_5_5_3  (
            .in0(N__18162),
            .in1(_gnd_net_),
            .in2(N__17948),
            .in3(N__29844),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_5_5_4 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_5_5_4 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \COUNTER.counter_2_LC_5_5_4  (
            .in0(N__18011),
            .in1(_gnd_net_),
            .in2(N__18005),
            .in3(N__29845),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_5_5_5 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_5_5_5 .LUT_INIT=16'b0001001000010010;
    LogicCell40 \COUNTER.counter_4_LC_5_5_5  (
            .in0(N__17984),
            .in1(N__29842),
            .in2(N__17978),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_5_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_5_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_5_5_6  (
            .in0(N__17959),
            .in1(N__17943),
            .in2(N__18347),
            .in3(N__17928),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_5_5_7 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_5_5_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_6_LC_5_5_7  (
            .in0(N__18346),
            .in1(N__29843),
            .in2(_gnd_net_),
            .in3(N__18353),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_6_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_5_6_0  (
            .in0(N__18325),
            .in1(N__18313),
            .in2(N__18302),
            .in3(N__18286),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_6_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_5_6_1  (
            .in0(N__18274),
            .in1(N__18262),
            .in2(N__18251),
            .in3(N__18235),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_6_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_6_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_6_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_6_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_5_6_5  (
            .in0(N__18223),
            .in1(N__18211),
            .in2(N__18200),
            .in3(N__18184),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_5_6_7 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_5_6_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \COUNTER.counter_0_LC_5_6_7  (
            .in0(N__29847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18172),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNII6BQ1_0_LC_5_7_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNII6BQ1_0_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNII6BQ1_0_LC_5_7_2 .LUT_INIT=16'b1000100010001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNII6BQ1_0_LC_5_7_2  (
            .in0(N__25319),
            .in1(N__33661),
            .in2(N__18146),
            .in3(N__18125),
            .lcout(\PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_7_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_5_7_3  (
            .in0(N__18103),
            .in1(N__18091),
            .in2(N__18080),
            .in3(N__18064),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_7_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_5_7_7  (
            .in0(N__18487),
            .in1(N__18475),
            .in2(N__18464),
            .in3(N__18448),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__22349),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__18567),
            .in2(N__22256),
            .in3(N__18437),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__18434),
            .in2(N__18572),
            .in3(N__18422),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__18419),
            .in2(N__18608),
            .in3(N__18407),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__18607),
            .in2(N__18404),
            .in3(N__18389),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_8_5  (
            .in0(N__21882),
            .in1(N__18571),
            .in2(N__18386),
            .in3(N__18371),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_8_6  (
            .in0(N__18368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18356),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_8_7  (
            .in0(N__18603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.VCCST_EN_i_1_i_LC_5_9_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.VCCST_EN_i_1_i_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.VCCST_EN_i_1_i_LC_5_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.VCCST_EN_i_1_i_LC_5_9_0  (
            .in0(N__32540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35131),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_12_LC_5_9_1 .C_ON=1'b0;
    defparam \POWERLED.G_12_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_12_LC_5_9_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.G_12_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__24505),
            .in2(_gnd_net_),
            .in3(N__29886),
            .lcout(G_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_LC_5_9_7 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_LC_5_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_0_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__24506),
            .in2(_gnd_net_),
            .in3(N__29887),
            .lcout(suswarn_n),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34701),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20421),
            .lcout(\POWERLED.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22742),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_5_10_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_5_10_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20684),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_10_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22397),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_10_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22427),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22531),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_10_6  (
            .in0(N__18694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__22396),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__18618),
            .in2(N__18653),
            .in3(N__18641),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__20195),
            .in2(N__18623),
            .in3(N__18638),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__20296),
            .in2(N__20186),
            .in3(N__18635),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__20174),
            .in2(N__20300),
            .in3(N__18632),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_11_5  (
            .in0(N__18730),
            .in1(N__18622),
            .in2(N__20165),
            .in3(N__18629),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_11_6  (
            .in0(N__20312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18626),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20295),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__22423),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__18705),
            .in2(N__18884),
            .in3(N__18863),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__18860),
            .in2(N__18710),
            .in3(N__18845),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__18732),
            .in2(N__18842),
            .in3(N__18821),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__18818),
            .in2(N__18737),
            .in3(N__18800),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_12_5  (
            .in0(N__18753),
            .in1(N__18709),
            .in2(N__18797),
            .in3(N__18779),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_12_6  (
            .in0(N__18776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18770),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18731),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_5_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__19057),
            .in2(N__19037),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_5_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_5_13_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_5_13_1  (
            .in0(N__19144),
            .in1(_gnd_net_),
            .in2(N__19022),
            .in3(N__18998),
            .lcout(\POWERLED.count_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18994),
            .in3(N__18962),
            .lcout(\POWERLED.un1_count_cry_2_c_RNICZ0Z419 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2 ),
            .carryout(\POWERLED.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNIEQUS_LC_5_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNIEQUS_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNIEQUS_LC_5_13_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNIEQUS_LC_5_13_3  (
            .in0(N__19145),
            .in1(_gnd_net_),
            .in2(N__18959),
            .in3(N__18932),
            .lcout(\POWERLED.count_1_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3 ),
            .carryout(\POWERLED.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_13_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18929),
            .in3(N__18896),
            .lcout(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNITFHE_LC_5_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNITFHE_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNITFHE_LC_5_13_5 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNITFHE_LC_5_13_5  (
            .in0(N__19146),
            .in1(_gnd_net_),
            .in2(N__19410),
            .in3(N__18893),
            .lcout(\POWERLED.count_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_5_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_5_13_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_5_13_6  (
            .in0(N__19160),
            .in1(_gnd_net_),
            .in2(N__20754),
            .in3(N__18890),
            .lcout(\POWERLED.count_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_5_13_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_5_13_7 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_5_13_7  (
            .in0(N__19147),
            .in1(_gnd_net_),
            .in2(N__20518),
            .in3(N__18887),
            .lcout(\POWERLED.count_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_5_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_5_14_0 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_5_14_0  (
            .in0(N__19172),
            .in1(_gnd_net_),
            .in2(N__20483),
            .in3(N__19283),
            .lcout(\POWERLED.count_1_9 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_5_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_5_14_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_5_14_1  (
            .in0(N__19161),
            .in1(_gnd_net_),
            .in2(N__19276),
            .in3(N__19253),
            .lcout(\POWERLED.count_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_5_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_5_14_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_5_14_2  (
            .in0(N__19173),
            .in1(_gnd_net_),
            .in2(N__19249),
            .in3(N__19205),
            .lcout(\POWERLED.count_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_5_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_5_14_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_5_14_3  (
            .in0(N__19162),
            .in1(_gnd_net_),
            .in2(N__19073),
            .in3(N__19202),
            .lcout(\POWERLED.count_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_5_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_5_14_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_5_14_4  (
            .in0(N__19174),
            .in1(_gnd_net_),
            .in2(N__20578),
            .in3(N__19199),
            .lcout(\POWERLED.count_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNICO0D_LC_5_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNICO0D_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNICO0D_LC_5_14_5 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNICO0D_LC_5_14_5  (
            .in0(N__19163),
            .in1(_gnd_net_),
            .in2(N__20802),
            .in3(N__19184),
            .lcout(\POWERLED.count_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_5_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_5_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_5_14_6  (
            .in0(N__19175),
            .in1(N__20841),
            .in2(_gnd_net_),
            .in3(N__19094),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICOIT_12_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNICOIT_12_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICOIT_12_LC_5_14_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNICOIT_12_LC_5_14_7  (
            .in0(N__20559),
            .in1(N__24664),
            .in2(_gnd_net_),
            .in3(N__20534),
            .lcout(\POWERLED.un1_count_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIO94T_9_LC_5_15_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIO94T_9_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIO94T_9_LC_5_15_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIO94T_9_LC_5_15_1  (
            .in0(N__24663),
            .in1(_gnd_net_),
            .in2(N__19457),
            .in3(N__19445),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_5_15_2 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_5_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_9_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19456),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34686),
            .ce(N__21208),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_5_15_3 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_5_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_10_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19435),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34686),
            .ce(N__21208),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNII01T_6_LC_5_15_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNII01T_6_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNII01T_6_LC_5_15_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNII01T_6_LC_5_15_4  (
            .in0(N__19358),
            .in1(N__24661),
            .in2(_gnd_net_),
            .in3(N__19377),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_5_15_5 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_5_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_6_LC_5_15_5  (
            .in0(N__19378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34686),
            .ce(N__21208),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIM63T_8_LC_5_15_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIM63T_8_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIM63T_8_LC_5_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNIM63T_8_LC_5_15_7  (
            .in0(N__24662),
            .in1(N__19325),
            .in2(_gnd_net_),
            .in3(N__19347),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_5_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_5_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_8_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19348),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34724),
            .ce(N__21213),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_6_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_6_1_0 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_6_1_0  (
            .in0(N__21371),
            .in1(N__21426),
            .in2(N__21349),
            .in3(N__21237),
            .lcout(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_6_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_6_1_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_6_1_2  (
            .in0(N__21480),
            .in1(N__19315),
            .in2(N__20981),
            .in3(N__21645),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_6_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_6_1_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIF7361_3_LC_6_1_3  (
            .in0(N__19304),
            .in1(_gnd_net_),
            .in2(N__19298),
            .in3(N__19953),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_1_5 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_1_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_6_1_5  (
            .in0(N__19543),
            .in1(N__21344),
            .in2(N__19820),
            .in3(N__19840),
            .lcout(\VPP_VDDQ.delayed_vddq_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34062),
            .ce(),
            .sr(N__19859));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI6JOT1_LC_6_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI6JOT1_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI6JOT1_LC_6_1_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNI6JOT1_LC_6_1_6  (
            .in0(N__19841),
            .in1(N__19819),
            .in2(N__21350),
            .in3(N__19544),
            .lcout(),
            .ltout(VPP_VDDQ_delayed_vddq_ok_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_PWRGD_LC_6_1_7 .C_ON=1'b0;
    defparam \POWERLED.VCCST_PWRGD_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_PWRGD_LC_6_1_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.VCCST_PWRGD_LC_6_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19535),
            .in3(N__25114),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_6_LC_6_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_6_LC_6_2_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_6_2_1  (
            .in0(N__21428),
            .in1(N__19492),
            .in2(N__20957),
            .in3(N__21648),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34264),
            .ce(N__20042),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_6_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_6_2_2 .LUT_INIT=16'b0000000000110101;
    LogicCell40 \VPP_VDDQ.count_2_RNI38QU_0_6_LC_6_2_2  (
            .in0(N__19472),
            .in1(N__19481),
            .in2(N__20048),
            .in3(N__19526),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_6_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_6_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIOUR33_1_LC_6_2_3  (
            .in0(N__19574),
            .in1(N__19511),
            .in2(N__19505),
            .in3(N__19502),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(\VPP_VDDQ.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_6_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_6_2_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_6_2_4  (
            .in0(N__19493),
            .in1(N__20895),
            .in2(N__19484),
            .in3(N__21427),
            .lcout(\VPP_VDDQ.count_2_1_6 ),
            .ltout(\VPP_VDDQ.count_2_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_6_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_6_2_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI38QU_6_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(N__19934),
            .in2(N__19475),
            .in3(N__19471),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_6_2_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_6_2_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_6_2_6  (
            .in0(N__19762),
            .in1(N__19739),
            .in2(N__19670),
            .in3(N__19720),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_SUSn_RNIN4K9_LC_6_2_7.C_ON=1'b0;
    defparam SLP_SUSn_RNIN4K9_LC_6_2_7.SEQ_MODE=4'b0000;
    defparam SLP_SUSn_RNIN4K9_LC_6_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 SLP_SUSn_RNIN4K9_LC_6_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19669),
            .lcout(v33a_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_6_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_6_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__19595),
            .in2(_gnd_net_),
            .in3(N__19622),
            .lcout(\VPP_VDDQ.count_2_RNIZ0Z_1 ),
            .ltout(\VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_6_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_6_3_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_1_LC_6_3_1  (
            .in0(N__21518),
            .in1(N__20986),
            .in2(N__19628),
            .in3(N__21632),
            .lcout(\VPP_VDDQ.count_2_1_1 ),
            .ltout(\VPP_VDDQ.count_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_6_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_6_3_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIU2QU_1_LC_6_3_2  (
            .in0(N__19960),
            .in1(_gnd_net_),
            .in2(N__19625),
            .in3(N__19561),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_6_3_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_6_3_3 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_6_3_3  (
            .in0(N__19562),
            .in1(N__19610),
            .in2(N__19603),
            .in3(N__20024),
            .lcout(\VPP_VDDQ.un9_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_6_3_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_1_LC_6_3_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_6_3_4  (
            .in0(N__21633),
            .in1(N__21522),
            .in2(N__21049),
            .in3(N__19568),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34198),
            .ce(N__20023),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_11_LC_6_3_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_11_LC_6_3_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_6_3_5  (
            .in0(N__19552),
            .in1(N__20987),
            .in2(N__21546),
            .in3(N__21634),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34198),
            .ce(N__20023),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_6_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_6_3_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_6_3_6  (
            .in0(N__21635),
            .in1(N__19553),
            .in2(N__21050),
            .in3(N__21523),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_6_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_6_3_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIDR4C1_11_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(N__19959),
            .in2(N__19880),
            .in3(N__19877),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_6_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_6_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNO_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19834),
            .lcout(\VPP_VDDQ.N_60_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_6_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_6_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20982),
            .lcout(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_6_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_6_4_4 .LUT_INIT=16'b1011101011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_6_4_4  (
            .in0(N__21516),
            .in1(N__21306),
            .in2(N__19844),
            .in3(N__24630),
            .lcout(\VPP_VDDQ.N_60 ),
            .ltout(\VPP_VDDQ.N_60_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_6_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_6_4_5 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNINI731_0_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(N__21517),
            .in2(N__19823),
            .in3(N__21238),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_6_5_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_6_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19805),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_6_5_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_6_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19796),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_6_5_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_6_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19787),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_6_5_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_6_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19778),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_6_5_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_6_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20108),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_6_5_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_6_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20099),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_6_5_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_6_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20087),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_6_5_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_6_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20075),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(COUNTER_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_6_0.C_ON=1'b0;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20060),
            .lcout(COUNTER_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_6_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25852),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_6_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_6_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__30417),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__20148),
            .in2(N__20057),
            .in3(N__22121),
            .lcout(G_2161),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__22037),
            .in2(N__20153),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__22122),
            .in2(N__22019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__21992),
            .in2(N__22129),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__20152),
            .in2(N__22196),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_7_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_7_6  (
            .in0(N__22154),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20138),
            .lcout(\POWERLED.mult1_un166_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_7_7  (
            .in0(N__22236),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_6_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_6_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_6_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23822),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34426),
            .ce(N__34002),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_52_and_i_o3_0_a2_0_LC_6_9_0 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_52_and_i_o3_0_a2_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_52_and_i_o3_0_a2_0_LC_6_9_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.un1_clk_100khz_52_and_i_o3_0_a2_0_LC_6_9_0  (
            .in0(N__35443),
            .in1(N__32541),
            .in2(_gnd_net_),
            .in3(N__35097),
            .lcout(\POWERLED.N_600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_6_9_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_6_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21883),
            .lcout(\POWERLED.mult1_un145_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5QAN_0_LC_6_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5QAN_0_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5QAN_0_LC_6_9_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \POWERLED.func_state_RNI5QAN_0_LC_6_9_2  (
            .in0(N__35442),
            .in1(N__32408),
            .in2(_gnd_net_),
            .in3(N__29314),
            .lcout(\POWERLED.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22621),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_9_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22700),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20422),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22718),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__22738),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__20201),
            .in2(N__20329),
            .in3(N__20189),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__20325),
            .in2(N__20255),
            .in3(N__20177),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__20417),
            .in2(N__20243),
            .in3(N__20168),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__20231),
            .in2(N__20423),
            .in3(N__20156),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_10_5  (
            .in0(N__20294),
            .in1(N__20222),
            .in2(N__20330),
            .in3(N__20306),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20438),
            .in3(N__20303),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(\POWERLED.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20279),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__22714),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__20264),
            .in2(N__20650),
            .in3(N__20246),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__20646),
            .in2(N__20384),
            .in3(N__20234),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__20372),
            .in2(N__20680),
            .in3(N__20225),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__20676),
            .in2(N__20363),
            .in3(N__20216),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5  (
            .in0(N__20416),
            .in1(N__20351),
            .in2(N__20651),
            .in3(N__20429),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20342),
            .in3(N__20426),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22666),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(N__22696),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(N__20390),
            .in2(N__22801),
            .in3(N__20375),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__22797),
            .in2(N__21146),
            .in3(N__20366),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(N__22900),
            .in2(N__21131),
            .in3(N__20354),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__21116),
            .in2(N__22904),
            .in3(N__20345),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_12_5  (
            .in0(N__20672),
            .in1(N__21104),
            .in2(N__22802),
            .in3(N__20333),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(N__21092),
            .in2(_gnd_net_),
            .in3(N__20687),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(\POWERLED.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20654),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICOIT_0_12_LC_6_13_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNICOIT_0_12_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICOIT_0_12_LC_6_13_0 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \POWERLED.count_RNICOIT_0_12_LC_6_13_0  (
            .in0(N__20561),
            .in1(N__20633),
            .in2(N__20543),
            .in3(N__24641),
            .lcout(\POWERLED.count_RNICOIT_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_6_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_6_13_2 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_12_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20542),
            .in3(_gnd_net_),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34557),
            .ce(N__21207),
            .sr(_gnd_net_));
    defparam \POWERLED.count_13_LC_6_13_3 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_6_13_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_13_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20594),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34557),
            .ce(N__21207),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIERJT_13_LC_6_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIERJT_13_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIERJT_13_LC_6_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIERJT_13_LC_6_13_4  (
            .in0(N__20600),
            .in1(N__24639),
            .in2(_gnd_net_),
            .in3(N__20590),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(\POWERLED.countZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICOIT_1_12_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNICOIT_1_12_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICOIT_1_12_LC_6_13_5 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \POWERLED.count_RNICOIT_1_12_LC_6_13_5  (
            .in0(N__24640),
            .in1(N__20560),
            .in2(N__20546),
            .in3(N__20535),
            .lcout(\POWERLED.un79_clk_100khzlto15_3 ),
            .ltout(\POWERLED.un79_clk_100khzlto15_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICOIT_5_12_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNICOIT_5_12_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICOIT_5_12_LC_6_13_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.count_RNICOIT_5_12_LC_6_13_6  (
            .in0(N__20517),
            .in1(N__20484),
            .in2(N__20450),
            .in3(N__20747),
            .lcout(\POWERLED.un79_clk_100khzlto15_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICOIT_4_12_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNICOIT_4_12_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICOIT_4_12_LC_6_13_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.count_RNICOIT_4_12_LC_6_13_7  (
            .in0(N__20849),
            .in1(N__20842),
            .in2(N__20755),
            .in3(N__20807),
            .lcout(\POWERLED.g1_i_o4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIK32T_7_LC_6_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIK32T_7_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIK32T_7_LC_6_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIK32T_7_LC_6_14_0  (
            .in0(N__20717),
            .in1(N__24631),
            .in2(_gnd_net_),
            .in3(N__20725),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_6_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_6_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_7_LC_6_14_1  (
            .in0(N__20726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34553),
            .ce(N__21212),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI12AS_8_LC_6_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI12AS_8_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI12AS_8_LC_6_14_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \POWERLED.dutycycle_RNI12AS_8_LC_6_14_3  (
            .in0(N__30291),
            .in1(N__32483),
            .in2(_gnd_net_),
            .in3(N__32960),
            .lcout(\POWERLED.un1_clk_100khz_32_and_i_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6SKJ1_0_LC_6_14_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6SKJ1_0_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6SKJ1_0_LC_6_14_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI6SKJ1_0_LC_6_14_4  (
            .in0(N__32484),
            .in1(N__20708),
            .in2(_gnd_net_),
            .in3(N__30290),
            .lcout(\POWERLED.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI4MHI4_4_LC_6_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI4MHI4_4_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI4MHI4_4_LC_6_14_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI4MHI4_4_LC_6_14_5  (
            .in0(N__23870),
            .in1(N__33986),
            .in2(_gnd_net_),
            .in3(N__23846),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINE7B4_0_10_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINE7B4_0_10_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINE7B4_0_10_LC_6_14_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \POWERLED.count_clk_RNINE7B4_0_10_LC_6_14_6  (
            .in0(N__33988),
            .in1(_gnd_net_),
            .in2(N__26651),
            .in3(N__26696),
            .lcout(\POWERLED.un1_count_clk_2_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8SJI4_6_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8SJI4_6_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8SJI4_6_LC_6_14_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI8SJI4_6_LC_6_14_7  (
            .in0(N__20699),
            .in1(N__33987),
            .in2(_gnd_net_),
            .in3(N__23821),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_6_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_6_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22670),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_6_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_6_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22817),
            .in3(N__21134),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_6_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_6_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__22844),
            .in2(N__22826),
            .in3(N__21119),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_6_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_6_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__23147),
            .in2(N__22976),
            .in3(N__21107),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_6_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_6_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__23148),
            .in2(N__22955),
            .in3(N__21095),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_6_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_6_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_6_15_5  (
            .in0(N__22898),
            .in1(N__22934),
            .in2(N__21077),
            .in3(N__21083),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_6_15_6 .C_ON=1'b0;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_6_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21080),
            .lcout(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_15_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_15_7  (
            .in0(N__22932),
            .in1(N__22933),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_7_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_7_1_0 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_7_1_0  (
            .in0(N__21274),
            .in1(N__21372),
            .in2(N__21348),
            .in3(N__21425),
            .lcout(\VPP_VDDQ.N_53 ),
            .ltout(\VPP_VDDQ.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_7_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_7_1_1 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_7_1_1  (
            .in0(N__24695),
            .in1(_gnd_net_),
            .in2(N__21068),
            .in3(N__21254),
            .lcout(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_7_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_7_1_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_7_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21722),
            .in3(N__21647),
            .lcout(\VPP_VDDQ.N_664 ),
            .ltout(\VPP_VDDQ.N_664_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_7_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_7_1_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_7_1_3  (
            .in0(N__21374),
            .in1(N__21481),
            .in2(N__21557),
            .in3(N__21337),
            .lcout(),
            .ltout(\VPP_VDDQ.m4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_7_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_7_1_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_7_1_4  (
            .in0(_gnd_net_),
            .in1(N__21266),
            .in2(N__21554),
            .in3(N__24694),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_0_LC_7_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_7_1_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_7_1_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_7_1_5  (
            .in0(N__21373),
            .in1(N__21336),
            .in2(N__21278),
            .in3(N__21275),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34061),
            .ce(N__21199),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_1_LC_7_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_7_1_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_7_1_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_7_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21260),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34061),
            .ce(N__21199),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_m0_0_0_a2_2_0_LC_7_2_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_m0_0_0_a2_2_0_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_1_m0_0_0_a2_2_0_LC_7_2_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.func_state_1_m0_0_0_a2_2_0_LC_7_2_0  (
            .in0(N__35474),
            .in1(N__32656),
            .in2(_gnd_net_),
            .in3(N__24675),
            .lcout(\POWERLED.N_627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI4MLK1_1_LC_7_2_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI4MLK1_1_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI4MLK1_1_LC_7_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNI4MLK1_1_LC_7_2_2  (
            .in0(N__23041),
            .in1(N__23257),
            .in2(N__23078),
            .in3(N__23059),
            .lcout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIVSS4_11_LC_7_2_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIVSS4_11_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIVSS4_11_LC_7_2_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIVSS4_11_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(N__23212),
            .in2(_gnd_net_),
            .in3(N__23227),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI5BM11_10_LC_7_2_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI5BM11_10_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI5BM11_10_LC_7_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNI5BM11_10_LC_7_2_4  (
            .in0(N__23242),
            .in1(N__23272),
            .in2(N__21149),
            .in3(N__23023),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIST215_10_LC_7_2_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIST215_10_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIST215_10_LC_7_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIST215_10_LC_7_2_5  (
            .in0(N__24338),
            .in1(N__21833),
            .in2(N__21827),
            .in3(N__21824),
            .lcout(\RSMRST_PWRGD.N_662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_7_2_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_7_2_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_7_2_7  (
            .in0(N__23182),
            .in1(N__23197),
            .in2(N__23093),
            .in3(N__23287),
            .lcout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_7_3_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_7_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_7_3_0  (
            .in0(_gnd_net_),
            .in1(N__30140),
            .in2(_gnd_net_),
            .in3(N__23422),
            .lcout(\POWERLED.N_613 ),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_3_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__21861),
            .in2(N__22073),
            .in3(N__21818),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_3_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__21815),
            .in2(N__21866),
            .in3(N__21800),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_3_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_3_3  (
            .in0(_gnd_net_),
            .in1(N__21895),
            .in2(N__21797),
            .in3(N__21779),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_3_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_3_4  (
            .in0(_gnd_net_),
            .in1(N__21776),
            .in2(N__21899),
            .in3(N__21761),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_3_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_3_5  (
            .in0(N__22212),
            .in1(N__21865),
            .in2(N__21758),
            .in3(N__21740),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_3_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_3_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_3_6  (
            .in0(_gnd_net_),
            .in1(N__21737),
            .in2(_gnd_net_),
            .in3(N__21902),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_7_3_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_7_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_7_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21894),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_7_4_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_7_4_0 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_7_4_0 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \POWERLED.dutycycle_2_LC_7_4_0  (
            .in0(N__21851),
            .in1(N__27551),
            .in2(N__23342),
            .in3(N__33589),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34293),
            .ce(),
            .sr(N__31539));
    defparam \POWERLED.dutycycle_RNIA8C49_2_LC_7_4_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIA8C49_2_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIA8C49_2_LC_7_4_1 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_RNIA8C49_2_LC_7_4_1  (
            .in0(N__27550),
            .in1(N__21850),
            .in2(N__33643),
            .in3(N__23338),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(\POWERLED.dutycycleZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_2_LC_7_4_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_7_4_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \POWERLED.dutycycle_RNI_1_2_LC_7_4_2  (
            .in0(_gnd_net_),
            .in1(N__33122),
            .in2(N__21842),
            .in3(N__32270),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_LC_7_4_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_LC_7_4_3 .LUT_INIT=16'b1100001110000111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_LC_7_4_3  (
            .in0(N__31407),
            .in1(N__25835),
            .in2(N__21839),
            .in3(N__31025),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_2_LC_7_4_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_7_4_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_2_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21836),
            .in3(N__30150),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_7_4_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_7_4_5 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_7_4_5  (
            .in0(N__31408),
            .in1(N__25836),
            .in2(N__30175),
            .in3(N__31026),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_1_LC_7_4_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_7_4_6 .LUT_INIT=16'b0000111101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_1_LC_7_4_6  (
            .in0(N__31024),
            .in1(_gnd_net_),
            .in2(N__25867),
            .in3(N__31406),
            .lcout(\POWERLED.un1_dutycycle_53_axb_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIER938_0_LC_7_5_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIER938_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIER938_0_LC_7_5_0 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \POWERLED.dutycycle_RNIER938_0_LC_7_5_0  (
            .in0(N__33600),
            .in1(N__21958),
            .in2(N__21971),
            .in3(N__23368),
            .lcout(\POWERLED.dutycycle ),
            .ltout(\POWERLED.dutycycle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_0_LC_7_5_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_0_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_0_LC_7_5_1 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_0_LC_7_5_1  (
            .in0(N__27339),
            .in1(N__33358),
            .in2(N__21974),
            .in3(N__27415),
            .lcout(\POWERLED.dutycycle_1_0_0 ),
            .ltout(\POWERLED.dutycycle_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_7_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_7_5_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_7_5_2 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \POWERLED.dutycycle_0_LC_7_5_2  (
            .in0(N__33602),
            .in1(N__23369),
            .in2(N__21962),
            .in3(N__21959),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34245),
            .ce(),
            .sr(N__31538));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_5_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_5_3 .LUT_INIT=16'b1110101011111011;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_5_3  (
            .in0(N__27340),
            .in1(N__33359),
            .in2(N__27421),
            .in3(N__25778),
            .lcout(\POWERLED.dutycycle_1_0_1 ),
            .ltout(\POWERLED.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNII6848_1_LC_7_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNII6848_1_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNII6848_1_LC_7_5_4 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \POWERLED.dutycycle_RNII6848_1_LC_7_5_4  (
            .in0(N__33601),
            .in1(N__21928),
            .in2(N__21950),
            .in3(N__21944),
            .lcout(dutycycle_RNII6848_0_1),
            .ltout(dutycycle_RNII6848_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITL8S5_1_LC_7_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITL8S5_1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITL8S5_1_LC_7_5_5 .LUT_INIT=16'b0101010011111111;
    LogicCell40 \POWERLED.dutycycle_RNITL8S5_1_LC_7_5_5  (
            .in0(N__23359),
            .in1(N__30712),
            .in2(N__21947),
            .in3(N__33739),
            .lcout(\POWERLED.dutycycle_eena_0 ),
            .ltout(\POWERLED.dutycycle_eena_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_7_5_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_7_5_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_7_5_6 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_1_LC_7_5_6  (
            .in0(N__21938),
            .in1(N__21929),
            .in2(N__21932),
            .in3(N__33603),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34245),
            .ce(),
            .sr(N__31538));
    defparam \POWERLED.func_state_RNI4R67A_1_LC_7_6_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4R67A_1_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4R67A_1_LC_7_6_0 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \POWERLED.func_state_RNI4R67A_1_LC_7_6_0  (
            .in0(N__22082),
            .in1(N__24413),
            .in2(N__21920),
            .in3(N__29247),
            .lcout(\POWERLED.N_13_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_2_LC_7_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_2_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_2_LC_7_6_1 .LUT_INIT=16'b0001110111011101;
    LogicCell40 \POWERLED.dutycycle_RNI_4_2_LC_7_6_1  (
            .in0(N__31017),
            .in1(N__22289),
            .in2(N__30204),
            .in3(N__30630),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_7_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_7_6_2 .LUT_INIT=16'b1010111010100100;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_2_LC_7_6_2  (
            .in0(N__22288),
            .in1(N__27341),
            .in2(N__21905),
            .in3(N__29559),
            .lcout(POWERLED_un1_dutycycle_172_m1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_0_LC_7_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_7_6_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_0_LC_7_6_3  (
            .in0(N__25848),
            .in1(N__23423),
            .in2(N__30400),
            .in3(N__33108),
            .lcout(),
            .ltout(\POWERLED.N_672_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_5_LC_7_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_7_6_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_5_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__35576),
            .in2(N__22058),
            .in3(N__31016),
            .lcout(dutycycle_RNI_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_1_LC_7_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_7_6_6 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_1_LC_7_6_6  (
            .in0(N__30629),
            .in1(N__22055),
            .in2(N__29572),
            .in3(N__23480),
            .lcout(),
            .ltout(dutycycle_RNI_3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNINCRN3_LC_7_6_7 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNINCRN3_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNINCRN3_LC_7_6_7 .LUT_INIT=16'b0000101100000000;
    LogicCell40 \COUNTER.tmp_0_fast_RNINCRN3_LC_7_6_7  (
            .in0(N__22054),
            .in1(N__22046),
            .in2(N__22040),
            .in3(N__25711),
            .lcout(G_11_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_7_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_7_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_1_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__25872),
            .in2(_gnd_net_),
            .in3(N__35642),
            .lcout(N_50),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__22179),
            .in2(N__22100),
            .in3(N__22031),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__22028),
            .in2(N__22184),
            .in3(N__22010),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__22232),
            .in2(N__22007),
            .in3(N__21986),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__21983),
            .in2(N__22240),
            .in3(N__22187),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_7_5  (
            .in0(N__22120),
            .in1(N__22183),
            .in2(N__22169),
            .in3(N__22148),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_7_6  (
            .in0(N__22145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22136),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30194),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_141_LC_7_8_1 .C_ON=1'b0;
    defparam \POWERLED.G_141_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_141_LC_7_8_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.G_141_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29945),
            .in3(N__29848),
            .lcout(G_141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_7_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_7_8_2 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_7_8_2  (
            .in0(N__22091),
            .in1(N__33124),
            .in2(N__22552),
            .in3(N__32272),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIT53D6_1_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIT53D6_1_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIT53D6_1_LC_7_8_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \POWERLED.func_state_RNIT53D6_1_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__22262),
            .in2(_gnd_net_),
            .in3(N__29849),
            .lcout(\POWERLED.g0_7_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_0_LC_7_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_7_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_0_LC_7_8_4  (
            .in0(N__30395),
            .in1(N__31409),
            .in2(_gnd_net_),
            .in3(N__25868),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_8_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22345),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_rep1_LC_7_8_6 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_rep1_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_rep1_LC_7_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \COUNTER.tmp_0_rep1_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29872),
            .in3(N__29928),
            .lcout(SUSWARN_N_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34425),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_0_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_7_8_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_0_LC_7_8_7  (
            .in0(N__25869),
            .in1(N__22274),
            .in2(N__35575),
            .in3(N__30396),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_7_9_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_7_9_0  (
            .in0(N__32959),
            .in1(N__23513),
            .in2(N__25907),
            .in3(N__28508),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_0_a2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_9_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_14_LC_7_9_1  (
            .in0(N__34969),
            .in1(N__22273),
            .in2(N__22277),
            .in3(N__22355),
            .lcout(\POWERLED.N_612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_7_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_7_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_7_9_2  (
            .in0(N__32274),
            .in1(N__31400),
            .in2(_gnd_net_),
            .in3(N__32846),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_LC_7_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_7_9_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_7_9_3  (
            .in0(N__26228),
            .in1(N__23609),
            .in2(N__26108),
            .in3(N__23579),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_3_LC_7_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_3_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_3_LC_7_9_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.dutycycle_RNI_13_3_LC_7_9_5  (
            .in0(N__32847),
            .in1(N__31386),
            .in2(_gnd_net_),
            .in3(N__32275),
            .lcout(\POWERLED.N_604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1O2V5_1_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1O2V5_1_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1O2V5_1_LC_7_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI1O2V5_1_LC_7_9_6  (
            .in0(N__30882),
            .in1(N__29939),
            .in2(N__32590),
            .in3(N__26918),
            .lcout(\POWERLED.func_state_RNI1O2V5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22309),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_8_LC_7_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_7_10_0 .LUT_INIT=16'b0000010101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_8_LC_7_10_0  (
            .in0(N__31410),
            .in1(_gnd_net_),
            .in2(N__31252),
            .in3(N__31820),
            .lcout(),
            .ltout(\POWERLED.N_9_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_7_10_1 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_7_10_1  (
            .in0(N__33144),
            .in1(N__31224),
            .in2(N__22376),
            .in3(N__32831),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_7_10_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_7_10_2  (
            .in0(N__31225),
            .in1(N__28529),
            .in2(N__22373),
            .in3(N__31821),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI14KO1_8_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI14KO1_8_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI14KO1_8_LC_7_10_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \POWERLED.dutycycle_RNI14KO1_8_LC_7_10_3  (
            .in0(N__27661),
            .in1(N__22370),
            .in2(N__31254),
            .in3(N__31892),
            .lcout(\POWERLED.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI02AS_1_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI02AS_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI02AS_1_LC_7_10_4 .LUT_INIT=16'b1100111111111111;
    LogicCell40 \POWERLED.func_state_RNI02AS_1_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__27660),
            .in2(N__27814),
            .in3(N__32529),
            .lcout(\POWERLED.N_421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_6_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_7_10_5 .LUT_INIT=16'b1101110011000100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_6_LC_7_10_5  (
            .in0(N__23552),
            .in1(N__33123),
            .in2(N__31826),
            .in3(N__32830),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_6 ),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_7_10_6 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_7_10_6  (
            .in0(N__32832),
            .in1(N__31230),
            .in2(N__22358),
            .in3(N__28202),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_10_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_7_10_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_10_LC_7_10_7  (
            .in0(N__28310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33173),
            .lcout(\POWERLED.un2_count_clk_17_0_0_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_11_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_0_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__32276),
            .in2(N__30416),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_53_axb_0 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__30394),
            .in2(N__22328),
            .in3(N__22292),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__22637),
            .in2(N__30195),
            .in3(N__22604),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__22601),
            .in2(N__30206),
            .in3(N__22568),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__22565),
            .in2(N__22553),
            .in3(N__22511),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__31027),
            .in2(N__30926),
            .in3(N__22490),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__31028),
            .in2(N__23435),
            .in3(N__22466),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__28309),
            .in2(N__23681),
            .in3(N__22442),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__28198),
            .in2(N__22439),
            .in3(N__22409),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__22406),
            .in2(N__28525),
            .in3(N__22379),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__26242),
            .in2(N__26171),
            .in3(N__22721),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__34934),
            .in2(N__26087),
            .in3(N__22703),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__31107),
            .in2(N__23693),
            .in3(N__22685),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__26237),
            .in2(N__22682),
            .in3(N__22652),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_12_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__34936),
            .in2(N__23666),
            .in3(N__22649),
            .lcout(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_12_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__31085),
            .in2(N__23738),
            .in3(N__22646),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__31108),
            .in2(N__22784),
            .in3(N__22643),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22640),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23002),
            .lcout(\POWERLED.un1_dutycycle_53_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22899),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_7_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_7_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__34935),
            .in2(_gnd_net_),
            .in3(N__23750),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIC2MI4_8_LC_7_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIC2MI4_8_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIC2MI4_8_LC_7_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNIC2MI4_8_LC_7_14_0  (
            .in0(N__22775),
            .in1(N__33955),
            .in2(_gnd_net_),
            .in3(N__23944),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_7_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_7_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_8_LC_7_14_1  (
            .in0(N__23945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34552),
            .ce(N__33933),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDTBQ11_7_LC_7_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDTBQ11_7_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDTBQ11_7_LC_7_14_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIDTBQ11_7_LC_7_14_3  (
            .in0(N__28589),
            .in1(N__29461),
            .in2(_gnd_net_),
            .in3(N__28613),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIF0DQ11_8_LC_7_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIF0DQ11_8_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIF0DQ11_8_LC_7_14_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \POWERLED.count_off_RNIF0DQ11_8_LC_7_14_4  (
            .in0(N__29462),
            .in1(_gnd_net_),
            .in2(N__28550),
            .in3(N__28574),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_14_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_14_5 .LUT_INIT=16'b1100110011000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__22768),
            .in2(N__22760),
            .in3(N__22873),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_14_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_14_6  (
            .in0(N__22769),
            .in1(_gnd_net_),
            .in2(N__22877),
            .in3(N__22758),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_14_7 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22759),
            .in3(N__22872),
            .lcout(\POWERLED.mult1_un47_sum_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23006),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22853),
            .in3(N__22988),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_15_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22985),
            .in3(N__22967),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__23163),
            .in2(N__22964),
            .in3(N__22946),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__22943),
            .in2(N__23168),
            .in3(N__22919),
            .lcout(\POWERLED.mult1_un47_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_15_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_15_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22916),
            .in3(N__22907),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22871),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7  (
            .in0(N__22842),
            .in1(N__22843),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_7_16_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_10_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26691),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34655),
            .ce(N__33992),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_8_1_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_8_1_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_8_1_0  (
            .in0(N__24138),
            .in1(N__23092),
            .in2(N__24323),
            .in3(N__24322),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_1_LC_8_1_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_8_1_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_8_1_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_8_1_1  (
            .in0(N__24134),
            .in1(N__23077),
            .in2(_gnd_net_),
            .in3(N__23063),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_2_LC_8_1_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_8_1_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_8_1_2  (
            .in0(N__24139),
            .in1(N__23060),
            .in2(_gnd_net_),
            .in3(N__23048),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_3_LC_8_1_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_8_1_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_8_1_3  (
            .in0(N__24135),
            .in1(N__24350),
            .in2(_gnd_net_),
            .in3(N__23045),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_4_LC_8_1_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_8_1_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_8_1_4  (
            .in0(N__24140),
            .in1(N__23042),
            .in2(_gnd_net_),
            .in3(N__23030),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_5_LC_8_1_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_8_1_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_8_1_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_8_1_5  (
            .in0(N__24136),
            .in1(N__24377),
            .in2(_gnd_net_),
            .in3(N__23027),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_6_LC_8_1_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_8_1_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_8_1_6  (
            .in0(N__24141),
            .in1(N__23024),
            .in2(_gnd_net_),
            .in3(N__23012),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_7_LC_8_1_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_8_1_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_8_1_7  (
            .in0(N__24137),
            .in1(N__24364),
            .in2(_gnd_net_),
            .in3(N__23009),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__34063),
            .ce(),
            .sr(N__24186));
    defparam \RSMRST_PWRGD.count_8_LC_8_2_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_8_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_8_2_0  (
            .in0(N__24148),
            .in1(N__23273),
            .in2(_gnd_net_),
            .in3(N__23261),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.count_9_LC_8_2_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_8_2_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_8_2_1  (
            .in0(N__24144),
            .in1(N__23258),
            .in2(_gnd_net_),
            .in3(N__23246),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.count_10_LC_8_2_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_8_2_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_8_2_2  (
            .in0(N__24145),
            .in1(N__23243),
            .in2(_gnd_net_),
            .in3(N__23231),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.count_11_LC_8_2_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_8_2_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_8_2_3  (
            .in0(N__24142),
            .in1(N__23228),
            .in2(_gnd_net_),
            .in3(N__23216),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.count_12_LC_8_2_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_8_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_8_2_4  (
            .in0(N__24146),
            .in1(N__23213),
            .in2(_gnd_net_),
            .in3(N__23201),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.count_13_LC_8_2_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_8_2_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_8_2_5  (
            .in0(N__24143),
            .in1(N__23198),
            .in2(_gnd_net_),
            .in3(N__23186),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.count_14_LC_8_2_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_8_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_8_2_6  (
            .in0(N__24147),
            .in1(N__23183),
            .in2(_gnd_net_),
            .in3(N__23171),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__34286),
            .ce(),
            .sr(N__24193));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__23134),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_3_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_3_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__23288),
            .in2(_gnd_net_),
            .in3(N__23291),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34333),
            .ce(N__23957),
            .sr(N__24194));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIHIN01_LC_8_4_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIHIN01_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIHIN01_LC_8_4_0 .LUT_INIT=16'b1111010111000101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIHIN01_LC_8_4_0  (
            .in0(N__25754),
            .in1(N__29714),
            .in2(N__35495),
            .in3(N__30559),
            .lcout(\POWERLED.N_452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_4_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__35491),
            .in2(_gnd_net_),
            .in3(N__30853),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_8_4_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_8_4_4 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__24260),
            .in2(N__24302),
            .in3(N__29119),
            .lcout(RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34465),
            .ce(N__24040),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_8_4_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_8_4_5 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_8_4_5  (
            .in0(N__24261),
            .in1(N__24283),
            .in2(N__29130),
            .in3(_gnd_net_),
            .lcout(RSMRSTn_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34465),
            .ce(N__24040),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_8_4_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_8_4_6 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(N__24262),
            .in2(N__24303),
            .in3(N__29123),
            .lcout(RSMRSTn_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34465),
            .ce(N__24040),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_8_4_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_8_4_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_8_4_7  (
            .in0(N__24263),
            .in1(N__24284),
            .in2(N__29131),
            .in3(N__24219),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34465),
            .ce(N__24040),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNI0RLU1_LC_8_5_0 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNI0RLU1_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNI0RLU1_LC_8_5_0 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \COUNTER.tmp_0_fast_RNI0RLU1_LC_8_5_0  (
            .in0(N__32385),
            .in1(N__27873),
            .in2(N__27799),
            .in3(N__23329),
            .lcout(\COUNTER.tmp_0_fast_RNI0RLUZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOI5P1_1_LC_8_5_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOI5P1_1_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOI5P1_1_LC_8_5_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \POWERLED.func_state_RNIOI5P1_1_LC_8_5_1  (
            .in0(N__23306),
            .in1(N__30033),
            .in2(N__23318),
            .in3(N__29679),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI81IE3_1_LC_8_5_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI81IE3_1_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI81IE3_1_LC_8_5_2 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \POWERLED.func_state_RNI81IE3_1_LC_8_5_2  (
            .in0(N__30710),
            .in1(_gnd_net_),
            .in2(N__23276),
            .in3(N__24877),
            .lcout(\POWERLED.N_413_N ),
            .ltout(\POWERLED.N_413_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITL8S5_0_LC_8_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITL8S5_0_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITL8S5_0_LC_8_5_3 .LUT_INIT=16'b0011111100111011;
    LogicCell40 \POWERLED.dutycycle_RNITL8S5_0_LC_8_5_3  (
            .in0(N__30390),
            .in1(N__33738),
            .in2(N__23372),
            .in3(N__30711),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_215_i_0_o2_LC_8_5_4 .C_ON=1'b0;
    defparam \POWERLED.N_215_i_0_o2_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_215_i_0_o2_LC_8_5_4 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \POWERLED.N_215_i_0_o2_LC_8_5_4  (
            .in0(N__32386),
            .in1(N__27874),
            .in2(N__27798),
            .in3(N__23328),
            .lcout(\POWERLED.N_430 ),
            .ltout(\POWERLED.N_430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITL8S5_2_LC_8_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITL8S5_2_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITL8S5_2_LC_8_5_5 .LUT_INIT=16'b0100111101011111;
    LogicCell40 \POWERLED.dutycycle_RNITL8S5_2_LC_8_5_5  (
            .in0(N__23360),
            .in1(N__30709),
            .in2(N__23345),
            .in3(N__27101),
            .lcout(\POWERLED.dutycycle_eena_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_en_LC_8_5_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_en_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_en_LC_8_5_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.func_state_en_LC_8_5_6  (
            .in0(N__24669),
            .in1(N__28055),
            .in2(_gnd_net_),
            .in3(N__29873),
            .lcout(\POWERLED.func_state_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_LC_8_5_7 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_fast_LC_8_5_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \COUNTER.tmp_0_fast_LC_8_5_7  (
            .in0(N__23330),
            .in1(_gnd_net_),
            .in2(N__29888),
            .in3(_gnd_net_),
            .lcout(SUSWARN_N_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34533),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_0_0_LC_8_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_0_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_0_0_LC_8_6_0 .LUT_INIT=16'b1100110111001111;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_0_0_LC_8_6_0  (
            .in0(N__24922),
            .in1(N__27338),
            .in2(N__35641),
            .in3(N__24718),
            .lcout(\POWERLED.un1_count_off_1_sqmuxa_8_m0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_7_1_LC_8_6_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_7_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_7_1_LC_8_6_1 .LUT_INIT=16'b0010011110101111;
    LogicCell40 \POWERLED.func_state_RNI_7_1_LC_8_6_1  (
            .in0(N__30002),
            .in1(N__24940),
            .in2(N__30658),
            .in3(N__24923),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_8_6_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_8_6_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \POWERLED.func_state_RNIMQ0F_1_LC_8_6_2  (
            .in0(N__27677),
            .in1(_gnd_net_),
            .in2(N__23309),
            .in3(N__31953),
            .lcout(\POWERLED.un1_count_off_1_sqmuxa_8_m1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNILKMD2_LC_8_6_3 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNILKMD2_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNILKMD2_LC_8_6_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \COUNTER.tmp_0_fast_RNILKMD2_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23300),
            .in3(N__30729),
            .lcout(N_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_0_LC_8_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_8_6_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_0_LC_8_6_4  (
            .in0(N__30358),
            .in1(N__30997),
            .in2(N__33056),
            .in3(N__25822),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNI_6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_0_LC_8_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_0_LC_8_6_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_0_LC_8_6_5  (
            .in0(N__30625),
            .in1(_gnd_net_),
            .in2(N__23399),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_10Z0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNI_10Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_8_6_6 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_8_6_6  (
            .in0(N__27396),
            .in1(N__24929),
            .in2(N__23396),
            .in3(N__24717),
            .lcout(\POWERLED.N_676 ),
            .ltout(\POWERLED.N_676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI99TE_1_LC_8_6_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI99TE_1_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI99TE_1_LC_8_6_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI99TE_1_LC_8_6_7  (
            .in0(N__32598),
            .in1(N__35085),
            .in2(N__23393),
            .in3(N__27676),
            .lcout(\POWERLED.N_492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_0_LC_8_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_0_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_0_LC_8_7_0 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \POWERLED.dutycycle_RNI_13_0_LC_8_7_0  (
            .in0(N__35635),
            .in1(N__23449),
            .in2(N__29681),
            .in3(N__30054),
            .lcout(\POWERLED.dutycycle_RNI_13Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNILKMD2_1_LC_8_7_1 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNILKMD2_1_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNILKMD2_1_LC_8_7_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \COUNTER.tmp_0_fast_RNILKMD2_1_LC_8_7_1  (
            .in0(N__23560),
            .in1(N__25710),
            .in2(_gnd_net_),
            .in3(N__35633),
            .lcout(G_11_i_a10_0_1),
            .ltout(G_11_i_a10_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNI2Q8O5_LC_8_7_2 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNI2Q8O5_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNI2Q8O5_LC_8_7_2 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \COUNTER.tmp_0_fast_RNI2Q8O5_LC_8_7_2  (
            .in0(N__25709),
            .in1(N__30089),
            .in2(N__23390),
            .in3(N__23378),
            .lcout(),
            .ltout(N_9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKJI1H_1_LC_8_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKJI1H_1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKJI1H_1_LC_8_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNIKJI1H_1_LC_8_7_3  (
            .in0(N__23387),
            .in1(N__23486),
            .in2(N__23381),
            .in3(N__24989),
            .lcout(\POWERLED.g0_i_o4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_0_LC_8_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_0_LC_8_7_4 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \POWERLED.dutycycle_RNI_12_0_LC_8_7_4  (
            .in0(N__35634),
            .in1(N__23448),
            .in2(N__29680),
            .in3(N__30053),
            .lcout(N_8_3),
            .ltout(N_8_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBFNS2_1_LC_8_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBFNS2_1_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBFNS2_1_LC_8_7_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNIBFNS2_1_LC_8_7_5  (
            .in0(N__27437),
            .in1(N__23495),
            .in2(N__23489),
            .in3(N__25874),
            .lcout(\POWERLED.N_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_0_LC_8_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_0_LC_8_7_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.dutycycle_RNI_14_0_LC_8_7_6  (
            .in0(N__35636),
            .in1(N__23450),
            .in2(_gnd_net_),
            .in3(N__30055),
            .lcout(\POWERLED.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_1_LC_8_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_8_7_7 .LUT_INIT=16'b0101010100000001;
    LogicCell40 \POWERLED.dutycycle_RNI_1_1_LC_8_7_7  (
            .in0(N__24958),
            .in1(N__25875),
            .in2(N__23564),
            .in3(N__35637),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_8_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_8_8_0 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_8_8_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \POWERLED.dutycycle_5_LC_8_8_0  (
            .in0(N__23474),
            .in1(N__24844),
            .in2(N__25010),
            .in3(N__23464),
            .lcout(\POWERLED.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__31543));
    defparam \POWERLED.dutycycle_RNIH61711_5_LC_8_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIH61711_5_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIH61711_5_LC_8_8_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \POWERLED.dutycycle_RNIH61711_5_LC_8_8_1  (
            .in0(N__24845),
            .in1(N__23473),
            .in2(N__23465),
            .in3(N__25000),
            .lcout(\POWERLED.dutycycleZ1Z_5 ),
            .ltout(\POWERLED.dutycycleZ1Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_0_LC_8_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_8_8_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_0_LC_8_8_2  (
            .in0(N__33089),
            .in1(N__30420),
            .in2(N__23453),
            .in3(N__25871),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_0_LC_8_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_8_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_0_LC_8_8_3  (
            .in0(N__23421),
            .in1(N__30419),
            .in2(N__33145),
            .in3(N__25870),
            .lcout(\POWERLED.N_546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_8_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_8_8_4 .LUT_INIT=16'b1110110011001000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_8_8_4  (
            .in0(N__32257),
            .in1(N__31415),
            .in2(N__31258),
            .in3(N__32849),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_LC_8_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_5_LC_8_8_5  (
            .in0(N__30984),
            .in1(N__33088),
            .in2(N__23438),
            .in3(N__31811),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_0_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_8_8_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_0_LC_8_8_6  (
            .in0(N__30418),
            .in1(N__33128),
            .in2(_gnd_net_),
            .in3(N__23420),
            .lcout(N_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_3_LC_8_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_3_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_3_LC_8_8_7 .LUT_INIT=16'b0100010101011101;
    LogicCell40 \POWERLED.dutycycle_RNI_11_3_LC_8_8_7  (
            .in0(N__31414),
            .in1(N__33087),
            .in2(N__32271),
            .in3(N__31245),
            .lcout(\POWERLED.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_8_9_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_13_LC_8_9_1  (
            .in0(N__23537),
            .in1(N__26036),
            .in2(N__23531),
            .in3(N__29531),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34592),
            .ce(),
            .sr(N__31556));
    defparam \POWERLED.dutycycle_RNI99TE_13_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI99TE_13_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI99TE_13_LC_8_9_2 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \POWERLED.dutycycle_RNI99TE_13_LC_8_9_2  (
            .in0(N__32591),
            .in1(N__23512),
            .in2(_gnd_net_),
            .in3(N__35126),
            .lcout(),
            .ltout(\POWERLED.N_598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI9B7B1_13_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI9B7B1_13_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI9B7B1_13_LC_8_9_3 .LUT_INIT=16'b1100111000000010;
    LogicCell40 \POWERLED.dutycycle_RNI9B7B1_13_LC_8_9_3  (
            .in0(N__31887),
            .in1(N__27683),
            .in2(N__23543),
            .in3(N__26227),
            .lcout(),
            .ltout(\POWERLED.N_450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5FJ65_13_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5FJ65_13_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5FJ65_13_LC_8_9_4 .LUT_INIT=16'b0010001010100010;
    LogicCell40 \POWERLED.dutycycle_RNI5FJ65_13_LC_8_9_4  (
            .in0(N__33544),
            .in1(N__33802),
            .in2(N__23540),
            .in3(N__30832),
            .lcout(\POWERLED.dutycycle_RNI5FJ65Z0Z_13 ),
            .ltout(\POWERLED.dutycycle_RNI5FJ65Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIT3QT5_13_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIT3QT5_13_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIT3QT5_13_LC_8_9_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \POWERLED.dutycycle_RNIT3QT5_13_LC_8_9_5  (
            .in0(N__23527),
            .in1(N__26035),
            .in2(N__23519),
            .in3(N__29530),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(\POWERLED.dutycycleZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_13_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_8_9_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_13_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23516),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2336_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIT70K5_8_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIT70K5_8_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIT70K5_8_LC_8_9_7 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \POWERLED.dutycycle_RNIT70K5_8_LC_8_9_7  (
            .in0(N__23501),
            .in1(N__33795),
            .in2(N__30833),
            .in3(N__33543),
            .lcout(\POWERLED.dutycycle_RNIT70K5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_8_10_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_12_LC_8_10_0  (
            .in0(N__26050),
            .in1(N__28436),
            .in2(N__33642),
            .in3(N__23603),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34582),
            .ce(),
            .sr(N__31589));
    defparam \POWERLED.dutycycle_RNI_6_8_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_8_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_8_LC_8_10_1 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \POWERLED.dutycycle_RNI_6_8_LC_8_10_1  (
            .in0(N__26119),
            .in1(N__31217),
            .in2(N__32853),
            .in3(N__27724),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_8_10_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_8_10_2  (
            .in0(N__28181),
            .in1(_gnd_net_),
            .in2(N__31809),
            .in3(N__28495),
            .lcout(),
            .ltout(\POWERLED.un1_m2_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_8_LC_8_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_8_10_3 .LUT_INIT=16'b1110000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_8_LC_8_10_3  (
            .in0(N__32837),
            .in1(N__23789),
            .in2(N__23612),
            .in3(N__31219),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIGQPC6_12_LC_8_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIGQPC6_12_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIGQPC6_12_LC_8_10_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNIGQPC6_12_LC_8_10_4  (
            .in0(N__33582),
            .in1(N__23602),
            .in2(N__26051),
            .in3(N__28435),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(\POWERLED.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_8_10_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__28180),
            .in2(N__23594),
            .in3(N__31769),
            .lcout(\POWERLED.un1_dutycycle_53_56_a1_2 ),
            .ltout(\POWERLED.un1_dutycycle_53_56_a1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_8_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_8_10_6 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_8_LC_8_10_6  (
            .in0(N__31218),
            .in1(N__27725),
            .in2(N__23591),
            .in3(N__32836),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_3Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_8_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_8_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_8_LC_8_10_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_8_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__23790),
            .in2(N__23588),
            .in3(N__23585),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM3TC6_15_LC_8_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM3TC6_15_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM3TC6_15_LC_8_11_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIM3TC6_15_LC_8_11_0  (
            .in0(N__23572),
            .in1(N__29508),
            .in2(N__33455),
            .in3(N__25930),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_8_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_8_11_1 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \POWERLED.dutycycle_15_LC_8_11_1  (
            .in0(N__25931),
            .in1(N__33451),
            .in2(N__29538),
            .in3(N__23573),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34678),
            .ce(),
            .sr(N__31569));
    defparam \POWERLED.dutycycle_8_LC_8_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_8_11_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \POWERLED.dutycycle_8_LC_8_11_2  (
            .in0(N__23642),
            .in1(N__29510),
            .in2(N__23654),
            .in3(N__25732),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34678),
            .ce(),
            .sr(N__31569));
    defparam \POWERLED.dutycycle_RNI_3_10_LC_8_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_8_11_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_10_LC_8_11_3  (
            .in0(N__33134),
            .in1(N__31402),
            .in2(N__32957),
            .in3(N__28278),
            .lcout(\POWERLED.g0_9_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_10_LC_8_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_8_11_4 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_10_LC_8_11_4  (
            .in0(N__33133),
            .in1(N__31215),
            .in2(N__28298),
            .in3(N__32942),
            .lcout(\POWERLED.N_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIT1OR5_8_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIT1OR5_8_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIT1OR5_8_LC_8_11_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \POWERLED.dutycycle_RNIT1OR5_8_LC_8_11_5  (
            .in0(N__29509),
            .in1(N__23650),
            .in2(N__25733),
            .in3(N__23641),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(\POWERLED.dutycycleZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_8_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_8_11_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_8_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23630),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_8 ),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_8_11_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__33132),
            .in2(N__23627),
            .in3(N__31401),
            .lcout(\POWERLED.N_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_8_12_0 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_8_12_0  (
            .in0(N__33136),
            .in1(N__31404),
            .in2(N__31253),
            .in3(N__32273),
            .lcout(),
            .ltout(\POWERLED.N_6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_8_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_8_12_1  (
            .in0(N__28166),
            .in1(N__31756),
            .in2(N__23624),
            .in3(N__32845),
            .lcout(),
            .ltout(\POWERLED.N_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_3_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_3_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_3_LC_8_12_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \POWERLED.dutycycle_RNI_15_3_LC_8_12_2  (
            .in0(N__23672),
            .in1(N__23621),
            .in2(N__23615),
            .in3(N__26315),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_15Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_8_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_8_12_3  (
            .in0(N__28167),
            .in1(N__31086),
            .in2(N__23696),
            .in3(N__28511),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_12_4 .LUT_INIT=16'b1100000011111100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_6_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__33135),
            .in2(N__31798),
            .in3(N__31121),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_10_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_8_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_10_LC_8_12_5  (
            .in0(N__28284),
            .in1(N__33137),
            .in2(N__23684),
            .in3(N__32844),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHDMC5_10_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHDMC5_10_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHDMC5_10_LC_8_12_6 .LUT_INIT=16'b0101010101110101;
    LogicCell40 \POWERLED.dutycycle_RNIHDMC5_10_LC_8_12_6  (
            .in0(N__33817),
            .in1(N__28214),
            .in2(N__27755),
            .in3(N__33437),
            .lcout(\POWERLED.dutycycle_RNIHDMC5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__32258),
            .in2(_gnd_net_),
            .in3(N__31226),
            .lcout(\POWERLED.N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_8_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_8_13_0 .LUT_INIT=16'b1100110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_8_13_0  (
            .in0(N__34937),
            .in1(N__26233),
            .in2(N__25922),
            .in3(N__23768),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_8_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_8_13_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \POWERLED.dutycycle_14_LC_8_13_1  (
            .in0(N__25949),
            .in1(N__23762),
            .in2(N__29571),
            .in3(N__28087),
            .lcout(\POWERLED.dutycycleZ1Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34676),
            .ce(),
            .sr(N__31570));
    defparam \POWERLED.dutycycle_RNI_7_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_LC_8_13_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32854),
            .in3(N__25899),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_12_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_13_LC_8_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_8_13_4 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_13_LC_8_13_4  (
            .in0(N__25918),
            .in1(N__26232),
            .in2(N__23657),
            .in3(N__23792),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_8_LC_8_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_8_13_5 .LUT_INIT=16'b0000010001001100;
    LogicCell40 \POWERLED.dutycycle_RNI_5_8_LC_8_13_5  (
            .in0(N__23791),
            .in1(N__25900),
            .in2(N__32855),
            .in3(N__31244),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIK0SC6_14_LC_8_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIK0SC6_14_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIK0SC6_14_LC_8_13_6 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIK0SC6_14_LC_8_13_6  (
            .in0(N__23761),
            .in1(N__29555),
            .in2(N__28088),
            .in3(N__25948),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(\POWERLED.dutycycleZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_15_LC_8_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_8_13_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_15_LC_8_13_7  (
            .in0(N__31109),
            .in1(_gnd_net_),
            .in2(N__23753),
            .in3(N__23749),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI4QQA4_13_LC_8_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI4QQA4_13_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI4QQA4_13_LC_8_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI4QQA4_13_LC_8_14_0  (
            .in0(N__23729),
            .in1(N__33956),
            .in2(_gnd_net_),
            .in3(N__23908),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_8_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_8_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_13_LC_8_14_1  (
            .in0(N__23909),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34656),
            .ce(N__33935),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIFIL44_1_LC_8_14_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFIL44_1_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFIL44_1_LC_8_14_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.func_state_RNIFIL44_1_LC_8_14_2  (
            .in0(N__27149),
            .in1(N__28022),
            .in2(N__33669),
            .in3(N__23723),
            .lcout(\POWERLED.count_clk_en ),
            .ltout(\POWERLED.count_clk_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI0GFI4_2_LC_8_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI0GFI4_2_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI0GFI4_2_LC_8_14_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \POWERLED.count_clk_RNI0GFI4_2_LC_8_14_3  (
            .in0(N__23861),
            .in1(_gnd_net_),
            .in2(N__23711),
            .in3(N__23708),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_8_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_8_14_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \POWERLED.count_clk_2_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__23860),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34656),
            .ce(N__33935),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_8_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_8_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_15_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23887),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34656),
            .ce(N__33935),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI80TA4_15_LC_8_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI80TA4_15_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI80TA4_15_LC_8_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_clk_RNI80TA4_15_LC_8_14_6  (
            .in0(N__23888),
            .in1(N__23702),
            .in2(_gnd_net_),
            .in3(N__33957),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_8_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_8_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_4_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23842),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34656),
            .ce(N__33935),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_8_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_8_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__28676),
            .in2(N__34880),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_8_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_8_15_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_8_15_1  (
            .in0(N__34815),
            .in1(N__26477),
            .in2(_gnd_net_),
            .in3(N__23852),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_8_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_8_15_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_8_15_2  (
            .in0(N__34809),
            .in1(N__26342),
            .in2(_gnd_net_),
            .in3(N__23849),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_8_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_8_15_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_8_15_3  (
            .in0(N__34812),
            .in1(N__26507),
            .in2(_gnd_net_),
            .in3(N__23828),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_8_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_8_15_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_8_15_4  (
            .in0(N__34810),
            .in1(N__26763),
            .in2(_gnd_net_),
            .in3(N__23825),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_8_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_8_15_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_8_15_5  (
            .in0(N__34813),
            .in1(N__26529),
            .in2(_gnd_net_),
            .in3(N__23798),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_8_15_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_8_15_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_8_15_6  (
            .in0(N__34811),
            .in1(N__26406),
            .in2(_gnd_net_),
            .in3(N__23795),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_8_15_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_8_15_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_8_15_7  (
            .in0(N__34814),
            .in1(N__26542),
            .in2(_gnd_net_),
            .in3(N__23936),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_8_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_8_16_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_8_16_0  (
            .in0(N__34830),
            .in1(N__26749),
            .in2(_gnd_net_),
            .in3(N__23933),
            .lcout(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_8_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_8_16_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_8_16_1  (
            .in0(N__34832),
            .in1(N__23930),
            .in2(_gnd_net_),
            .in3(N__23918),
            .lcout(\POWERLED.count_clk_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_8_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_8_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__28363),
            .in2(_gnd_net_),
            .in3(N__23915),
            .lcout(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_8_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_8_16_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_8_16_3  (
            .in0(N__34833),
            .in1(N__26579),
            .in2(_gnd_net_),
            .in3(N__23912),
            .lcout(\POWERLED.count_clk_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_8_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_8_16_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_8_16_4  (
            .in0(N__34831),
            .in1(N__26710),
            .in2(_gnd_net_),
            .in3(N__23897),
            .lcout(\POWERLED.count_clk_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI6TRA4_LC_8_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI6TRA4_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI6TRA4_LC_8_16_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNI6TRA4_LC_8_16_5  (
            .in0(N__34834),
            .in1(N__23876),
            .in2(_gnd_net_),
            .in3(N__23894),
            .lcout(\POWERLED.count_clk_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_8_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_8_16_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_8_16_6  (
            .in0(N__26668),
            .in1(N__34835),
            .in2(_gnd_net_),
            .in3(N__23891),
            .lcout(\POWERLED.count_clk_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIUMD84_0_14_LC_8_16_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIUMD84_0_14_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIUMD84_0_14_LC_8_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIUMD84_0_14_LC_8_16_7  (
            .in0(N__33978),
            .in1(N__26797),
            .in2(_gnd_net_),
            .in3(N__26571),
            .lcout(\POWERLED.un1_count_clk_2_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIN0RE1_3_LC_9_1_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIN0RE1_3_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIN0RE1_3_LC_9_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIN0RE1_3_LC_9_1_0  (
            .in0(N__24376),
            .in1(N__24304),
            .in2(N__24365),
            .in3(N__24349),
            .lcout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_1_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_1_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_1_1  (
            .in0(N__24307),
            .in1(N__29116),
            .in2(_gnd_net_),
            .in3(N__24245),
            .lcout(),
            .ltout(\RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_1_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_1_2 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_9_1_2  (
            .in0(N__24247),
            .in1(_gnd_net_),
            .in2(N__24326),
            .in3(N__24221),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34399),
            .ce(N__24028),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_1_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_1_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_1_3  (
            .in0(N__24305),
            .in1(N__29118),
            .in2(_gnd_net_),
            .in3(N__24243),
            .lcout(\RSMRST_PWRGD.N_264_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_1_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_1_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_LC_9_1_4  (
            .in0(N__24246),
            .in1(N__29115),
            .in2(_gnd_net_),
            .in3(N__24308),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34399),
            .ce(N__24028),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_1_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_1_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_1_5  (
            .in0(N__24306),
            .in1(N__29117),
            .in2(_gnd_net_),
            .in3(N__24242),
            .lcout(),
            .ltout(\RSMRST_PWRGD.N_555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__G_14_LC_9_1_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__G_14_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__G_14_LC_9_1_6 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__G_14_LC_9_1_6  (
            .in0(N__24244),
            .in1(N__24220),
            .in2(N__24197),
            .in3(N__24130),
            .lcout(\RSMRST_PWRGD.G_14 ),
            .ltout(\RSMRST_PWRGD.G_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_1_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_1_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_1_7  (
            .in0(N__24131),
            .in1(_gnd_net_),
            .in2(N__23960),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.N_92_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIB4D36_1_LC_9_2_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIB4D36_1_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIB4D36_1_LC_9_2_0 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \POWERLED.func_state_RNIB4D36_1_LC_9_2_0  (
            .in0(N__35472),
            .in1(N__32676),
            .in2(N__26907),
            .in3(N__29186),
            .lcout(\POWERLED.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIOTGO_10_LC_9_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIOTGO_10_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIOTGO_10_LC_9_2_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \POWERLED.count_off_RNIOTGO_10_LC_9_2_1  (
            .in0(N__32394),
            .in1(N__30742),
            .in2(N__30577),
            .in3(N__29261),
            .lcout(\POWERLED.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_0_0_o2_0_LC_9_2_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_0_0_o2_0_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_0_0_o2_0_LC_9_2_2 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_0_0_o2_0_LC_9_2_2  (
            .in0(N__35470),
            .in1(N__32674),
            .in2(_gnd_net_),
            .in3(N__27806),
            .lcout(\POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_18_LC_9_2_3 .C_ON=1'b0;
    defparam \POWERLED.g0_18_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_18_LC_9_2_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.g0_18_LC_9_2_3  (
            .in0(N__27807),
            .in1(N__35473),
            .in2(N__32681),
            .in3(N__32395),
            .lcout(),
            .ltout(\POWERLED.N_423_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI7KPT2_1_LC_9_2_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI7KPT2_1_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI7KPT2_1_LC_9_2_4 .LUT_INIT=16'b1101000000000000;
    LogicCell40 \POWERLED.func_state_RNI7KPT2_1_LC_9_2_4  (
            .in0(N__30561),
            .in1(N__27316),
            .in2(N__24401),
            .in3(N__33369),
            .lcout(\POWERLED.N_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_LC_9_2_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_9_2_5 .LUT_INIT=16'b0110011001000100;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_LC_9_2_5  (
            .in0(N__32675),
            .in1(N__35471),
            .in2(_gnd_net_),
            .in3(N__29294),
            .lcout(),
            .ltout(\POWERLED.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJ2SL7_1_LC_9_2_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJ2SL7_1_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJ2SL7_1_LC_9_2_6 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \POWERLED.func_state_RNIJ2SL7_1_LC_9_2_6  (
            .in0(N__29961),
            .in1(N__30277),
            .in2(N__24398),
            .in3(N__24395),
            .lcout(),
            .ltout(\POWERLED.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICVMGB_1_LC_9_2_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICVMGB_1_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICVMGB_1_LC_9_2_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.func_state_RNICVMGB_1_LC_9_2_7  (
            .in0(N__24389),
            .in1(N__32003),
            .in2(N__24383),
            .in3(N__29889),
            .lcout(\POWERLED.g0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDNS62_1_LC_9_3_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDNS62_1_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDNS62_1_LC_9_3_0 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \POWERLED.func_state_RNIDNS62_1_LC_9_3_0  (
            .in0(N__29185),
            .in1(N__27317),
            .in2(N__28067),
            .in3(N__30560),
            .lcout(),
            .ltout(\POWERLED.N_541_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6NN75_1_LC_9_3_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6NN75_1_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6NN75_1_LC_9_3_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.func_state_RNI6NN75_1_LC_9_3_1  (
            .in0(N__24797),
            .in1(N__33776),
            .in2(N__24380),
            .in3(N__24806),
            .lcout(\POWERLED.N_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_9_3_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_9_3_2 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \POWERLED.func_state_0_LC_9_3_2  (
            .in0(N__24737),
            .in1(N__24752),
            .in2(N__24776),
            .in3(N__24782),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34326),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIP4521_1_LC_9_3_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIP4521_1_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIP4521_1_LC_9_3_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.func_state_RNIP4521_1_LC_9_3_3  (
            .in0(N__24683),
            .in1(N__35049),
            .in2(N__27896),
            .in3(N__33364),
            .lcout(\POWERLED.N_542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8KQ72_0_LC_9_3_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8KQ72_0_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8KQ72_0_LC_9_3_4 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \POWERLED.func_state_RNI8KQ72_0_LC_9_3_4  (
            .in0(N__24791),
            .in1(N__24824),
            .in2(_gnd_net_),
            .in3(N__29885),
            .lcout(\POWERLED.g2 ),
            .ltout(\POWERLED.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIGC9OO_0_LC_9_3_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIGC9OO_0_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIGC9OO_0_LC_9_3_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \POWERLED.func_state_RNIGC9OO_0_LC_9_3_5  (
            .in0(N__24763),
            .in1(N__24751),
            .in2(N__24740),
            .in3(N__24736),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(\POWERLED.func_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_9_3_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_9_3_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24722),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2291_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_9_3_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_9_3_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_9_3_7  (
            .in0(N__27389),
            .in1(N__24928),
            .in2(_gnd_net_),
            .in3(N__24719),
            .lcout(\POWERLED.func_state_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_430_i_LC_9_4_0 .C_ON=1'b0;
    defparam \POWERLED.N_430_i_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_430_i_LC_9_4_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.N_430_i_LC_9_4_0  (
            .in0(N__32352),
            .in1(N__24698),
            .in2(N__27895),
            .in3(N__35050),
            .lcout(\POWERLED.N_430_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_7_o3_LC_9_4_1 .C_ON=1'b0;
    defparam \POWERLED.g0_7_o3_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_7_o3_LC_9_4_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.g0_7_o3_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__35481),
            .in2(_gnd_net_),
            .in3(N__27797),
            .lcout(),
            .ltout(\POWERLED.N_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1PE62_1_LC_9_4_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1PE62_1_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1PE62_1_LC_9_4_2 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \POWERLED.func_state_RNI1PE62_1_LC_9_4_2  (
            .in0(N__27332),
            .in1(N__33366),
            .in2(N__24416),
            .in3(N__30539),
            .lcout(\POWERLED.N_16_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8H551_9_LC_9_4_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8H551_9_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8H551_9_LC_9_4_3 .LUT_INIT=16'b0011101100110011;
    LogicCell40 \POWERLED.dutycycle_RNI8H551_9_LC_9_4_3  (
            .in0(N__32657),
            .in1(N__35480),
            .in2(N__32384),
            .in3(N__31822),
            .lcout(),
            .ltout(\POWERLED.dutycycle_e_N_3L4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_9_LC_9_4_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_9_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_9_LC_9_4_4 .LUT_INIT=16'b1011000010111010;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_9_LC_9_4_4  (
            .in0(N__31823),
            .in1(N__33368),
            .in2(N__24827),
            .in3(N__30271),
            .lcout(\POWERLED.dutycycle_RNI6SKJ1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_8_0_LC_9_4_5 .C_ON=1'b0;
    defparam \POWERLED.g0_8_0_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_8_0_LC_9_4_5 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \POWERLED.g0_8_0_LC_9_4_5  (
            .in0(N__32658),
            .in1(N__29960),
            .in2(N__35490),
            .in3(N__30260),
            .lcout(\POWERLED.g0_8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_9_4_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_9_4_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(N__33367),
            .in2(_gnd_net_),
            .in3(N__30540),
            .lcout(\POWERLED.N_435 ),
            .ltout(\POWERLED.N_435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_1_LC_9_4_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_9_4_7 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_9_4_7  (
            .in0(N__33365),
            .in1(N__24924),
            .in2(N__24818),
            .in3(N__24815),
            .lcout(\POWERLED.func_state_1_m2s2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_9_5_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_9_5_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_9_5_0  (
            .in0(N__33361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29262),
            .lcout(\POWERLED.func_state_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_5_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_5_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_5_1  (
            .in0(N__27348),
            .in1(N__27985),
            .in2(N__30644),
            .in3(N__33363),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_m1_0_a2_LC_9_5_2 .C_ON=1'b0;
    defparam \POWERLED.un1_m1_0_a2_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_m1_0_a2_LC_9_5_2 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \POWERLED.un1_m1_0_a2_LC_9_5_2  (
            .in0(N__32655),
            .in1(N__35450),
            .in2(N__32402),
            .in3(N__30264),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_0_a2_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_215_i_0_o2_0_LC_9_5_3 .C_ON=1'b0;
    defparam \POWERLED.N_215_i_0_o2_0_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_215_i_0_o2_0_LC_9_5_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.N_215_i_0_o2_0_LC_9_5_3  (
            .in0(N__35449),
            .in1(N__32654),
            .in2(N__35144),
            .in3(N__32387),
            .lcout(),
            .ltout(\POWERLED.N_423_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRQ4D3_0_LC_9_5_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRQ4D3_0_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRQ4D3_0_LC_9_5_4 .LUT_INIT=16'b1010111100101111;
    LogicCell40 \POWERLED.func_state_RNIRQ4D3_0_LC_9_5_4  (
            .in0(N__30576),
            .in1(N__27347),
            .in2(N__24800),
            .in3(N__28056),
            .lcout(\POWERLED.N_688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDNFD1_1_LC_9_5_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDNFD1_1_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDNFD1_1_LC_9_5_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.func_state_RNIDNFD1_1_LC_9_5_5  (
            .in0(N__29710),
            .in1(N__33360),
            .in2(N__27886),
            .in3(N__30574),
            .lcout(\POWERLED.N_545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.VCCST_EN_i_0_o2_LC_9_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.VCCST_EN_i_0_o2_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.VCCST_EN_i_0_o2_LC_9_5_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \PCH_PWRGD.VCCST_EN_i_0_o2_LC_9_5_6  (
            .in0(N__32653),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30854),
            .lcout(VCCST_EN_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRKB61_1_LC_9_5_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRKB61_1_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRKB61_1_LC_9_5_7 .LUT_INIT=16'b0000101100001010;
    LogicCell40 \POWERLED.func_state_RNIRKB61_1_LC_9_5_7  (
            .in0(N__35213),
            .in1(N__33362),
            .in2(N__30797),
            .in3(N__30575),
            .lcout(\POWERLED.N_252_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_6_LC_9_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_9_6_0 .LUT_INIT=16'b0000100100000101;
    LogicCell40 \POWERLED.dutycycle_RNI_3_6_LC_9_6_0  (
            .in0(N__33052),
            .in1(N__24944),
            .in2(N__33371),
            .in3(N__24921),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI12AS_6_LC_9_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI12AS_6_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI12AS_6_LC_9_6_1 .LUT_INIT=16'b1000000001111111;
    LogicCell40 \POWERLED.dutycycle_RNI12AS_6_LC_9_6_1  (
            .in0(N__32633),
            .in1(N__30275),
            .in2(N__24881),
            .in3(N__33051),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI9S7D5_6_LC_9_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI9S7D5_6_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI9S7D5_6_LC_9_6_2 .LUT_INIT=16'b0000001011111111;
    LogicCell40 \POWERLED.dutycycle_RNI9S7D5_6_LC_9_6_2  (
            .in0(N__27254),
            .in1(N__24878),
            .in2(N__24863),
            .in3(N__33735),
            .lcout(\POWERLED.dutycycle_eena_13 ),
            .ltout(\POWERLED.dutycycle_eena_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIH1T5A_6_LC_9_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIH1T5A_6_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIH1T5A_6_LC_9_6_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \POWERLED.dutycycle_RNIH1T5A_6_LC_9_6_3  (
            .in0(N__25052),
            .in1(N__25036),
            .in2(N__24860),
            .in3(N__33634),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIIFNR3_LC_9_6_4 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIIFNR3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIIFNR3_LC_9_6_4 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIIFNR3_LC_9_6_4  (
            .in0(N__24833),
            .in1(N__24857),
            .in2(_gnd_net_),
            .in3(N__33736),
            .lcout(\POWERLED.dutycycle_set_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI12AS_1_LC_9_6_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI12AS_1_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI12AS_1_LC_9_6_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \POWERLED.func_state_RNI12AS_1_LC_9_6_5  (
            .in0(N__32634),
            .in1(N__33349),
            .in2(_gnd_net_),
            .in3(N__30276),
            .lcout(\POWERLED.func_state_RNI12ASZ0Z_1 ),
            .ltout(\POWERLED.func_state_RNI12ASZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHOR3_LC_9_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHOR3_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHOR3_LC_9_6_6 .LUT_INIT=16'b0000001111111111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHOR3_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__27116),
            .in2(N__25055),
            .in3(N__33737),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3 ),
            .ltout(\POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_9_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_9_6_7 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_9_6_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_6_LC_9_6_7  (
            .in0(N__25046),
            .in1(N__25037),
            .in2(N__25040),
            .in3(N__33635),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34451),
            .ce(),
            .sr(N__31563));
    defparam \POWERLED.dutycycle_RNI_1_0_LC_9_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_9_7_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_0_LC_9_7_0  (
            .in0(N__30415),
            .in1(N__27269),
            .in2(N__25880),
            .in3(N__25028),
            .lcout(\POWERLED.N_2363_0 ),
            .ltout(\POWERLED.N_2363_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_0_LC_9_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_0_LC_9_7_1 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_15_0_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25022),
            .in3(N__35625),
            .lcout(\POWERLED.N_12_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNILKMD2_0_LC_9_7_2 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNILKMD2_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNILKMD2_0_LC_9_7_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \COUNTER.tmp_0_fast_RNILKMD2_0_LC_9_7_2  (
            .in0(N__30311),
            .in1(N__25712),
            .in2(_gnd_net_),
            .in3(N__25876),
            .lcout(),
            .ltout(G_11_i_a10_2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO453C_5_LC_9_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO453C_5_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO453C_5_LC_9_7_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \POWERLED.dutycycle_RNIO453C_5_LC_9_7_3  (
            .in0(N__29624),
            .in1(N__25019),
            .in2(N__25013),
            .in3(N__25682),
            .lcout(\POWERLED.g2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNIGTMK4_LC_9_7_4 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNIGTMK4_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNIGTMK4_LC_9_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.tmp_0_fast_RNIGTMK4_LC_9_7_4  (
            .in0(N__25708),
            .in1(N__24983),
            .in2(N__24977),
            .in3(N__29623),
            .lcout(N_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_17_0_LC_9_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_17_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_17_0_LC_9_7_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_17_0_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__29641),
            .in2(_gnd_net_),
            .in3(N__29672),
            .lcout(N_7),
            .ltout(N_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_0_LC_9_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_0_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_0_LC_9_7_6 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_11_0_LC_9_7_6  (
            .in0(N__24976),
            .in1(N__30310),
            .in2(N__24962),
            .in3(N__24959),
            .lcout(),
            .ltout(\POWERLED.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI87EE7_5_LC_9_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI87EE7_5_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI87EE7_5_LC_9_7_7 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \POWERLED.dutycycle_RNI87EE7_5_LC_9_7_7  (
            .in0(N__29777),
            .in1(N__27436),
            .in2(N__25715),
            .in3(N__25707),
            .lcout(\POWERLED.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_1_LC_9_8_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_9_8_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_9_8_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \PCH_PWRGD.count_1_LC_9_8_0  (
            .in0(N__25676),
            .in1(N__25631),
            .in2(_gnd_net_),
            .in3(N__25407),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(N__25583),
            .sr(N__25408));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_9_8_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_9_8_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__25175),
            .in2(_gnd_net_),
            .in3(N__25214),
            .lcout(\POWERLED.mult1_un124_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25174),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_0_LC_9_8_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_0_LC_9_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_0_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25118),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_9_8_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_9_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27703),
            .lcout(\POWERLED.func_state_RNI_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_1_LC_9_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_1_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_1_LC_9_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_5_1_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30052),
            .lcout(\POWERLED.N_435_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_9_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30424),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__25873),
            .in2(N__26005),
            .in3(N__25766),
            .lcout(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__25983),
            .in2(N__30205),
            .in3(N__25763),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_9_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_9_3  (
            .in0(N__29570),
            .in1(N__32250),
            .in2(N__26006),
            .in3(N__25760),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__25987),
            .in2(N__31405),
            .in3(N__25757),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__25989),
            .in2(N__30996),
            .in3(N__25742),
            .lcout(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_9_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__33106),
            .in2(N__26007),
            .in3(N__25739),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_9_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__25988),
            .in2(N__32822),
            .in3(N__25736),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__26008),
            .in2(N__31234),
            .in3(N__25721),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_10_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_10_1  (
            .in0(N__29568),
            .in1(N__26019),
            .in2(N__31807),
            .in3(N__25718),
            .lcout(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_10_2  (
            .in0(N__29567),
            .in1(N__26010),
            .in2(N__28308),
            .in3(N__26057),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_10_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_10_3  (
            .in0(N__29569),
            .in1(N__26020),
            .in2(N__28179),
            .in3(N__26054),
            .lcout(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_10_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_10_4  (
            .in0(N__29566),
            .in1(N__26009),
            .in2(N__28509),
            .in3(N__26039),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__26021),
            .in2(N__26238),
            .in3(N__26024),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__26011),
            .in2(N__34970),
            .in3(N__25937),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_10_7  (
            .in0(N__31104),
            .in1(N__30068),
            .in2(_gnd_net_),
            .in3(N__25934),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_12_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_9_11_0 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_12_LC_9_11_0  (
            .in0(N__28272),
            .in1(N__28163),
            .in2(N__28510),
            .in3(N__26156),
            .lcout(\POWERLED.un1_dutycycle_53_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_9_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_9_11_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.dutycycle_11_LC_9_11_1  (
            .in0(N__28325),
            .in1(N__33658),
            .in2(N__26150),
            .in3(N__26137),
            .lcout(\POWERLED.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34596),
            .ce(),
            .sr(N__31568));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_11_2 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31810),
            .in3(N__28162),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_9_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_9_11_3 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__31773),
            .in2(N__28183),
            .in3(N__32940),
            .lcout(\POWERLED.un1_dutycycle_53_59_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6G5Q6_11_LC_9_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6G5Q6_11_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6G5Q6_11_LC_9_11_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNI6G5Q6_11_LC_9_11_4  (
            .in0(N__33657),
            .in1(N__26146),
            .in2(N__26138),
            .in3(N__28324),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_9_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_9_11_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_9_11_5  (
            .in0(N__31216),
            .in1(N__28491),
            .in2(N__26126),
            .in3(N__31774),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_12_LC_9_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_12_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_12_LC_9_11_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.dutycycle_RNI_6_12_LC_9_11_6  (
            .in0(N__32941),
            .in1(N__26093),
            .in2(N__26123),
            .in3(N__26120),
            .lcout(\POWERLED.un1_dutycycle_53_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_9_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_9_11_7 .LUT_INIT=16'b0000001111000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__28271),
            .in2(N__28182),
            .in3(N__28490),
            .lcout(\POWERLED.un1_dutycycle_53_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_9_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_9_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_9_12_0  (
            .in0(N__28280),
            .in1(N__28165),
            .in2(N__34967),
            .in3(N__26063),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_4_LC_9_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_9_12_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_4_LC_9_12_1  (
            .in0(N__31403),
            .in1(N__33107),
            .in2(N__32958),
            .in3(N__31750),
            .lcout(),
            .ltout(\POWERLED.G_7_i_a5_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_10_LC_9_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_10_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_10_LC_9_12_2 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_10_LC_9_12_2  (
            .in0(N__28279),
            .in1(N__32690),
            .in2(N__26075),
            .in3(N__31220),
            .lcout(),
            .ltout(\POWERLED.N_16_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_9_LC_9_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_9_12_3 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \POWERLED.dutycycle_RNI_1_9_LC_9_12_3  (
            .in0(N__26072),
            .in1(N__31751),
            .in2(N__26066),
            .in3(N__26348),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITRJC6_10_LC_9_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITRJC6_10_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITRJC6_10_LC_9_12_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \POWERLED.dutycycle_RNITRJC6_10_LC_9_12_4  (
            .in0(N__26284),
            .in1(N__26269),
            .in2(N__26302),
            .in3(N__33659),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(\POWERLED.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_9_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_9_12_5 .LUT_INIT=16'b1111100011100000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_9_12_5  (
            .in0(N__28164),
            .in1(N__31752),
            .in2(N__26318),
            .in3(N__26309),
            .lcout(\POWERLED.g0_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_9_LC_9_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_9_12_6 .LUT_INIT=16'b0000000011111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_9_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__32848),
            .in2(N__31797),
            .in3(N__32946),
            .lcout(\POWERLED.g0_9_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_9_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_9_12_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.dutycycle_10_LC_9_12_7  (
            .in0(N__26303),
            .in1(N__33660),
            .in2(N__26273),
            .in3(N__26285),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34708),
            .ce(),
            .sr(N__31585));
    defparam \POWERLED.dutycycle_RNI_0_8_LC_9_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_9_13_0 .LUT_INIT=16'b1111110111000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_8_LC_9_13_0  (
            .in0(N__27740),
            .in1(N__32852),
            .in2(N__31796),
            .in3(N__31243),
            .lcout(\POWERLED.un1_dutycycle_53_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHDMC5_9_LC_9_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHDMC5_9_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHDMC5_9_LC_9_13_1 .LUT_INIT=16'b0011001100111011;
    LogicCell40 \POWERLED.dutycycle_RNIHDMC5_9_LC_9_13_1  (
            .in0(N__26261),
            .in1(N__33818),
            .in2(N__31646),
            .in3(N__33436),
            .lcout(\POWERLED.dutycycle_RNIHDMC5Z0Z_9 ),
            .ltout(\POWERLED.dutycycle_RNIHDMC5Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_9_LC_9_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_9_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_9_LC_9_13_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_9_LC_9_13_2  (
            .in0(N__26393),
            .in1(N__26383),
            .in2(N__26246),
            .in3(N__33673),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34742),
            .ce(),
            .sr(N__31580));
    defparam \POWERLED.dutycycle_RNI_1_10_LC_9_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_9_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_10_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__28274),
            .in2(_gnd_net_),
            .in3(N__31746),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_9_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_9_13_4 .LUT_INIT=16'b1111000000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_9_13_4  (
            .in0(N__26243),
            .in1(N__26180),
            .in2(N__26174),
            .in3(N__31427),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKUPA6_9_LC_9_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKUPA6_9_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKUPA6_9_LC_9_13_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNIKUPA6_9_LC_9_13_5  (
            .in0(N__33672),
            .in1(N__26392),
            .in2(N__26384),
            .in3(N__26369),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_10_LC_9_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_10_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_10_LC_9_13_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_10_LC_9_13_6  (
            .in0(N__28273),
            .in1(N__32850),
            .in2(N__26363),
            .in3(N__31242),
            .lcout(),
            .ltout(\POWERLED.N_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_LC_9_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_LC_9_13_7 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \POWERLED.dutycycle_RNI_9_LC_9_13_7  (
            .in0(N__32851),
            .in1(N__31742),
            .in2(N__26360),
            .in3(N__26357),
            .lcout(\POWERLED.G_7_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINSEUC_7_LC_9_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINSEUC_7_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINSEUC_7_LC_9_14_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \POWERLED.count_clk_RNINSEUC_7_LC_9_14_0  (
            .in0(N__26462),
            .in1(N__26408),
            .in2(_gnd_net_),
            .in3(N__26450),
            .lcout(\POWERLED.count_clk_RNINSEUCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_9_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_9_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_3_LC_9_14_1  (
            .in0(N__26329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34737),
            .ce(N__33936),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2JGI4_3_LC_9_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2JGI4_3_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2JGI4_3_LC_9_14_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI2JGI4_3_LC_9_14_2  (
            .in0(N__26557),
            .in1(N__33944),
            .in2(_gnd_net_),
            .in3(N__26328),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(\POWERLED.count_clkZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_3_LC_9_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_3_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_3_LC_9_14_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \POWERLED.count_clk_RNI_3_LC_9_14_3  (
            .in0(N__26476),
            .in1(N__26549),
            .in2(N__26336),
            .in3(N__26506),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINSEUC_6_LC_9_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINSEUC_6_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINSEUC_6_LC_9_14_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.count_clk_RNINSEUC_6_LC_9_14_4  (
            .in0(N__26531),
            .in1(N__26407),
            .in2(N__26333),
            .in3(N__26449),
            .lcout(count_clk_RNINSEUC_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2JGI4_0_3_LC_9_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2JGI4_0_3_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2JGI4_0_3_LC_9_14_5 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \POWERLED.count_clk_RNI2JGI4_0_3_LC_9_14_5  (
            .in0(N__26330),
            .in1(N__26558),
            .in2(N__33985),
            .in3(N__26548),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2JGI4_1_3_LC_9_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2JGI4_1_3_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2JGI4_1_3_LC_9_14_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNI2JGI4_1_3_LC_9_14_6  (
            .in0(N__26530),
            .in1(N__26505),
            .in2(N__26480),
            .in3(N__26475),
            .lcout(\POWERLED.N_625 ),
            .ltout(\POWERLED.N_625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINSEUC_1_10_LC_9_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINSEUC_1_10_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINSEUC_1_10_LC_9_14_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \POWERLED.count_clk_RNINSEUC_1_10_LC_9_14_7  (
            .in0(N__26735),
            .in1(_gnd_net_),
            .in2(N__26456),
            .in3(N__26621),
            .lcout(\POWERLED.N_668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_9_15_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_9_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_5_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26417),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__33934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIE5NI4_9_LC_9_15_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIE5NI4_9_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIE5NI4_9_LC_9_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIE5NI4_9_LC_9_15_1  (
            .in0(N__33917),
            .in1(N__26432),
            .in2(_gnd_net_),
            .in3(N__26440),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(\POWERLED.count_clkZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINSEUC_0_10_LC_9_15_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINSEUC_0_10_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINSEUC_0_10_LC_9_15_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \POWERLED.count_clk_RNINSEUC_0_10_LC_9_15_2  (
            .in0(N__26764),
            .in1(N__26617),
            .in2(N__26453),
            .in3(N__28674),
            .lcout(\POWERLED.count_clk_RNINSEUC_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_9_15_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_9_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_9_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26441),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__33934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI6PII4_5_LC_9_15_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI6PII4_5_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI6PII4_5_LC_9_15_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI6PII4_5_LC_9_15_4  (
            .in0(N__26426),
            .in1(N__33915),
            .in2(_gnd_net_),
            .in3(N__26416),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAVKI4_7_LC_9_15_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAVKI4_7_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAVKI4_7_LC_9_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIAVKI4_7_LC_9_15_5  (
            .in0(N__33916),
            .in1(N__26720),
            .in2(_gnd_net_),
            .in3(N__26728),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(\POWERLED.count_clkZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_9_15_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_9_15_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_9_15_6  (
            .in0(N__26765),
            .in1(N__26750),
            .in2(N__26738),
            .in3(N__28675),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_9_15_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_9_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_7_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26729),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__33934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2NPA4_12_LC_9_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2NPA4_12_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2NPA4_12_LC_9_16_0 .LUT_INIT=16'b1110111111101100;
    LogicCell40 \POWERLED.count_clk_RNI2NPA4_12_LC_9_16_0  (
            .in0(N__26591),
            .in1(N__26714),
            .in2(N__33997),
            .in3(N__26600),
            .lcout(\POWERLED.un2_count_clk_17_0_o2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_9_16_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_9_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_12_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26590),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34738),
            .ce(N__34004),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINE7B4_10_LC_9_16_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINE7B4_10_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINE7B4_10_LC_9_16_2 .LUT_INIT=16'b1110111111101100;
    LogicCell40 \POWERLED.count_clk_RNINE7B4_10_LC_9_16_2  (
            .in0(N__26692),
            .in1(N__26672),
            .in2(N__33998),
            .in3(N__26650),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_o2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINSEUC_10_LC_9_16_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINSEUC_10_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINSEUC_10_LC_9_16_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNINSEUC_10_LC_9_16_3  (
            .in0(N__26630),
            .in1(N__26606),
            .in2(N__26624),
            .in3(N__28364),
            .lcout(\POWERLED.count_clk_RNINSEUCZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIUMD84_14_LC_9_16_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIUMD84_14_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIUMD84_14_LC_9_16_4 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \POWERLED.count_clk_RNIUMD84_14_LC_9_16_4  (
            .in0(N__33977),
            .in1(N__26798),
            .in2(N__34879),
            .in3(N__26573),
            .lcout(\POWERLED.un2_count_clk_17_0_o2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2NPA4_0_12_LC_9_16_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2NPA4_0_12_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2NPA4_0_12_LC_9_16_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI2NPA4_0_12_LC_9_16_5  (
            .in0(N__26599),
            .in1(N__33970),
            .in2(_gnd_net_),
            .in3(N__26589),
            .lcout(\POWERLED.un1_count_clk_2_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_9_16_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_9_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_14_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26572),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34738),
            .ce(N__34004),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_11_2_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_11_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_9_LC_11_2_0  (
            .in0(N__26846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34423),
            .ce(N__29412),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIH3EQ11_9_LC_11_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIH3EQ11_9_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIH3EQ11_9_LC_11_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIH3EQ11_9_LC_11_2_1  (
            .in0(N__29446),
            .in1(N__26786),
            .in2(_gnd_net_),
            .in3(N__26845),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(\POWERLED.count_offZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_10_LC_11_2_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_10_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_10_LC_11_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_10_LC_11_2_2  (
            .in0(N__26980),
            .in1(N__28699),
            .in2(N__26780),
            .in3(N__26827),
            .lcout(\POWERLED.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIQDJO11_10_LC_11_2_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIQDJO11_10_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIQDJO11_10_LC_11_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIQDJO11_10_LC_11_2_3  (
            .in0(N__29447),
            .in1(N__26777),
            .in2(_gnd_net_),
            .in3(N__26812),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_11_2_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_11_2_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_10_LC_11_2_4  (
            .in0(N__26813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34423),
            .ce(N__29412),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI5O1N11_12_LC_11_2_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI5O1N11_12_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI5O1N11_12_LC_11_2_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNI5O1N11_12_LC_11_2_5  (
            .in0(N__29448),
            .in1(N__26771),
            .in2(_gnd_net_),
            .in3(N__26965),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_11_2_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_11_2_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_12_LC_11_2_6  (
            .in0(N__26966),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34423),
            .ce(N__29412),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI9U3N11_14_LC_11_2_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI9U3N11_14_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI9U3N11_14_LC_11_2_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \POWERLED.count_off_RNI9U3N11_14_LC_11_2_7  (
            .in0(N__28619),
            .in1(_gnd_net_),
            .in2(N__29460),
            .in3(N__28636),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_11_3_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_11_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__28838),
            .in2(N__28964),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI3666G_LC_11_3_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI3666G_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI3666G_LC_11_3_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNI3666G_LC_11_3_1  (
            .in0(N__28926),
            .in1(_gnd_net_),
            .in2(N__28748),
            .in3(N__26876),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_11_3_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_11_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__27014),
            .in2(_gnd_net_),
            .in3(N__26873),
            .lcout(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_11_3_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_11_3_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27005),
            .in3(N__26870),
            .lcout(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI6C96G_LC_11_3_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI6C96G_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI6C96G_LC_11_3_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNI6C96G_LC_11_3_4  (
            .in0(N__28929),
            .in1(_gnd_net_),
            .in2(N__28763),
            .in3(N__26867),
            .lcout(\POWERLED.count_off_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI7EA6G_LC_11_3_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI7EA6G_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI7EA6G_LC_11_3_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNI7EA6G_LC_11_3_5  (
            .in0(N__28927),
            .in1(_gnd_net_),
            .in2(N__28772),
            .in3(N__26864),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI8GB6G_LC_11_3_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI8GB6G_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI8GB6G_LC_11_3_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNI8GB6G_LC_11_3_6  (
            .in0(N__28930),
            .in1(_gnd_net_),
            .in2(N__27236),
            .in3(N__26861),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI9IC6G_LC_11_3_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI9IC6G_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI9IC6G_LC_11_3_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNI9IC6G_LC_11_3_7  (
            .in0(N__28928),
            .in1(_gnd_net_),
            .in2(N__27203),
            .in3(N__26858),
            .lcout(\POWERLED.count_off_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIAKD6G_LC_11_4_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIAKD6G_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIAKD6G_LC_11_4_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNIAKD6G_LC_11_4_0  (
            .in0(N__28931),
            .in1(N__26855),
            .in2(_gnd_net_),
            .in3(N__26834),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIBME6G_LC_11_4_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIBME6G_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIBME6G_LC_11_4_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNIBME6G_LC_11_4_1  (
            .in0(N__28922),
            .in1(_gnd_net_),
            .in2(N__26831),
            .in3(N__26801),
            .lcout(\POWERLED.count_off_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIJSR4G_LC_11_4_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIJSR4G_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIJSR4G_LC_11_4_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNIJSR4G_LC_11_4_2  (
            .in0(N__28932),
            .in1(_gnd_net_),
            .in2(N__28700),
            .in3(N__26987),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIKUS4G_LC_11_4_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIKUS4G_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIKUS4G_LC_11_4_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNIKUS4G_LC_11_4_3  (
            .in0(N__28923),
            .in1(_gnd_net_),
            .in2(N__26984),
            .in3(N__26954),
            .lcout(\POWERLED.count_off_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIL0U4G_LC_11_4_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIL0U4G_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIL0U4G_LC_11_4_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNIL0U4G_LC_11_4_4  (
            .in0(N__28933),
            .in1(_gnd_net_),
            .in2(N__29042),
            .in3(N__26951),
            .lcout(\POWERLED.count_off_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIM2V4G_LC_11_4_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIM2V4G_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIM2V4G_LC_11_4_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNIM2V4G_LC_11_4_5  (
            .in0(N__28924),
            .in1(_gnd_net_),
            .in2(N__29033),
            .in3(N__26948),
            .lcout(\POWERLED.count_off_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIN405G_LC_11_4_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIN405G_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIN405G_LC_11_4_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIN405G_LC_11_4_6  (
            .in0(N__29009),
            .in1(N__28925),
            .in2(_gnd_net_),
            .in3(N__26945),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNIN405GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBH2F5_1_LC_11_5_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBH2F5_1_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBH2F5_1_LC_11_5_0 .LUT_INIT=16'b1110111110101010;
    LogicCell40 \POWERLED.func_state_RNIBH2F5_1_LC_11_5_0  (
            .in0(N__27092),
            .in1(N__26942),
            .in2(N__26930),
            .in3(N__33287),
            .lcout(),
            .ltout(\POWERLED.N_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIVO7PG_1_LC_11_5_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIVO7PG_1_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIVO7PG_1_LC_11_5_1 .LUT_INIT=16'b1100100011111011;
    LogicCell40 \POWERLED.func_state_RNIVO7PG_1_LC_11_5_1  (
            .in0(N__29327),
            .in1(N__26917),
            .in2(N__26885),
            .in3(N__27155),
            .lcout(\POWERLED.func_state_1_m2_1 ),
            .ltout(\POWERLED.func_state_1_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIFFPVI_1_LC_11_5_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFFPVI_1_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFFPVI_1_LC_11_5_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \POWERLED.func_state_RNIFFPVI_1_LC_11_5_2  (
            .in0(N__27061),
            .in1(N__31954),
            .in2(N__26882),
            .in3(N__27082),
            .lcout(\POWERLED.func_state ),
            .ltout(\POWERLED.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_2_LC_11_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_11_5_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_2_LC_11_5_3  (
            .in0(N__30197),
            .in1(_gnd_net_),
            .in2(N__26879),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_426_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_5_4 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_5_4 .LUT_INIT=16'b0011001010001000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_5_4  (
            .in0(N__27944),
            .in1(N__33288),
            .in2(N__29260),
            .in3(N__27416),
            .lcout(\POWERLED.un1_func_state25_6_0_0_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIT3R01_10_LC_11_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIT3R01_10_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIT3R01_10_LC_11_5_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \POWERLED.count_off_RNIT3R01_10_LC_11_5_5  (
            .in0(N__29703),
            .in1(N__29241),
            .in2(N__30798),
            .in3(N__30640),
            .lcout(\POWERLED.N_562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_11_5_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_11_5_6 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.func_state_1_LC_11_5_6  (
            .in0(N__27062),
            .in1(N__31955),
            .in2(N__27086),
            .in3(N__27068),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34398),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_11_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_11_5_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_11_5_7  (
            .in0(N__32668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35444),
            .lcout(N_247),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_11_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_11_6_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_3_LC_11_6_0  (
            .in0(N__27026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28917),
            .lcout(\POWERLED.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34573),
            .ce(N__29389),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_11_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_11_6_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.count_off_4_LC_11_6_1  (
            .in0(N__28916),
            .in1(_gnd_net_),
            .in2(N__27047),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34573),
            .ce(N__29389),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI7K8Q11_4_LC_11_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI7K8Q11_4_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI7K8Q11_4_LC_11_6_2 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.count_off_RNI7K8Q11_4_LC_11_6_2  (
            .in0(N__27053),
            .in1(N__28915),
            .in2(N__29413),
            .in3(N__27043),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI5H7Q11_3_LC_11_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI5H7Q11_3_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI5H7Q11_3_LC_11_6_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.count_off_RNI5H7Q11_3_LC_11_6_3  (
            .in0(N__27032),
            .in1(N__29385),
            .in2(N__28934),
            .in3(N__27025),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(\POWERLED.count_offZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_3_LC_11_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_3_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_3_LC_11_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_3_LC_11_6_4  (
            .in0(N__27001),
            .in1(N__27235),
            .in2(N__27206),
            .in3(N__27202),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_10_LC_11_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_10_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_10_LC_11_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_10_LC_11_6_5  (
            .in0(N__28730),
            .in1(N__27176),
            .in2(N__27164),
            .in3(N__28982),
            .lcout(\POWERLED.count_off_RNI_0Z0Z_10 ),
            .ltout(\POWERLED.count_off_RNI_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI8AQH_10_LC_11_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI8AQH_10_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI8AQH_10_LC_11_6_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \POWERLED.count_off_RNI8AQH_10_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27161),
            .in3(N__29697),
            .lcout(\POWERLED.count_off_RNI8AQHZ0Z_10 ),
            .ltout(\POWERLED.count_off_RNI8AQHZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIU30A4_1_LC_11_6_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIU30A4_1_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIU30A4_1_LC_11_6_7 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \POWERLED.func_state_RNIU30A4_1_LC_11_6_7  (
            .in0(N__30101),
            .in1(_gnd_net_),
            .in2(N__27158),
            .in3(N__29144),
            .lcout(\POWERLED.func_state_1_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_11_7_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_11_7_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_1_LC_11_7_0  (
            .in0(N__33293),
            .in1(N__29240),
            .in2(N__27353),
            .in3(N__30631),
            .lcout(\POWERLED.N_494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIA61DE_10_LC_11_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIA61DE_10_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIA61DE_10_LC_11_7_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.count_clk_RNIA61DE_10_LC_11_7_1  (
            .in0(N__27868),
            .in1(N__35111),
            .in2(N__27943),
            .in3(N__28384),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICU5NF_1_LC_11_7_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICU5NF_1_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICU5NF_1_LC_11_7_2 .LUT_INIT=16'b1101110011101100;
    LogicCell40 \POWERLED.func_state_RNICU5NF_1_LC_11_7_2  (
            .in0(N__33292),
            .in1(N__27275),
            .in2(N__27134),
            .in3(N__27420),
            .lcout(\POWERLED.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_0_LC_11_7_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_0_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_0_LC_11_7_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \POWERLED.func_state_RNI34G9_0_LC_11_7_3  (
            .in0(N__30632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32376),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_i_m2_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIIKO01_LC_11_7_4 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIIKO01_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIIKO01_LC_11_7_4 .LUT_INIT=16'b0001101110111011;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIIKO01_LC_11_7_4  (
            .in0(N__35379),
            .in1(N__27131),
            .in2(N__27119),
            .in3(N__29969),
            .lcout(\POWERLED.N_453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMQ0F_5_LC_11_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMQ0F_5_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMQ0F_5_LC_11_7_5 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \POWERLED.dutycycle_RNIMQ0F_5_LC_11_7_5  (
            .in0(N__31996),
            .in1(N__27682),
            .in2(N__30660),
            .in3(N__31035),
            .lcout(\POWERLED.N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_11_7_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_11_7_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_1_LC_11_7_6  (
            .in0(N__33294),
            .in1(N__27869),
            .in2(N__27422),
            .in3(N__30639),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2O4A1_7_LC_11_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2O4A1_7_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2O4A1_7_LC_11_7_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNI2O4A1_7_LC_11_7_7  (
            .in0(N__27986),
            .in1(N__29189),
            .in2(N__30659),
            .in3(N__27352),
            .lcout(\POWERLED.N_490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_3_LC_11_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_3_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_3_LC_11_8_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_3_LC_11_8_0  (
            .in0(N__31352),
            .in1(N__30070),
            .in2(N__35568),
            .in3(N__32215),
            .lcout(\POWERLED.g1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2MQD_5_LC_11_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2MQD_5_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2MQD_5_LC_11_8_1 .LUT_INIT=16'b0001101100010001;
    LogicCell40 \POWERLED.dutycycle_RNI2MQD_5_LC_11_8_1  (
            .in0(N__31018),
            .in1(N__35377),
            .in2(N__27681),
            .in3(N__30661),
            .lcout(\POWERLED.un1_dutycycle_172_m0_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_0_LC_11_8_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_11_8_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.func_state_RNI2MQD_0_LC_11_8_2  (
            .in0(N__35378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29318),
            .lcout(),
            .ltout(\POWERLED.func_state_RNI2MQDZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIDASB1_6_LC_11_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIDASB1_6_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIDASB1_6_LC_11_8_3 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \POWERLED.dutycycle_RNIDASB1_6_LC_11_8_3  (
            .in0(N__30794),
            .in1(N__27242),
            .in2(N__27257),
            .in3(N__27611),
            .lcout(\POWERLED.dutycycle_eena_13_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_6_LC_11_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_11_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_6_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__33299),
            .in2(_gnd_net_),
            .in3(N__33143),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_8_5 .LUT_INIT=16'b1100010011110100;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_8_5  (
            .in0(N__33300),
            .in1(N__32105),
            .in2(N__32249),
            .in3(N__30283),
            .lcout(\POWERLED.dutycycle_RNI6SKJ1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9S7D5_1_LC_11_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9S7D5_1_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9S7D5_1_LC_11_8_6 .LUT_INIT=16'b0011001101110011;
    LogicCell40 \POWERLED.func_state_RNI9S7D5_1_LC_11_8_6  (
            .in0(N__27532),
            .in1(N__33803),
            .in2(N__27587),
            .in3(N__33402),
            .lcout(\POWERLED.func_state_RNI9S7D5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJ17U4_1_LC_11_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJ17U4_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJ17U4_1_LC_11_8_7 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \POWERLED.func_state_RNIJ17U4_1_LC_11_8_7  (
            .in0(N__33403),
            .in1(N__27533),
            .in2(N__29603),
            .in3(N__33804),
            .lcout(\POWERLED.func_state_RNIJ17U4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILC2B6_4_LC_11_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILC2B6_4_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILC2B6_4_LC_11_9_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_RNILC2B6_4_LC_11_9_0  (
            .in0(N__27490),
            .in1(N__27509),
            .in2(N__33671),
            .in3(N__27500),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNIFPUF_LC_11_9_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNIFPUF_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNIFPUF_LC_11_9_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNIFPUF_LC_11_9_1  (
            .in0(N__27518),
            .in1(N__35118),
            .in2(N__32647),
            .in3(N__27655),
            .lcout(\POWERLED.dutycycle_e_1_4 ),
            .ltout(\POWERLED.dutycycle_e_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_11_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_11_9_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_4_LC_11_9_2  (
            .in0(N__33651),
            .in1(N__27491),
            .in2(N__27503),
            .in3(N__27499),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34741),
            .ce(),
            .sr(N__31567));
    defparam \POWERLED.dutycycle_7_LC_11_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_11_9_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_7_LC_11_9_3  (
            .in0(N__27464),
            .in1(N__27470),
            .in2(N__33670),
            .in3(N__27449),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34741),
            .ce(),
            .sr(N__31567));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_11_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_11_9_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_11_9_4  (
            .in0(N__27656),
            .in1(N__35119),
            .in2(N__32646),
            .in3(N__27479),
            .lcout(\POWERLED.dutycycle_e_1_7 ),
            .ltout(\POWERLED.dutycycle_e_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHG6Q6_7_LC_11_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHG6Q6_7_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHG6Q6_7_LC_11_9_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNIHG6Q6_7_LC_11_9_5  (
            .in0(N__33644),
            .in1(N__27463),
            .in2(N__27452),
            .in3(N__27448),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(\POWERLED.dutycycleZ1Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_3_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_3_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_3_LC_11_9_6 .LUT_INIT=16'b0000010101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_10_3_LC_11_9_6  (
            .in0(N__31340),
            .in1(_gnd_net_),
            .in2(N__27440),
            .in3(N__32192),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_25_0_tz_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_4_LC_11_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_11_9_7 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_4_LC_11_9_7  (
            .in0(N__33142),
            .in1(N__31341),
            .in2(N__27728),
            .in3(N__31808),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2MQD_7_LC_11_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2MQD_7_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2MQD_7_LC_11_10_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \POWERLED.dutycycle_RNI2MQD_7_LC_11_10_0  (
            .in0(N__32773),
            .in1(N__35344),
            .in2(_gnd_net_),
            .in3(N__33298),
            .lcout(\POWERLED.dutycycle_RNI2MQDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_1_LC_11_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_1_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_1_LC_11_10_1 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \POWERLED.func_state_RNI_2_1_LC_11_10_1  (
            .in0(N__33297),
            .in1(N__29263),
            .in2(N__27707),
            .in3(N__30657),
            .lcout(\POWERLED.N_2075_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMQ0F_7_LC_11_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMQ0F_7_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMQ0F_7_LC_11_10_2 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \POWERLED.dutycycle_RNIMQ0F_7_LC_11_10_2  (
            .in0(N__32063),
            .in1(N__32578),
            .in2(N__32821),
            .in3(N__30901),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_1_LC_11_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_1_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_1_LC_11_10_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \POWERLED.func_state_RNI2MQD_1_LC_11_10_3  (
            .in0(N__35345),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33289),
            .lcout(\POWERLED.func_state_RNI2MQDZ0Z_1 ),
            .ltout(\POWERLED.func_state_RNI2MQDZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_8_1_LC_11_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_8_1_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_8_1_LC_11_10_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_8_1_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27617),
            .in3(_gnd_net_),
            .lcout(\POWERLED.func_state_RNI_8Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI_8Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMQ0F_0_1_LC_11_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMQ0F_0_1_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMQ0F_0_1_LC_11_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNIMQ0F_0_1_LC_11_10_5  (
            .in0(N__32579),
            .in1(N__30899),
            .in2(N__27614),
            .in3(N__35541),
            .lcout(\POWERLED.func_state_RNIMQ0F_0Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNIMQ0F_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEBSB1_7_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEBSB1_7_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEBSB1_7_LC_11_10_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.dutycycle_RNIEBSB1_7_LC_11_10_6  (
            .in0(N__27602),
            .in1(_gnd_net_),
            .in2(N__27596),
            .in3(N__27593),
            .lcout(\POWERLED.dutycycle_RNIEBSB1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_11_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_11_10_7 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_11_10_7  (
            .in0(N__27575),
            .in1(N__32062),
            .in2(N__28010),
            .in3(N__27563),
            .lcout(\POWERLED.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3T8L1_0_1_LC_11_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3T8L1_0_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3T8L1_0_1_LC_11_11_0 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \POWERLED.func_state_RNI3T8L1_0_1_LC_11_11_0  (
            .in0(N__30809),
            .in1(N__28073),
            .in2(N__32407),
            .in3(N__28066),
            .lcout(\POWERLED.count_clk_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_11_11_1 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_11_11_1 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_11_11_1  (
            .in0(N__35325),
            .in1(N__32524),
            .in2(_gnd_net_),
            .in3(N__35142),
            .lcout(\POWERLED.N_443 ),
            .ltout(\POWERLED.N_443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIH37EG_1_LC_11_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIH37EG_1_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIH37EG_1_LC_11_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_RNIH37EG_1_LC_11_11_2  (
            .in0(N__27998),
            .in1(N__27821),
            .in2(N__27989),
            .in3(N__27902),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIS94QD_1_LC_11_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIS94QD_1_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIS94QD_1_LC_11_11_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \POWERLED.func_state_RNIS94QD_1_LC_11_11_4  (
            .in0(N__27891),
            .in1(N__33290),
            .in2(N__27981),
            .in3(N__27927),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_LC_11_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_11_11_5 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_LC_11_11_5  (
            .in0(N__33291),
            .in1(N__27890),
            .in2(N__35551),
            .in3(N__29264),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI02AS_6_LC_11_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI02AS_6_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI02AS_6_LC_11_11_6 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \POWERLED.count_clk_RNI02AS_6_LC_11_11_6  (
            .in0(N__32523),
            .in1(N__27815),
            .in2(_gnd_net_),
            .in3(N__35533),
            .lcout(\POWERLED.N_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_10_LC_11_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_10_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_10_LC_11_12_0 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_10_LC_11_12_0  (
            .in0(N__35340),
            .in1(N__35207),
            .in2(N__30296),
            .in3(N__28303),
            .lcout(),
            .ltout(\POWERLED.N_506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_0_10_LC_11_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_0_10_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_0_10_LC_11_12_1 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_0_10_LC_11_12_1  (
            .in0(N__28302),
            .in1(_gnd_net_),
            .in2(N__27758),
            .in3(N__33301),
            .lcout(\POWERLED.dutycycle_RNI6SKJ1_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_3_LC_11_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_11_12_2 .LUT_INIT=16'b0001111100111111;
    LogicCell40 \POWERLED.dutycycle_RNI_9_3_LC_11_12_2  (
            .in0(N__32228),
            .in1(N__31387),
            .in2(N__33146),
            .in3(N__32813),
            .lcout(\POWERLED.g0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_11_LC_11_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_11_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_11_LC_11_12_3 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_11_LC_11_12_3  (
            .in0(N__28201),
            .in1(N__31869),
            .in2(N__32026),
            .in3(N__32085),
            .lcout(),
            .ltout(\POWERLED.N_514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHDMC5_11_LC_11_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHDMC5_11_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHDMC5_11_LC_11_12_4 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \POWERLED.dutycycle_RNIHDMC5_11_LC_11_12_4  (
            .in0(N__33819),
            .in1(N__28103),
            .in2(N__28328),
            .in3(N__33435),
            .lcout(\POWERLED.dutycycle_RNIHDMC5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_10_LC_11_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_10_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_10_LC_11_12_5 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_10_LC_11_12_5  (
            .in0(N__28304),
            .in1(N__31868),
            .in2(N__32025),
            .in3(N__32084),
            .lcout(\POWERLED.N_508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_11_LC_11_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_11_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_11_LC_11_12_6 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_11_LC_11_12_6  (
            .in0(N__30295),
            .in1(N__28200),
            .in2(N__35390),
            .in3(N__35208),
            .lcout(),
            .ltout(\POWERLED.N_512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_0_11_LC_11_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_0_11_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_0_11_LC_11_12_7 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_0_11_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__33302),
            .in2(N__28205),
            .in3(N__28199),
            .lcout(\POWERLED.dutycycle_RNI6SKJ1_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3T8L1_14_LC_11_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3T8L1_14_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3T8L1_14_LC_11_13_0 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \POWERLED.dutycycle_RNI3T8L1_14_LC_11_13_0  (
            .in0(N__33295),
            .in1(N__34886),
            .in2(N__34968),
            .in3(N__33434),
            .lcout(\POWERLED.un1_clk_100khz_47_and_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_14_LC_11_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_14_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_14_LC_11_13_1 .LUT_INIT=16'b0111000000110000;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_14_LC_11_13_1  (
            .in0(N__34959),
            .in1(N__31886),
            .in2(N__32093),
            .in3(N__32014),
            .lcout(),
            .ltout(\POWERLED.N_526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQ8KL5_14_LC_11_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQ8KL5_14_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQ8KL5_14_LC_11_13_2 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \POWERLED.dutycycle_RNIQ8KL5_14_LC_11_13_2  (
            .in0(N__33666),
            .in1(N__33821),
            .in2(N__28097),
            .in3(N__28094),
            .lcout(\POWERLED.dutycycle_en_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE3861_12_LC_11_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE3861_12_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE3861_12_LC_11_13_3 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \POWERLED.dutycycle_RNIE3861_12_LC_11_13_3  (
            .in0(N__28527),
            .in1(N__35324),
            .in2(N__35148),
            .in3(N__35209),
            .lcout(),
            .ltout(\POWERLED.N_518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE3861_0_12_LC_11_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE3861_0_12_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE3861_0_12_LC_11_13_4 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \POWERLED.dutycycle_RNIE3861_0_12_LC_11_13_4  (
            .in0(N__33296),
            .in1(_gnd_net_),
            .in2(N__28532),
            .in3(N__28526),
            .lcout(\POWERLED.dutycycle_RNIE3861_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_12_LC_11_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_12_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_12_LC_11_13_5 .LUT_INIT=16'b0111000000110000;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_12_LC_11_13_5  (
            .in0(N__28528),
            .in1(N__31885),
            .in2(N__32092),
            .in3(N__32013),
            .lcout(),
            .ltout(\POWERLED.N_520_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIPK9V4_12_LC_11_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIPK9V4_12_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIPK9V4_12_LC_11_13_6 .LUT_INIT=16'b0011001100111011;
    LogicCell40 \POWERLED.dutycycle_RNIPK9V4_12_LC_11_13_6  (
            .in0(N__28445),
            .in1(N__33820),
            .in2(N__28439),
            .in3(N__33433),
            .lcout(\POWERLED.dutycycle_RNIPK9V4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIB15N11_15_LC_11_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIB15N11_15_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIB15N11_15_LC_11_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIB15N11_15_LC_11_13_7  (
            .in0(N__29458),
            .in1(N__28403),
            .in2(_gnd_net_),
            .in3(N__28420),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_11_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_11_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_15_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28421),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34720),
            .ce(N__29459),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIUQMRH_1_LC_11_15_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIUQMRH_1_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIUQMRH_1_LC_11_15_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \POWERLED.func_state_RNIUQMRH_1_LC_11_15_4  (
            .in0(N__32528),
            .in1(N__35272),
            .in2(N__28397),
            .in3(N__28373),
            .lcout(\POWERLED.func_state_RNIUQMRH_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI0KOA4_11_LC_11_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI0KOA4_11_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI0KOA4_11_LC_11_16_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.count_clk_RNI0KOA4_11_LC_11_16_0  (
            .in0(N__34783),
            .in1(N__28348),
            .in2(N__28337),
            .in3(N__33983),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_11_16_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_11_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_clk_11_LC_11_16_1  (
            .in0(N__28349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34784),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34739),
            .ce(N__33996),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_16_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_16_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__34865),
            .in2(_gnd_net_),
            .in3(N__34786),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI92UF4_0_LC_11_16_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI92UF4_0_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI92UF4_0_LC_11_16_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNI92UF4_0_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__34754),
            .in2(N__28685),
            .in3(N__33982),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(\POWERLED.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_11_16_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_11_16_5 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__28665),
            .in2(N__28682),
            .in3(N__34782),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIA3UF4_1_LC_11_16_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIA3UF4_1_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIA3UF4_1_LC_11_16_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIA3UF4_1_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__28646),
            .in2(N__28679),
            .in3(N__33984),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(\POWERLED.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_11_16_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_11_16_7 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_clk_1_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__34864),
            .in2(N__28649),
            .in3(N__34785),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34739),
            .ce(N__33996),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_12_2_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_12_2_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_12_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_11_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28715),
            .lcout(\POWERLED.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__29411),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_12_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_12_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_13_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29057),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__29411),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_12_2_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_12_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_14_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28640),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__29411),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_12_2_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_12_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_7_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28603),
            .lcout(\POWERLED.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__29411),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_12_2_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_12_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_8_LC_12_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28564),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__29411),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_12_3_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_12_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_6_LC_12_3_0  (
            .in0(N__28781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34583),
            .ce(N__29452),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI3E6Q11_2_LC_12_3_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI3E6Q11_2_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI3E6Q11_2_LC_12_3_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \POWERLED.count_off_RNI3E6Q11_2_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__28808),
            .in2(N__29435),
            .in3(N__28816),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_12_3_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_12_3_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_2_LC_12_3_2  (
            .in0(N__28817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34583),
            .ce(N__29452),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI9N9Q11_5_LC_12_3_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI9N9Q11_5_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI9N9Q11_5_LC_12_3_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNI9N9Q11_5_LC_12_3_3  (
            .in0(N__29406),
            .in1(N__28793),
            .in2(_gnd_net_),
            .in3(N__28801),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_12_3_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_12_3_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_5_LC_12_3_4  (
            .in0(N__28802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34583),
            .ce(N__29452),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIBQAQ11_6_LC_12_3_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBQAQ11_6_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBQAQ11_6_LC_12_3_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIBQAQ11_6_LC_12_3_5  (
            .in0(N__29407),
            .in1(N__28787),
            .in2(_gnd_net_),
            .in3(N__28780),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(\POWERLED.count_offZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_1_LC_12_3_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_1_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_1_LC_12_3_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_off_RNI_0_1_LC_12_3_6  (
            .in0(N__28762),
            .in1(N__28747),
            .in2(N__28733),
            .in3(N__28833),
            .lcout(\POWERLED.un34_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI3L0N11_11_LC_12_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI3L0N11_11_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI3L0N11_11_LC_12_3_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \POWERLED.count_off_RNI3L0N11_11_LC_12_3_7  (
            .in0(N__28721),
            .in1(_gnd_net_),
            .in2(N__29436),
            .in3(N__28711),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_12_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_12_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_1_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(N__28940),
            .in2(_gnd_net_),
            .in3(N__28920),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34532),
            .ce(N__29369),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI7R2N11_13_LC_12_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI7R2N11_13_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI7R2N11_13_LC_12_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNI7R2N11_13_LC_12_4_1  (
            .in0(N__29402),
            .in1(N__29066),
            .in2(_gnd_net_),
            .in3(N__29053),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(\POWERLED.count_offZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_12_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_12_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_12_4_2  (
            .in0(N__28961),
            .in1(N__29032),
            .in2(N__29012),
            .in3(N__29008),
            .lcout(\POWERLED.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_12_4_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_12_4_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_off_0_LC_12_4_3  (
            .in0(N__28919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28962),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34532),
            .ce(N__29369),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNICU5NF_0_LC_12_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNICU5NF_0_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNICU5NF_0_LC_12_4_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_off_RNICU5NF_0_LC_12_4_4  (
            .in0(N__28963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28918),
            .lcout(),
            .ltout(\POWERLED.count_off_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIA46B11_0_LC_12_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIA46B11_0_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIA46B11_0_LC_12_4_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNIA46B11_0_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(N__28973),
            .in2(N__28967),
            .in3(N__29368),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(\POWERLED.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_12_4_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_12_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28943),
            .in3(N__28837),
            .lcout(\POWERLED.count_off_RNIZ0Z_1 ),
            .ltout(\POWERLED.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIB56B11_1_LC_12_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIB56B11_1_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIB56B11_1_LC_12_4_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \POWERLED.count_off_RNIB56B11_1_LC_12_4_7  (
            .in0(N__28921),
            .in1(N__28847),
            .in2(N__28841),
            .in3(N__29367),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_0_LC_12_5_0 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_0_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_0_LC_12_5_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_0_LC_12_5_0  (
            .in0(N__35447),
            .in1(N__32307),
            .in2(_gnd_net_),
            .in3(N__30616),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_0_a6_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_12_5_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_12_5_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_12_5_1  (
            .in0(N__31987),
            .in1(N__33280),
            .in2(N__29594),
            .in3(N__29246),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_o_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_12_5_2 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_12_5_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_12_5_2  (
            .in0(N__29591),
            .in1(N__29582),
            .in2(N__29576),
            .in3(N__29138),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI31IBH_0_LC_12_5_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI31IBH_0_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI31IBH_0_LC_12_5_3 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \POWERLED.func_state_RNI31IBH_0_LC_12_5_3  (
            .in0(N__29573),
            .in1(N__29310),
            .in2(N__29465),
            .in3(N__33668),
            .lcout(\POWERLED.func_state_RNI31IBHZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIGCDO1_1_LC_12_5_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIGCDO1_1_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIGCDO1_1_LC_12_5_4 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \POWERLED.func_state_RNIGCDO1_1_LC_12_5_4  (
            .in0(N__35446),
            .in1(N__32670),
            .in2(N__29273),
            .in3(N__29187),
            .lcout(\POWERLED.N_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_LC_12_5_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_12_5_5 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_LC_12_5_5  (
            .in0(N__32669),
            .in1(N__35445),
            .in2(N__35135),
            .in3(N__29309),
            .lcout(\POWERLED.func_state_RNIBVNSZ0Z_0 ),
            .ltout(\POWERLED.func_state_RNIBVNSZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBQDR2_1_LC_12_5_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBQDR2_1_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBQDR2_1_LC_12_5_6 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \POWERLED.func_state_RNIBQDR2_1_LC_12_5_6  (
            .in0(N__29245),
            .in1(N__29188),
            .in2(N__29147),
            .in3(N__33794),
            .lcout(\POWERLED.func_state_1_m0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_12_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_12_5_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_12_5_7  (
            .in0(N__32308),
            .in1(N__35448),
            .in2(N__32680),
            .in3(N__35110),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_12_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_12_6_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__35561),
            .in2(_gnd_net_),
            .in3(N__32244),
            .lcout(\POWERLED.G_11_i_o10_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_1_LC_12_6_3 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_1_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_1_LC_12_6_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \VCCIN_PWRGD.un10_output_1_LC_12_6_3  (
            .in0(N__30796),
            .in1(N__29132),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\VCCIN_PWRGD.un10_outputZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_12_6_4 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_12_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_12_6_4  (
            .in0(N__29765),
            .in1(N__29759),
            .in2(N__29747),
            .in3(N__29744),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_0_o2_2_LC_12_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_0_o2_2_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_0_o2_2_LC_12_6_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_0_o2_2_LC_12_6_7  (
            .in0(N__32375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29968),
            .lcout(\POWERLED.N_253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMQ0F_4_LC_12_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMQ0F_4_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMQ0F_4_LC_12_7_0 .LUT_INIT=16'b0001001110110011;
    LogicCell40 \POWERLED.dutycycle_RNIMQ0F_4_LC_12_7_0  (
            .in0(N__32652),
            .in1(N__31411),
            .in2(N__30905),
            .in3(N__35557),
            .lcout(\POWERLED.dutycycle_e_N_6L11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_1_LC_12_7_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_1_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_1_LC_12_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_6_1_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29995),
            .lcout(\POWERLED.func_state_RNI_6Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI_6Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_18_0_LC_12_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_18_0_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_18_0_LC_12_7_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.dutycycle_RNI_18_0_LC_12_7_2  (
            .in0(N__29645),
            .in1(_gnd_net_),
            .in2(N__29630),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.N_2361_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIR8072_5_LC_12_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIR8072_5_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIR8072_5_LC_12_7_3 .LUT_INIT=16'b0011000000110101;
    LogicCell40 \POWERLED.dutycycle_RNIR8072_5_LC_12_7_3  (
            .in0(N__31046),
            .in1(N__30082),
            .in2(N__29627),
            .in3(N__30107),
            .lcout(N_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2MQD_4_LC_12_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2MQD_4_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2MQD_4_LC_12_7_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \POWERLED.dutycycle_RNI2MQD_4_LC_12_7_4  (
            .in0(N__35457),
            .in1(N__31412),
            .in2(_gnd_net_),
            .in3(N__33345),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI2MQDZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOGRS_4_LC_12_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOGRS_4_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOGRS_4_LC_12_7_5 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \POWERLED.dutycycle_RNIOGRS_4_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__29612),
            .in2(N__29606),
            .in3(N__32082),
            .lcout(\POWERLED.dutycycle_RNIOGRSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_12_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_12_7_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_12_7_6  (
            .in0(N__30069),
            .in1(N__31413),
            .in2(N__30434),
            .in3(N__30425),
            .lcout(N_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3O4A1_2_LC_12_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3O4A1_2_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3O4A1_2_LC_12_7_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.dutycycle_RNI3O4A1_2_LC_12_7_7  (
            .in0(N__32651),
            .in1(N__30289),
            .in2(N__35476),
            .in3(N__30196),
            .lcout(\POWERLED.N_488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_12_8_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_12_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_0_LC_12_8_1  (
            .in0(N__32649),
            .in1(N__35127),
            .in2(N__35475),
            .in3(N__30662),
            .lcout(\POWERLED.N_540_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOGRS_5_LC_12_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOGRS_5_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOGRS_5_LC_12_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.dutycycle_RNIOGRS_5_LC_12_8_2  (
            .in0(N__31020),
            .in1(N__29975),
            .in2(_gnd_net_),
            .in3(N__30900),
            .lcout(POWERLED_un1_dutycycle_172_m0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_1_LC_12_8_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_1_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_1_LC_12_8_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.func_state_RNI_4_1_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__30071),
            .in2(_gnd_net_),
            .in3(N__35540),
            .lcout(\POWERLED.func_state_RNI_4Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI_4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5DLR_5_LC_12_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5DLR_5_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5DLR_5_LC_12_8_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.dutycycle_RNI5DLR_5_LC_12_8_4  (
            .in0(N__31019),
            .in1(N__29984),
            .in2(N__29978),
            .in3(N__32648),
            .lcout(\POWERLED.dutycycle_RNI5DLRZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI7ABC3_5_LC_12_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI7ABC3_5_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI7ABC3_5_LC_12_8_5 .LUT_INIT=16'b1011111100111111;
    LogicCell40 \POWERLED.dutycycle_RNI7ABC3_5_LC_12_8_5  (
            .in0(N__31052),
            .in1(N__29958),
            .in2(N__29894),
            .in3(N__33793),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI7ABC3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITNMH4_5_LC_12_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITNMH4_5_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITNMH4_5_LC_12_8_6 .LUT_INIT=16'b0111010011111100;
    LogicCell40 \POWERLED.dutycycle_RNITNMH4_5_LC_12_8_6  (
            .in0(N__29959),
            .in1(N__30795),
            .in2(N__29897),
            .in3(N__29893),
            .lcout(\POWERLED.g2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_12_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_12_8_7 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_12_8_7  (
            .in0(N__32650),
            .in1(N__32377),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6RAN_5_LC_12_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6RAN_5_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6RAN_5_LC_12_9_0 .LUT_INIT=16'b1100111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI6RAN_5_LC_12_9_0  (
            .in0(N__30663),
            .in1(N__35175),
            .in2(N__33377),
            .in3(N__31044),
            .lcout(\POWERLED.g1_1cf0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_12_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_12_9_1 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_12_9_1  (
            .in0(N__32208),
            .in1(N__31347),
            .in2(_gnd_net_),
            .in3(N__32772),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_5_LC_12_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_12_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_5_LC_12_9_2  (
            .in0(N__31348),
            .in1(N__31045),
            .in2(N__30929),
            .in3(N__31259),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6RAN_1_LC_12_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6RAN_1_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6RAN_1_LC_12_9_3 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \POWERLED.func_state_RNI6RAN_1_LC_12_9_3  (
            .in0(N__35176),
            .in1(N__33372),
            .in2(N__30664),
            .in3(N__30465),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_32_and_i_0cf0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRKB61_0_1_LC_12_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRKB61_0_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRKB61_0_1_LC_12_9_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.func_state_RNIRKB61_0_1_LC_12_9_4  (
            .in0(N__30466),
            .in1(N__35403),
            .in2(N__30908),
            .in3(N__30898),
            .lcout(\POWERLED.un1_clk_100khz_32_and_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNILP0F_1_LC_12_9_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNILP0F_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNILP0F_1_LC_12_9_5 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \POWERLED.func_state_RNILP0F_1_LC_12_9_5  (
            .in0(N__33376),
            .in1(N__30790),
            .in2(N__30665),
            .in3(N__30467),
            .lcout(\POWERLED.func_state_RNILP0FZ0Z_1 ),
            .ltout(\POWERLED.func_state_RNILP0FZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHDMC5_3_LC_12_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHDMC5_3_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHDMC5_3_LC_12_9_6 .LUT_INIT=16'b0000010011111111;
    LogicCell40 \POWERLED.dutycycle_RNIHDMC5_3_LC_12_9_6  (
            .in0(N__30440),
            .in1(N__30449),
            .in2(N__30443),
            .in3(N__33789),
            .lcout(\POWERLED.dutycycle_RNIHDMC5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_3_LC_12_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_3_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_3_LC_12_9_7 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_3_LC_12_9_7  (
            .in0(N__31997),
            .in1(N__31891),
            .in2(N__32248),
            .in3(N__32081),
            .lcout(\POWERLED.N_523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8CJA6_3_LC_12_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8CJA6_3_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8CJA6_3_LC_12_10_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \POWERLED.dutycycle_RNI8CJA6_3_LC_12_10_0  (
            .in0(N__31618),
            .in1(N__31627),
            .in2(N__31601),
            .in3(N__33662),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(\POWERLED.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_3_LC_12_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_12_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_3_LC_12_10_1  (
            .in0(N__31812),
            .in1(N__32769),
            .in2(N__31631),
            .in3(N__31255),
            .lcout(\POWERLED.N_12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_12_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_12_10_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_3_LC_12_10_2  (
            .in0(N__31600),
            .in1(N__31628),
            .in2(N__33674),
            .in3(N__31619),
            .lcout(\POWERLED.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34719),
            .ce(),
            .sr(N__31581));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__32193),
            .in2(_gnd_net_),
            .in3(N__31256),
            .lcout(),
            .ltout(\POWERLED.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_6_LC_12_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_12_10_4 .LUT_INIT=16'b0000010100111111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_6_LC_12_10_4  (
            .in0(N__32771),
            .in1(N__33115),
            .in2(N__31439),
            .in3(N__31813),
            .lcout(),
            .ltout(\POWERLED.g0_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_4_LC_12_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_4_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_4_LC_12_10_5 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \POWERLED.dutycycle_RNI_2_4_LC_12_10_5  (
            .in0(N__31346),
            .in1(N__31436),
            .in2(N__31430),
            .in3(N__32900),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_3_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_3_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_3_LC_12_10_7 .LUT_INIT=16'b0001010101010111;
    LogicCell40 \POWERLED.dutycycle_RNI_12_3_LC_12_10_7  (
            .in0(N__31345),
            .in1(N__32770),
            .in2(N__32237),
            .in3(N__31257),
            .lcout(\POWERLED.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE3861_15_LC_12_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE3861_15_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE3861_15_LC_12_11_0 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \POWERLED.dutycycle_RNIE3861_15_LC_12_11_0  (
            .in0(N__31106),
            .in1(N__35458),
            .in2(N__35206),
            .in3(N__35143),
            .lcout(\POWERLED.N_527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_12_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_12_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31105),
            .lcout(\POWERLED.N_2341_i ),
            .ltout(\POWERLED.N_2341_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_15_LC_12_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_15_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_15_LC_12_11_2 .LUT_INIT=16'b1010001000100010;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_15_LC_12_11_2  (
            .in0(N__32064),
            .in1(N__31864),
            .in2(N__33824),
            .in3(N__32007),
            .lcout(),
            .ltout(\POWERLED.N_529_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQ8KL5_1_LC_12_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQ8KL5_1_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQ8KL5_1_LC_12_11_3 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \POWERLED.func_state_RNIQ8KL5_1_LC_12_11_3  (
            .in0(N__33152),
            .in1(N__33811),
            .in2(N__33677),
            .in3(N__33667),
            .lcout(\POWERLED.dutycycle_en_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3T8L1_1_LC_12_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3T8L1_1_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3T8L1_1_LC_12_11_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \POWERLED.func_state_RNI3T8L1_1_LC_12_11_4  (
            .in0(N__33432),
            .in1(N__33370),
            .in2(N__33182),
            .in3(N__33169),
            .lcout(\POWERLED.un1_clk_100khz_48_and_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_LC_12_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_LC_12_11_6 .LUT_INIT=16'b1010100011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_LC_12_11_6  (
            .in0(N__33141),
            .in1(N__32814),
            .in2(N__31825),
            .in3(N__32953),
            .lcout(\POWERLED.g0_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_12_11_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_12_11_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_12_11_7  (
            .in0(N__32008),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32894),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_3_LC_12_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_3_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_3_LC_12_12_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_8_3_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__32229),
            .in2(_gnd_net_),
            .in3(N__32812),
            .lcout(\POWERLED.G_7_i_o5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8H551_3_LC_12_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8H551_3_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8H551_3_LC_12_12_4 .LUT_INIT=16'b0011101100110011;
    LogicCell40 \POWERLED.dutycycle_RNI8H551_3_LC_12_12_4  (
            .in0(N__32645),
            .in1(N__35409),
            .in2(N__32406),
            .in3(N__32230),
            .lcout(\POWERLED.dutycycle_e_N_3L4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMSAB1_9_LC_12_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMSAB1_9_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMSAB1_9_LC_12_12_6 .LUT_INIT=16'b0000101010001010;
    LogicCell40 \POWERLED.dutycycle_RNIMSAB1_9_LC_12_12_6  (
            .in0(N__32083),
            .in1(N__32012),
            .in2(N__31884),
            .in3(N__31824),
            .lcout(\POWERLED.N_505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_6_LC_12_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_6_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_6_LC_12_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.count_clk_RNI_6_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35629),
            .lcout(\POWERLED.N_412_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE3861_14_LC_12_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE3861_14_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE3861_14_LC_12_13_1 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIE3861_14_LC_12_13_1  (
            .in0(N__35351),
            .in1(N__35194),
            .in2(N__35153),
            .in3(N__34960),
            .lcout(\POWERLED.N_524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_12_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_12_14_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_clk_0_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__34872),
            .in2(_gnd_net_),
            .in3(N__34808),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34716),
            .ce(N__34003),
            .sr(_gnd_net_));
endmodule // TOP
