-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Aug 9 2022 16:48:19

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__18893\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PCH_PWROK_c\ : std_logic;
signal \PCH_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \PCH_PWRGD.un4_count_11\ : std_logic;
signal \PCH_PWRGD.un4_count_8\ : std_logic;
signal \PCH_PWRGD.un4_count_10\ : std_logic;
signal \POWERLED.count_i_0_0\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \POWERLED.count_i_1\ : std_logic;
signal \POWERLED.un1_count_2_cry_0\ : std_logic;
signal \POWERLED.un1_count_2_2\ : std_logic;
signal \POWERLED.count_i_2\ : std_logic;
signal \POWERLED.un1_count_2_cry_1\ : std_logic;
signal \POWERLED.count_i_3\ : std_logic;
signal \POWERLED.un1_count_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_2_4\ : std_logic;
signal \POWERLED.count_i_4\ : std_logic;
signal \POWERLED.un1_count_2_cry_3\ : std_logic;
signal \POWERLED.count_i_5\ : std_logic;
signal \POWERLED.un1_count_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_2_6\ : std_logic;
signal \POWERLED.count_i_6\ : std_logic;
signal \POWERLED.un1_count_2_cry_5\ : std_logic;
signal \POWERLED.count_i_7\ : std_logic;
signal \POWERLED.un1_count_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_2_cry_7\ : std_logic;
signal \POWERLED.count_i_8\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \POWERLED.un1_count_2_9\ : std_logic;
signal \POWERLED.count_i_9\ : std_logic;
signal \POWERLED.un1_count_2_cry_8\ : std_logic;
signal \POWERLED.count_i_10\ : std_logic;
signal \POWERLED.un1_count_2_cry_9\ : std_logic;
signal \POWERLED.count_i_11\ : std_logic;
signal \POWERLED.un1_count_2_cry_10\ : std_logic;
signal \POWERLED.un1_count_2_12\ : std_logic;
signal \POWERLED.count_i_12\ : std_logic;
signal \POWERLED.un1_count_2_cry_11\ : std_logic;
signal \POWERLED.count_i_13\ : std_logic;
signal \POWERLED.un1_count_2_cry_12\ : std_logic;
signal \POWERLED.count_i_14\ : std_logic;
signal \POWERLED.un1_count_2_cry_13\ : std_logic;
signal \POWERLED.count_i_15\ : std_logic;
signal \POWERLED.un1_count_2_cry_14\ : std_logic;
signal \POWERLED.un1_count_2_cry_15\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \VCCST_EN_c_i\ : std_logic;
signal \POWERLED.un1_countlto15_5_cascade_\ : std_logic;
signal \POWERLED.un1_countlto15_4_cascade_\ : std_logic;
signal \POWERLED.un1_countlto15_7\ : std_logic;
signal \POWERLED.count_RNIOVT24Z0Z_11\ : std_logic;
signal \POWERLED.count_RNIOVT24Z0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_countlt6\ : std_logic;
signal \VPP_OK_c\ : std_logic;
signal \VDDQ_EN_c\ : std_logic;
signal \PCH_PWRGD.curr_state_RNICTB05Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_3_i\ : std_logic;
signal \PCH_PWRGD.N_3_i_cascade_\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.un1_curr_state_0_sqmuxa_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \VR_READY_VCCIN_c\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.un1_curr_state10_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.N_39_4\ : std_logic;
signal \PCH_PWRGD.curr_state_RNICTB05Z0Z_0\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_386\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un1_count_2_0\ : std_logic;
signal \POWERLED.un1_count_2_5\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7_cascade_\ : std_logic;
signal \POWERLED.un1_count_2_1\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.g0_0_4\ : std_logic;
signal \POWERLED.g0_0_7_cascade_\ : std_logic;
signal \POWERLED.un1_countlt6_0\ : std_logic;
signal \POWERLED.g0_0_5\ : std_logic;
signal \tmp_RNIRH3P\ : std_logic;
signal \POWERLED.un1_count_2_cry_15_THRU_CO\ : std_logic;
signal \tmp_RNIRH3P_cascade_\ : std_logic;
signal \POWERLED.un1_count_0\ : std_logic;
signal \COUNTER.tmp_i\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \PWRBTN_LED_c\ : std_logic;
signal \POWERLED.pwm_out_RNOZ0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_1_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_1_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_1_cry_3\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_1_cry_4\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_1_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_1_cry_6\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.un1_count_1_cry_7\ : std_logic;
signal \POWERLED.un1_count_1_cry_8\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_1_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_1_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_1_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_1_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_39_6\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \POWERLED.un1_count_2_11\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un1_count_2_3\ : std_logic;
signal \POWERLED.un1_count_2_15\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.curr_state_RNI75RB5Z0Z_0\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER.un4_counter_7\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.un4_counter_7_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \VPP_VDDQ.N_39_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.un1_count_2_14\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.un1_count_2_13\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \VPP_VDDQ.G_110_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_RNIQINR7Z0Z_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8_cascade_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un6_count_11_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_8\ : std_logic;
signal \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \POWERLED.un1_count_2_10\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.un1_count_2_8\ : std_logic;
signal \POWERLED.func_state_RNI9L40BZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.un1_count_2_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \VPP_VDDQ.N_32_i\ : std_logic;
signal \POWERLED.count_off_0_sqmuxa\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un4_count_8_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_1_i\ : std_logic;
signal \RSMRST_PWRGD.N_1_i_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_85\ : std_logic;
signal \RSMRST_PWRGD.N_85_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.un4_count_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.un4_count_9\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.N_51_i\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un4_count_11\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0\ : std_logic;
signal \RSMRST_PWRGD.N_39_3\ : std_logic;
signal \V5A_EN_c\ : std_logic;
signal \V5A_OK_c\ : std_logic;
signal \V33A_OK_c\ : std_logic;
signal \V1P8A_OK_c\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_7_l_fx\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_0\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_1\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_0\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_1\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_9\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_10\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_15\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ_un2_vpp_en_0_i\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_i_29\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_axb_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_i_28\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \POWERLED.dutycycle_1_sqmuxa_i_o6_0_0_cascade_\ : std_logic;
signal \POWERLED.N_68_i\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_0\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_1\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_2\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_5\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_7\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_8\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_9\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_10\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_11\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_12\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.N_39_0\ : std_logic;
signal \POWERLED.func_state_RNI9L40BZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIQAI81Z0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNIOQLJZ0Z_4\ : std_logic;
signal \POWERLED.dutycycle_fastZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fast_RNILMLMZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIJL1R1Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNIC8C11Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNIO18NZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNIO18NZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIQ09G1Z0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNIB1FLZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI84C11Z0Z_14\ : std_logic;
signal \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNIJNBA1Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNIE4FLZ0Z_9\ : std_logic;
signal \POWERLED.N_165\ : std_logic;
signal \POWERLED.dutycycle_RNI2V0PZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI712I1Z0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_1_44_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIF3561Z0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI53MGZ0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNI31MGZ0Z_12\ : std_logic;
signal \POWERLED.dutycycle_RNI73C11Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNI31MG_0Z0Z_12\ : std_logic;
signal \POWERLED.dutycycle_RNI75MGZ0Z_15\ : std_logic;
signal \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa\ : std_logic;
signal \VCCIN_EN_c\ : std_logic;
signal \ALL_SYS_PWRGD.N_44_cascade_\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_5\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_3\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_11\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_2\ : std_logic;
signal \ALL_SYS_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \ALL_SYS_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.un1_curr_state10_0\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_9\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_1\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_10\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_10\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \ALL_SYS_PWRGD.N_1_i\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_7\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_6\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_8\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_4\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_8\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_14\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_13\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_15\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_12\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_11\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o2_10_1\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o2_9_1\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o2_8_1\ : std_logic;
signal \POWERLED.un1_func_state11_2_i_o6_0_2\ : std_logic;
signal \POWERLED.N_100_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_sqmuxa_i_o6_1_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_sqmuxa_i_o6_1_6\ : std_logic;
signal \ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.N_39_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_7\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_11\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \POWERLED.dutycycle_s_0\ : std_logic;
signal \POWERLED.dutycycle_cry_c_0_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_s_1\ : std_logic;
signal \POWERLED.dutycycle_cry_0\ : std_logic;
signal \POWERLED.dutycycle_cry_1\ : std_logic;
signal \POWERLED.dutycycle_cry_2\ : std_logic;
signal \POWERLED.dutycycle_cry_3\ : std_logic;
signal \POWERLED.dutycycle_cry_4\ : std_logic;
signal \POWERLED.dutycycle_cry_5\ : std_logic;
signal \POWERLED.dutycycle_cry_6\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \POWERLED.dutycycle_cry_7\ : std_logic;
signal \POWERLED.dutycycle_cry_8\ : std_logic;
signal \POWERLED.dutycycle_cry_9\ : std_logic;
signal \POWERLED.dutycycle_cry_10\ : std_logic;
signal \POWERLED.dutycycle_cry_11\ : std_logic;
signal \POWERLED.dutycycle_cry_12\ : std_logic;
signal \POWERLED.dutycycle_cry_13\ : std_logic;
signal \POWERLED.dutycycle_cry_14\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o3_5_0_cascade_\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o3_6_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o3_7_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.un1_dutycycle_1_39_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI34C41Z0Z_8\ : std_logic;
signal \POWERLED.N_78\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.func_state_ns_0_i_o2_11_1\ : std_logic;
signal \POWERLED.dutycycle_RNIFHLJZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI16B71Z0Z_5\ : std_logic;
signal \POWERLED.N_126\ : std_logic;
signal \POWERLED.N_168_cascade_\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_2_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNI95RKLZ0Z_8\ : std_logic;
signal \POWERLED.count_clk_RNI95RKLZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.N_39_1\ : std_logic;
signal \POWERLED.N_167\ : std_logic;
signal \POWERLED.dutycycle_s_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI6NI81Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIK4I81Z0Z_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNIEJ021Z0Z_4\ : std_logic;
signal \POWERLED.N_173_cascade_\ : std_logic;
signal \POWERLED.N_84_cascade_\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.N_119\ : std_logic;
signal \POWERLED.N_65_i\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.N_84\ : std_logic;
signal \POWERLED.N_116\ : std_logic;
signal \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_2\ : std_logic;
signal \POWERLED.N_197\ : std_logic;
signal \POWERLED.dutycycle_cnst_1_i_o2_0_a3_2_5\ : std_logic;
signal \POWERLED.N_196_cascade_\ : std_logic;
signal \POWERLED.N_115\ : std_logic;
signal \POWERLED.N_92\ : std_logic;
signal \POWERLED.N_120_cascade_\ : std_logic;
signal \POWERLED.N_100\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_0_0\ : std_logic;
signal \POWERLED.N_171_cascade_\ : std_logic;
signal \POWERLED.N_163\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_i\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal \V33S_OK_c\ : std_logic;
signal \VCCST_CPU_OK_c\ : std_logic;
signal \ALL_SYS_PWRGD.N_194\ : std_logic;
signal \V5S_OK_c\ : std_logic;
signal \ALL_SYS_PWRGD.m4_0_0_a3_1\ : std_logic;
signal \POWERLED.dutycycle_s_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.un1_dutycycle_4_sqmuxa_0\ : std_logic;
signal \POWERLED.dutycycle_s_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_1_34_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_fastZ0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_1_19_0\ : std_logic;
signal \POWERLED.un45_slp_s3n\ : std_logic;
signal \POWERLED.N_174\ : std_logic;
signal \POWERLED.N_77\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_1_sqmuxa_i_1\ : std_logic;
signal \SLP_S3n_c\ : std_logic;
signal \VCCST_EN_c\ : std_logic;
signal \VCCST_EN_c_cascade_\ : std_logic;
signal \POWERLED.N_162\ : std_logic;
signal \SLP_S4n_c\ : std_logic;
signal \RSMRSTn_c\ : std_logic;
signal \slp_s4n_signal_i_0_cascade_\ : std_logic;
signal \VDDQ_OK_c\ : std_logic;
signal \VPP_VDDQ.N_181\ : std_logic;
signal slp_s4n_signal_i_0 : std_logic;
signal \POWERLED.func_state_ns_0_i_0_0_0\ : std_logic;
signal \POWERLED.N_120\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \FPGA_OSC_0_c_g\ : std_logic;
signal \N_39_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \FPGA_OSC_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;

begin
    \FPGA_OSC_wire\ <= FPGA_OSC;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \V5A_OK_wire\ <= V5A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    VDDQ_EN <= \VDDQ_EN_wire\;
    V5S_ENn <= \V5S_ENn_wire\;
    V5A_EN <= \V5A_EN_wire\;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    \SLP_S4n_wire\ <= SLP_S4n;
    \SLP_S3n_wire\ <= SLP_S3n;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    VCCST_EN <= \VCCST_EN_wire\;
    \VPP_OK_wire\ <= VPP_OK;
    V33A_ENn <= \V33A_ENn_wire\;
    \V5S_OK_wire\ <= V5S_OK;
    \V33A_OK_wire\ <= V33A_OK;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VPP_EN <= \VPP_EN_wire\;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    V33S_ENn <= \V33S_ENn_wire\;
    RSMRSTn <= \RSMRSTn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    SUSWARN_N <= \SUSWARN_N_wire\;
    DSW_PWROK <= \DSW_PWROK_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;

    \FPGA_OSC_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__18891\,
            GLOBALBUFFEROUTPUT => \FPGA_OSC_0_c_g\
        );

    \FPGA_OSC_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18893\,
            DIN => \N__18892\,
            DOUT => \N__18891\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \FPGA_OSC_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18893\,
            PADOUT => \N__18892\,
            PADIN => \N__18891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V1P8A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__18882\,
            DIN => \N__18881\,
            DOUT => \N__18880\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \V1P8A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18882\,
            PADOUT => \N__18881\,
            PADIN => \N__18880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V1P8A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__18873\,
            DIN => \N__18872\,
            DOUT => \N__18871\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \V5A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18873\,
            PADOUT => \N__18872\,
            PADIN => \N__18871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCH_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18864\,
            DIN => \N__18863\,
            DOUT => \N__18862\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \PCH_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18864\,
            PADOUT => \N__18863\,
            PADIN => \N__18862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7855\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCINAUX_VR_PE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18855\,
            DIN => \N__18854\,
            DOUT => \N__18853\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \VCCINAUX_VR_PE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18855\,
            PADOUT => \N__18854\,
            PADIN => \N__18853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCIN_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18846\,
            DIN => \N__18845\,
            DOUT => \N__18844\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \VCCIN_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18846\,
            PADOUT => \N__18845\,
            PADIN => \N__18844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14255\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33S_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18837\,
            DIN => \N__18836\,
            DOUT => \N__18835\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \V33S_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18837\,
            PADOUT => \N__18836\,
            PADIN => \N__18835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33S_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VDDQ_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18828\,
            DIN => \N__18827\,
            DOUT => \N__18826\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \VDDQ_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18828\,
            PADOUT => \N__18827\,
            PADIN => \N__18826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8078\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5S_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18819\,
            DIN => \N__18818\,
            DOUT => \N__18817\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \V5S_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18819\,
            PADOUT => \N__18818\,
            PADIN => \N__18817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18810\,
            DIN => \N__18809\,
            DOUT => \N__18808\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \V5A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18810\,
            PADOUT => \N__18809\,
            PADIN => \N__18808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12150\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCINAUX_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18801\,
            DIN => \N__18800\,
            DOUT => \N__18799\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \VCCINAUX_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18801\,
            PADOUT => \N__18800\,
            PADIN => \N__18799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12080\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCIN_VR_PE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18792\,
            DIN => \N__18791\,
            DOUT => \N__18790\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \VCCIN_VR_PE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18792\,
            PADOUT => \N__18791\,
            PADIN => \N__18790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_S4n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18783\,
            DIN => \N__18782\,
            DOUT => \N__18781\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \SLP_S4n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18783\,
            PADOUT => \N__18782\,
            PADIN => \N__18781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SLP_S4n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_S3n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18774\,
            DIN => \N__18773\,
            DOUT => \N__18772\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \SLP_S3n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18774\,
            PADOUT => \N__18773\,
            PADIN => \N__18772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SLP_S3n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_PWRGD_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18765\,
            DIN => \N__18764\,
            DOUT => \N__18763\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \VCCST_PWRGD_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18765\,
            PADOUT => \N__18764\,
            PADIN => \N__18763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_SUSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18756\,
            DIN => \N__18755\,
            DOUT => \N__18754\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \SLP_SUSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18756\,
            PADOUT => \N__18755\,
            PADIN => \N__18754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5A_EN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HDA_SDO_ATP_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18747\,
            DIN => \N__18746\,
            DOUT => \N__18745\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \HDA_SDO_ATP_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18747\,
            PADOUT => \N__18746\,
            PADIN => \N__18745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18738\,
            DIN => \N__18737\,
            DOUT => \N__18736\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \VCCST_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18738\,
            PADOUT => \N__18737\,
            PADIN => \N__18736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VPP_OK_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__18729\,
            DIN => \N__18728\,
            DOUT => \N__18727\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \VPP_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18729\,
            PADOUT => \N__18728\,
            PADIN => \N__18727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VPP_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33A_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18720\,
            DIN => \N__18719\,
            DOUT => \N__18718\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \V33A_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18720\,
            PADOUT => \N__18719\,
            PADIN => \N__18718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5S_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18711\,
            DIN => \N__18710\,
            DOUT => \N__18709\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \V5S_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18711\,
            PADOUT => \N__18710\,
            PADIN => \N__18709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5S_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18702\,
            DIN => \N__18701\,
            DOUT => \N__18700\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \V33A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18702\,
            PADOUT => \N__18701\,
            PADIN => \N__18700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_CPU_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18693\,
            DIN => \N__18692\,
            DOUT => \N__18691\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \VCCST_CPU_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18693\,
            PADOUT => \N__18692\,
            PADIN => \N__18691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VCCST_CPU_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VPP_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18684\,
            DIN => \N__18683\,
            DOUT => \N__18682\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \VPP_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18684\,
            PADOUT => \N__18683\,
            PADIN => \N__18682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13139\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWRBTN_LED_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18675\,
            DIN => \N__18674\,
            DOUT => \N__18673\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \PWRBTN_LED_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18675\,
            PADOUT => \N__18674\,
            PADIN => \N__18673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33S_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18666\,
            DIN => \N__18665\,
            DOUT => \N__18664\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \V33S_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18666\,
            PADOUT => \N__18665\,
            PADIN => \N__18664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RSMRSTn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18657\,
            DIN => \N__18656\,
            DOUT => \N__18655\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \RSMRSTn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18657\,
            PADOUT => \N__18656\,
            PADIN => \N__18655\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18518\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V1P8A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18648\,
            DIN => \N__18647\,
            DOUT => \N__18646\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \V1P8A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18648\,
            PADOUT => \N__18647\,
            PADIN => \N__18646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12151\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VDDQ_OK_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__18639\,
            DIN => \N__18638\,
            DOUT => \N__18637\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \VDDQ_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18639\,
            PADOUT => \N__18638\,
            PADIN => \N__18637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VDDQ_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SUSWARN_N_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18630\,
            DIN => \N__18629\,
            DOUT => \N__18628\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \SUSWARN_N_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18630\,
            PADOUT => \N__18629\,
            PADIN => \N__18628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14254\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DSW_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18621\,
            DIN => \N__18620\,
            DOUT => \N__18619\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \DSW_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18621\,
            PADOUT => \N__18620\,
            PADIN => \N__18619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14946\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SYS_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18612\,
            DIN => \N__18611\,
            DOUT => \N__18610\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \SYS_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18612\,
            PADOUT => \N__18611\,
            PADIN => \N__18610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7865\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VR_READY_VCCIN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18603\,
            DIN => \N__18602\,
            DOUT => \N__18601\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \VR_READY_VCCIN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18603\,
            PADOUT => \N__18602\,
            PADIN => \N__18601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VR_READY_VCCIN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4260\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18577\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18574\
        );

    \I__4258\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18568\
        );

    \I__4257\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18568\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18565\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18558\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18574\,
            I => \N__18558\
        );

    \I__4253\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18555\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__18568\,
            I => \N__18550\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__18565\,
            I => \N__18550\
        );

    \I__4250\ : InMux
    port map (
            O => \N__18564\,
            I => \N__18547\
        );

    \I__4249\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18544\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__18558\,
            I => \N__18541\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__18555\,
            I => \N__18538\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__18550\,
            I => \N__18531\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18531\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__18544\,
            I => \N__18531\
        );

    \I__4243\ : Span4Mux_h
    port map (
            O => \N__18541\,
            I => \N__18524\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__18538\,
            I => \N__18524\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__18531\,
            I => \N__18524\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__18521\,
            I => \SLP_S4n_c\
        );

    \I__4238\ : IoInMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__4236\ : IoSpan4Mux
    port map (
            O => \N__18512\,
            I => \N__18507\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__18511\,
            I => \N__18503\
        );

    \I__4234\ : InMux
    port map (
            O => \N__18510\,
            I => \N__18498\
        );

    \I__4233\ : Span4Mux_s2_v
    port map (
            O => \N__18507\,
            I => \N__18493\
        );

    \I__4232\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18490\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18487\
        );

    \I__4230\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18482\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18482\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18498\,
            I => \N__18479\
        );

    \I__4227\ : InMux
    port map (
            O => \N__18497\,
            I => \N__18474\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18474\
        );

    \I__4225\ : Span4Mux_h
    port map (
            O => \N__18493\,
            I => \N__18469\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__18490\,
            I => \N__18469\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18487\,
            I => \N__18460\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18460\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__18479\,
            I => \N__18460\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__18474\,
            I => \N__18460\
        );

    \I__4219\ : Span4Mux_v
    port map (
            O => \N__18469\,
            I => \N__18457\
        );

    \I__4218\ : Span4Mux_v
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__18454\,
            I => \N__18448\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__18451\,
            I => \N__18445\
        );

    \I__4214\ : Span4Mux_v
    port map (
            O => \N__18448\,
            I => \N__18442\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__18445\,
            I => \RSMRSTn_c\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__18442\,
            I => \RSMRSTn_c\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \slp_s4n_signal_i_0_cascade_\
        );

    \I__4210\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__4208\ : Span4Mux_s0_h
    port map (
            O => \N__18428\,
            I => \N__18424\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__4206\ : Span4Mux_v
    port map (
            O => \N__18424\,
            I => \N__18416\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18421\,
            I => \N__18416\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__18413\,
            I => \VDDQ_OK_c\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__4201\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18402\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18399\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18396\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__18402\,
            I => \N__18392\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__18399\,
            I => \N__18389\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__18396\,
            I => \N__18386\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18383\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__18392\,
            I => \N__18377\
        );

    \I__4193\ : Span4Mux_v
    port map (
            O => \N__18389\,
            I => \N__18377\
        );

    \I__4192\ : Span4Mux_v
    port map (
            O => \N__18386\,
            I => \N__18374\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18371\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18368\
        );

    \I__4189\ : Sp12to4
    port map (
            O => \N__18377\,
            I => \N__18359\
        );

    \I__4188\ : Sp12to4
    port map (
            O => \N__18374\,
            I => \N__18359\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__18371\,
            I => \N__18359\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__18368\,
            I => \N__18359\
        );

    \I__4185\ : Odrv12
    port map (
            O => \N__18359\,
            I => \VPP_VDDQ.N_181\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18352\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18349\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18346\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__18349\,
            I => \N__18343\
        );

    \I__4180\ : Span4Mux_v
    port map (
            O => \N__18346\,
            I => \N__18336\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__18343\,
            I => \N__18330\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18327\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18320\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18320\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18320\
        );

    \I__4174\ : Span4Mux_h
    port map (
            O => \N__18336\,
            I => \N__18317\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18312\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18312\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18308\
        );

    \I__4170\ : Span4Mux_h
    port map (
            O => \N__18330\,
            I => \N__18301\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18301\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__18320\,
            I => \N__18301\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__18317\,
            I => \N__18296\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18312\,
            I => \N__18296\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18293\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__18308\,
            I => slp_s4n_signal_i_0
        );

    \I__4163\ : Odrv4
    port map (
            O => \N__18301\,
            I => slp_s4n_signal_i_0
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__18296\,
            I => slp_s4n_signal_i_0
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__18293\,
            I => slp_s4n_signal_i_0
        );

    \I__4160\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18281\,
            I => \POWERLED.func_state_ns_0_i_0_0_0\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__18278\,
            I => \N__18274\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18271\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18271\,
            I => \POWERLED.N_120\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__18268\,
            I => \POWERLED.N_120\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__18263\,
            I => \N__18255\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18249\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18249\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18244\
        );

    \I__4149\ : InMux
    port map (
            O => \N__18259\,
            I => \N__18244\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__18258\,
            I => \N__18240\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18235\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18232\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18249\,
            I => \N__18227\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__18244\,
            I => \N__18227\
        );

    \I__4143\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18218\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18218\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18218\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18218\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18235\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18232\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__18227\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__18218\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4135\ : ClkMux
    port map (
            O => \N__18209\,
            I => \N__18074\
        );

    \I__4134\ : ClkMux
    port map (
            O => \N__18208\,
            I => \N__18074\
        );

    \I__4133\ : ClkMux
    port map (
            O => \N__18207\,
            I => \N__18074\
        );

    \I__4132\ : ClkMux
    port map (
            O => \N__18206\,
            I => \N__18074\
        );

    \I__4131\ : ClkMux
    port map (
            O => \N__18205\,
            I => \N__18074\
        );

    \I__4130\ : ClkMux
    port map (
            O => \N__18204\,
            I => \N__18074\
        );

    \I__4129\ : ClkMux
    port map (
            O => \N__18203\,
            I => \N__18074\
        );

    \I__4128\ : ClkMux
    port map (
            O => \N__18202\,
            I => \N__18074\
        );

    \I__4127\ : ClkMux
    port map (
            O => \N__18201\,
            I => \N__18074\
        );

    \I__4126\ : ClkMux
    port map (
            O => \N__18200\,
            I => \N__18074\
        );

    \I__4125\ : ClkMux
    port map (
            O => \N__18199\,
            I => \N__18074\
        );

    \I__4124\ : ClkMux
    port map (
            O => \N__18198\,
            I => \N__18074\
        );

    \I__4123\ : ClkMux
    port map (
            O => \N__18197\,
            I => \N__18074\
        );

    \I__4122\ : ClkMux
    port map (
            O => \N__18196\,
            I => \N__18074\
        );

    \I__4121\ : ClkMux
    port map (
            O => \N__18195\,
            I => \N__18074\
        );

    \I__4120\ : ClkMux
    port map (
            O => \N__18194\,
            I => \N__18074\
        );

    \I__4119\ : ClkMux
    port map (
            O => \N__18193\,
            I => \N__18074\
        );

    \I__4118\ : ClkMux
    port map (
            O => \N__18192\,
            I => \N__18074\
        );

    \I__4117\ : ClkMux
    port map (
            O => \N__18191\,
            I => \N__18074\
        );

    \I__4116\ : ClkMux
    port map (
            O => \N__18190\,
            I => \N__18074\
        );

    \I__4115\ : ClkMux
    port map (
            O => \N__18189\,
            I => \N__18074\
        );

    \I__4114\ : ClkMux
    port map (
            O => \N__18188\,
            I => \N__18074\
        );

    \I__4113\ : ClkMux
    port map (
            O => \N__18187\,
            I => \N__18074\
        );

    \I__4112\ : ClkMux
    port map (
            O => \N__18186\,
            I => \N__18074\
        );

    \I__4111\ : ClkMux
    port map (
            O => \N__18185\,
            I => \N__18074\
        );

    \I__4110\ : ClkMux
    port map (
            O => \N__18184\,
            I => \N__18074\
        );

    \I__4109\ : ClkMux
    port map (
            O => \N__18183\,
            I => \N__18074\
        );

    \I__4108\ : ClkMux
    port map (
            O => \N__18182\,
            I => \N__18074\
        );

    \I__4107\ : ClkMux
    port map (
            O => \N__18181\,
            I => \N__18074\
        );

    \I__4106\ : ClkMux
    port map (
            O => \N__18180\,
            I => \N__18074\
        );

    \I__4105\ : ClkMux
    port map (
            O => \N__18179\,
            I => \N__18074\
        );

    \I__4104\ : ClkMux
    port map (
            O => \N__18178\,
            I => \N__18074\
        );

    \I__4103\ : ClkMux
    port map (
            O => \N__18177\,
            I => \N__18074\
        );

    \I__4102\ : ClkMux
    port map (
            O => \N__18176\,
            I => \N__18074\
        );

    \I__4101\ : ClkMux
    port map (
            O => \N__18175\,
            I => \N__18074\
        );

    \I__4100\ : ClkMux
    port map (
            O => \N__18174\,
            I => \N__18074\
        );

    \I__4099\ : ClkMux
    port map (
            O => \N__18173\,
            I => \N__18074\
        );

    \I__4098\ : ClkMux
    port map (
            O => \N__18172\,
            I => \N__18074\
        );

    \I__4097\ : ClkMux
    port map (
            O => \N__18171\,
            I => \N__18074\
        );

    \I__4096\ : ClkMux
    port map (
            O => \N__18170\,
            I => \N__18074\
        );

    \I__4095\ : ClkMux
    port map (
            O => \N__18169\,
            I => \N__18074\
        );

    \I__4094\ : ClkMux
    port map (
            O => \N__18168\,
            I => \N__18074\
        );

    \I__4093\ : ClkMux
    port map (
            O => \N__18167\,
            I => \N__18074\
        );

    \I__4092\ : ClkMux
    port map (
            O => \N__18166\,
            I => \N__18074\
        );

    \I__4091\ : ClkMux
    port map (
            O => \N__18165\,
            I => \N__18074\
        );

    \I__4090\ : GlobalMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__4089\ : gio2CtrlBuf
    port map (
            O => \N__18071\,
            I => \FPGA_OSC_0_c_g\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__18068\,
            I => \N__18010\
        );

    \I__4087\ : InMux
    port map (
            O => \N__18067\,
            I => \N__17937\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18066\,
            I => \N__17937\
        );

    \I__4085\ : InMux
    port map (
            O => \N__18065\,
            I => \N__17937\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18064\,
            I => \N__17937\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18063\,
            I => \N__17928\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18062\,
            I => \N__17928\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18061\,
            I => \N__17928\
        );

    \I__4080\ : InMux
    port map (
            O => \N__18060\,
            I => \N__17928\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18059\,
            I => \N__17919\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18058\,
            I => \N__17919\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18057\,
            I => \N__17919\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18056\,
            I => \N__17919\
        );

    \I__4075\ : InMux
    port map (
            O => \N__18055\,
            I => \N__17910\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18054\,
            I => \N__17910\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18053\,
            I => \N__17910\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18052\,
            I => \N__17910\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18051\,
            I => \N__17901\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18050\,
            I => \N__17901\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18049\,
            I => \N__17901\
        );

    \I__4068\ : InMux
    port map (
            O => \N__18048\,
            I => \N__17901\
        );

    \I__4067\ : InMux
    port map (
            O => \N__18047\,
            I => \N__17892\
        );

    \I__4066\ : InMux
    port map (
            O => \N__18046\,
            I => \N__17892\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18045\,
            I => \N__17892\
        );

    \I__4064\ : InMux
    port map (
            O => \N__18044\,
            I => \N__17892\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18043\,
            I => \N__17883\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18042\,
            I => \N__17883\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18041\,
            I => \N__17883\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18040\,
            I => \N__17883\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18039\,
            I => \N__17874\
        );

    \I__4058\ : InMux
    port map (
            O => \N__18038\,
            I => \N__17874\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18037\,
            I => \N__17874\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18036\,
            I => \N__17874\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18035\,
            I => \N__17865\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18034\,
            I => \N__17865\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18033\,
            I => \N__17865\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18032\,
            I => \N__17865\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18031\,
            I => \N__17856\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18030\,
            I => \N__17856\
        );

    \I__4049\ : InMux
    port map (
            O => \N__18029\,
            I => \N__17856\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18028\,
            I => \N__17856\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18027\,
            I => \N__17847\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18026\,
            I => \N__17847\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18025\,
            I => \N__17847\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18024\,
            I => \N__17847\
        );

    \I__4043\ : InMux
    port map (
            O => \N__18023\,
            I => \N__17838\
        );

    \I__4042\ : InMux
    port map (
            O => \N__18022\,
            I => \N__17838\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18021\,
            I => \N__17838\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18020\,
            I => \N__17838\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18019\,
            I => \N__17829\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18018\,
            I => \N__17829\
        );

    \I__4037\ : InMux
    port map (
            O => \N__18017\,
            I => \N__17829\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18016\,
            I => \N__17829\
        );

    \I__4035\ : InMux
    port map (
            O => \N__18015\,
            I => \N__17822\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18014\,
            I => \N__17822\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18013\,
            I => \N__17822\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18010\,
            I => \N__17817\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18009\,
            I => \N__17817\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18008\,
            I => \N__17808\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17808\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18006\,
            I => \N__17808\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18005\,
            I => \N__17808\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17799\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17799\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17799\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18001\,
            I => \N__17799\
        );

    \I__4022\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17792\
        );

    \I__4021\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17792\
        );

    \I__4020\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17792\
        );

    \I__4019\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17783\
        );

    \I__4018\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17783\
        );

    \I__4017\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17783\
        );

    \I__4016\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17783\
        );

    \I__4015\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17776\
        );

    \I__4014\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17776\
        );

    \I__4013\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17776\
        );

    \I__4012\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17769\
        );

    \I__4011\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17769\
        );

    \I__4010\ : InMux
    port map (
            O => \N__17988\,
            I => \N__17769\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17987\,
            I => \N__17760\
        );

    \I__4008\ : InMux
    port map (
            O => \N__17986\,
            I => \N__17760\
        );

    \I__4007\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17760\
        );

    \I__4006\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17760\
        );

    \I__4005\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17751\
        );

    \I__4004\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17751\
        );

    \I__4003\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17751\
        );

    \I__4002\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17751\
        );

    \I__4001\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17744\
        );

    \I__4000\ : InMux
    port map (
            O => \N__17978\,
            I => \N__17744\
        );

    \I__3999\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17744\
        );

    \I__3998\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17737\
        );

    \I__3997\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17737\
        );

    \I__3996\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17737\
        );

    \I__3995\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17728\
        );

    \I__3994\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17728\
        );

    \I__3993\ : InMux
    port map (
            O => \N__17971\,
            I => \N__17728\
        );

    \I__3992\ : InMux
    port map (
            O => \N__17970\,
            I => \N__17728\
        );

    \I__3991\ : InMux
    port map (
            O => \N__17969\,
            I => \N__17721\
        );

    \I__3990\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17721\
        );

    \I__3989\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17721\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17714\
        );

    \I__3987\ : InMux
    port map (
            O => \N__17965\,
            I => \N__17714\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17714\
        );

    \I__3985\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17707\
        );

    \I__3984\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17707\
        );

    \I__3983\ : InMux
    port map (
            O => \N__17961\,
            I => \N__17707\
        );

    \I__3982\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17704\
        );

    \I__3981\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17701\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17958\,
            I => \N__17698\
        );

    \I__3979\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17695\
        );

    \I__3978\ : InMux
    port map (
            O => \N__17956\,
            I => \N__17692\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17955\,
            I => \N__17687\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17687\
        );

    \I__3975\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17682\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17682\
        );

    \I__3973\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17677\
        );

    \I__3972\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17677\
        );

    \I__3971\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17674\
        );

    \I__3970\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17671\
        );

    \I__3969\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17668\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17665\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__17937\,
            I => \N__17648\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__17928\,
            I => \N__17645\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__17919\,
            I => \N__17642\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__17910\,
            I => \N__17639\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__17901\,
            I => \N__17636\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__17892\,
            I => \N__17633\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__17883\,
            I => \N__17630\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__17874\,
            I => \N__17627\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__17865\,
            I => \N__17624\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__17856\,
            I => \N__17621\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17618\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17615\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17829\,
            I => \N__17612\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17609\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__17817\,
            I => \N__17606\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17603\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__17799\,
            I => \N__17600\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__17792\,
            I => \N__17597\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17594\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__17776\,
            I => \N__17591\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__17769\,
            I => \N__17588\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__17760\,
            I => \N__17585\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__17751\,
            I => \N__17582\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__17744\,
            I => \N__17579\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__17737\,
            I => \N__17576\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17573\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__17721\,
            I => \N__17570\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17567\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__17707\,
            I => \N__17564\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__17704\,
            I => \N__17561\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__17701\,
            I => \N__17558\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__17698\,
            I => \N__17555\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17695\,
            I => \N__17552\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17549\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17546\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__17682\,
            I => \N__17543\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__17677\,
            I => \N__17540\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__17674\,
            I => \N__17537\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17534\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17531\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__17665\,
            I => \N__17528\
        );

    \I__3926\ : CEMux
    port map (
            O => \N__17664\,
            I => \N__17417\
        );

    \I__3925\ : CEMux
    port map (
            O => \N__17663\,
            I => \N__17417\
        );

    \I__3924\ : CEMux
    port map (
            O => \N__17662\,
            I => \N__17417\
        );

    \I__3923\ : CEMux
    port map (
            O => \N__17661\,
            I => \N__17417\
        );

    \I__3922\ : CEMux
    port map (
            O => \N__17660\,
            I => \N__17417\
        );

    \I__3921\ : CEMux
    port map (
            O => \N__17659\,
            I => \N__17417\
        );

    \I__3920\ : CEMux
    port map (
            O => \N__17658\,
            I => \N__17417\
        );

    \I__3919\ : CEMux
    port map (
            O => \N__17657\,
            I => \N__17417\
        );

    \I__3918\ : CEMux
    port map (
            O => \N__17656\,
            I => \N__17417\
        );

    \I__3917\ : CEMux
    port map (
            O => \N__17655\,
            I => \N__17417\
        );

    \I__3916\ : CEMux
    port map (
            O => \N__17654\,
            I => \N__17417\
        );

    \I__3915\ : CEMux
    port map (
            O => \N__17653\,
            I => \N__17417\
        );

    \I__3914\ : CEMux
    port map (
            O => \N__17652\,
            I => \N__17417\
        );

    \I__3913\ : CEMux
    port map (
            O => \N__17651\,
            I => \N__17417\
        );

    \I__3912\ : Glb2LocalMux
    port map (
            O => \N__17648\,
            I => \N__17417\
        );

    \I__3911\ : Glb2LocalMux
    port map (
            O => \N__17645\,
            I => \N__17417\
        );

    \I__3910\ : Glb2LocalMux
    port map (
            O => \N__17642\,
            I => \N__17417\
        );

    \I__3909\ : Glb2LocalMux
    port map (
            O => \N__17639\,
            I => \N__17417\
        );

    \I__3908\ : Glb2LocalMux
    port map (
            O => \N__17636\,
            I => \N__17417\
        );

    \I__3907\ : Glb2LocalMux
    port map (
            O => \N__17633\,
            I => \N__17417\
        );

    \I__3906\ : Glb2LocalMux
    port map (
            O => \N__17630\,
            I => \N__17417\
        );

    \I__3905\ : Glb2LocalMux
    port map (
            O => \N__17627\,
            I => \N__17417\
        );

    \I__3904\ : Glb2LocalMux
    port map (
            O => \N__17624\,
            I => \N__17417\
        );

    \I__3903\ : Glb2LocalMux
    port map (
            O => \N__17621\,
            I => \N__17417\
        );

    \I__3902\ : Glb2LocalMux
    port map (
            O => \N__17618\,
            I => \N__17417\
        );

    \I__3901\ : Glb2LocalMux
    port map (
            O => \N__17615\,
            I => \N__17417\
        );

    \I__3900\ : Glb2LocalMux
    port map (
            O => \N__17612\,
            I => \N__17417\
        );

    \I__3899\ : Glb2LocalMux
    port map (
            O => \N__17609\,
            I => \N__17417\
        );

    \I__3898\ : Glb2LocalMux
    port map (
            O => \N__17606\,
            I => \N__17417\
        );

    \I__3897\ : Glb2LocalMux
    port map (
            O => \N__17603\,
            I => \N__17417\
        );

    \I__3896\ : Glb2LocalMux
    port map (
            O => \N__17600\,
            I => \N__17417\
        );

    \I__3895\ : Glb2LocalMux
    port map (
            O => \N__17597\,
            I => \N__17417\
        );

    \I__3894\ : Glb2LocalMux
    port map (
            O => \N__17594\,
            I => \N__17417\
        );

    \I__3893\ : Glb2LocalMux
    port map (
            O => \N__17591\,
            I => \N__17417\
        );

    \I__3892\ : Glb2LocalMux
    port map (
            O => \N__17588\,
            I => \N__17417\
        );

    \I__3891\ : Glb2LocalMux
    port map (
            O => \N__17585\,
            I => \N__17417\
        );

    \I__3890\ : Glb2LocalMux
    port map (
            O => \N__17582\,
            I => \N__17417\
        );

    \I__3889\ : Glb2LocalMux
    port map (
            O => \N__17579\,
            I => \N__17417\
        );

    \I__3888\ : Glb2LocalMux
    port map (
            O => \N__17576\,
            I => \N__17417\
        );

    \I__3887\ : Glb2LocalMux
    port map (
            O => \N__17573\,
            I => \N__17417\
        );

    \I__3886\ : Glb2LocalMux
    port map (
            O => \N__17570\,
            I => \N__17417\
        );

    \I__3885\ : Glb2LocalMux
    port map (
            O => \N__17567\,
            I => \N__17417\
        );

    \I__3884\ : Glb2LocalMux
    port map (
            O => \N__17564\,
            I => \N__17417\
        );

    \I__3883\ : Glb2LocalMux
    port map (
            O => \N__17561\,
            I => \N__17417\
        );

    \I__3882\ : Glb2LocalMux
    port map (
            O => \N__17558\,
            I => \N__17417\
        );

    \I__3881\ : Glb2LocalMux
    port map (
            O => \N__17555\,
            I => \N__17417\
        );

    \I__3880\ : Glb2LocalMux
    port map (
            O => \N__17552\,
            I => \N__17417\
        );

    \I__3879\ : Glb2LocalMux
    port map (
            O => \N__17549\,
            I => \N__17417\
        );

    \I__3878\ : Glb2LocalMux
    port map (
            O => \N__17546\,
            I => \N__17417\
        );

    \I__3877\ : Glb2LocalMux
    port map (
            O => \N__17543\,
            I => \N__17417\
        );

    \I__3876\ : Glb2LocalMux
    port map (
            O => \N__17540\,
            I => \N__17417\
        );

    \I__3875\ : Glb2LocalMux
    port map (
            O => \N__17537\,
            I => \N__17417\
        );

    \I__3874\ : Glb2LocalMux
    port map (
            O => \N__17534\,
            I => \N__17417\
        );

    \I__3873\ : Glb2LocalMux
    port map (
            O => \N__17531\,
            I => \N__17417\
        );

    \I__3872\ : Glb2LocalMux
    port map (
            O => \N__17528\,
            I => \N__17417\
        );

    \I__3871\ : GlobalMux
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3870\ : gio2CtrlBuf
    port map (
            O => \N__17414\,
            I => \N_39_g\
        );

    \I__3869\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17393\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17388\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17379\
        );

    \I__3866\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17379\
        );

    \I__3865\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17379\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17379\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17405\,
            I => \N__17376\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17367\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17367\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17367\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17367\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17362\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17362\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17359\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17354\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17354\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17393\,
            I => \N__17351\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17348\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17345\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__17388\,
            I => \N__17342\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17379\,
            I => \N__17337\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17376\,
            I => \N__17337\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17334\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17362\,
            I => \N__17331\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17328\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17325\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__17351\,
            I => \N__17322\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17348\,
            I => \N__17319\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17345\,
            I => \N__17314\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__17342\,
            I => \N__17314\
        );

    \I__3839\ : Span4Mux_h
    port map (
            O => \N__17337\,
            I => \N__17311\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__17334\,
            I => \N__17306\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__17331\,
            I => \N__17306\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__17328\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__17325\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__17322\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3833\ : Odrv12
    port map (
            O => \N__17319\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__17314\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__17311\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__17306\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3829\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17288\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__17288\,
            I => \N__17284\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17287\,
            I => \N__17281\
        );

    \I__3826\ : Span4Mux_s2_h
    port map (
            O => \N__17284\,
            I => \N__17278\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__17281\,
            I => \N__17275\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__17278\,
            I => \POWERLED.dutycycle_s_5\
        );

    \I__3823\ : Odrv12
    port map (
            O => \N__17275\,
            I => \POWERLED.dutycycle_s_5\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \N__17265\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__17269\,
            I => \N__17262\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17268\,
            I => \N__17254\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17251\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17246\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17246\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__17260\,
            I => \N__17243\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__17259\,
            I => \N__17240\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__17258\,
            I => \N__17237\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__17257\,
            I => \N__17233\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17254\,
            I => \N__17226\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17251\,
            I => \N__17226\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__17246\,
            I => \N__17226\
        );

    \I__3809\ : InMux
    port map (
            O => \N__17243\,
            I => \N__17223\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17240\,
            I => \N__17220\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17213\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17213\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17213\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__17226\,
            I => \N__17208\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__17223\,
            I => \N__17208\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__17220\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17213\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__17208\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__17198\,
            I => \POWERLED.un1_dutycycle_1_34_0\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17188\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__17194\,
            I => \N__17185\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17178\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17173\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17173\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17188\,
            I => \N__17170\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17165\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17165\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17162\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17157\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17181\,
            I => \N__17157\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17178\,
            I => \N__17152\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17152\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__17170\,
            I => \N__17149\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17146\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17162\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__17157\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__17152\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__17149\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__17146\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__17135\,
            I => \N__17132\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17127\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17131\,
            I => \N__17124\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17130\,
            I => \N__17121\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17127\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17124\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17121\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__3770\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__17111\,
            I => \POWERLED.un1_dutycycle_1_19_0\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__17108\,
            I => \N__17104\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__17107\,
            I => \N__17101\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17097\
        );

    \I__3765\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17094\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__17100\,
            I => \N__17091\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17097\,
            I => \N__17087\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17094\,
            I => \N__17084\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17080\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17077\
        );

    \I__3759\ : Span4Mux_h
    port map (
            O => \N__17087\,
            I => \N__17074\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__17084\,
            I => \N__17071\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17068\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__17080\,
            I => \POWERLED.un45_slp_s3n\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17077\,
            I => \POWERLED.un45_slp_s3n\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__17074\,
            I => \POWERLED.un45_slp_s3n\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__17071\,
            I => \POWERLED.un45_slp_s3n\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17068\,
            I => \POWERLED.un45_slp_s3n\
        );

    \I__3751\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17054\,
            I => \POWERLED.N_174\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17045\,
            I => \N__17041\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17038\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__17041\,
            I => \POWERLED.N_77\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17038\,
            I => \POWERLED.N_77\
        );

    \I__3743\ : InMux
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__17024\,
            I => \POWERLED.un2_slp_s3n_2_0_0\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__17021\,
            I => \N__17016\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__17020\,
            I => \N__17013\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17006\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17016\,
            I => \N__17001\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17001\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17012\,
            I => \N__16996\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17011\,
            I => \N__16996\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17010\,
            I => \N__16993\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17009\,
            I => \N__16990\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__17006\,
            I => \N__16987\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17001\,
            I => \N__16980\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16980\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__16993\,
            I => \N__16980\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__16990\,
            I => \N__16973\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__16987\,
            I => \N__16973\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__16980\,
            I => \N__16973\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__16973\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__16967\,
            I => \POWERLED.dutycycle_1_sqmuxa_i_1\
        );

    \I__3720\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16957\
        );

    \I__3719\ : InMux
    port map (
            O => \N__16963\,
            I => \N__16957\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__16962\,
            I => \N__16954\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__16957\,
            I => \N__16949\
        );

    \I__3716\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16946\
        );

    \I__3715\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16943\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__16952\,
            I => \N__16940\
        );

    \I__3713\ : Span4Mux_s0_h
    port map (
            O => \N__16949\,
            I => \N__16932\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__16946\,
            I => \N__16932\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__16943\,
            I => \N__16932\
        );

    \I__3710\ : InMux
    port map (
            O => \N__16940\,
            I => \N__16929\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__16939\,
            I => \N__16925\
        );

    \I__3708\ : Span4Mux_v
    port map (
            O => \N__16932\,
            I => \N__16921\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16918\
        );

    \I__3706\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16913\
        );

    \I__3705\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16913\
        );

    \I__3704\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16910\
        );

    \I__3703\ : IoSpan4Mux
    port map (
            O => \N__16921\,
            I => \N__16907\
        );

    \I__3702\ : Span4Mux_h
    port map (
            O => \N__16918\,
            I => \N__16904\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__16913\,
            I => \N__16899\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__16910\,
            I => \N__16899\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__16907\,
            I => \SLP_S3n_c\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__16904\,
            I => \SLP_S3n_c\
        );

    \I__3697\ : Odrv12
    port map (
            O => \N__16899\,
            I => \SLP_S3n_c\
        );

    \I__3696\ : IoInMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__3694\ : IoSpan4Mux
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__3693\ : Span4Mux_s2_h
    port map (
            O => \N__16883\,
            I => \N__16878\
        );

    \I__3692\ : InMux
    port map (
            O => \N__16882\,
            I => \N__16875\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__16881\,
            I => \N__16871\
        );

    \I__3690\ : Sp12to4
    port map (
            O => \N__16878\,
            I => \N__16864\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__16875\,
            I => \N__16864\
        );

    \I__3688\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16861\
        );

    \I__3687\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16858\
        );

    \I__3686\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16855\
        );

    \I__3685\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16852\
        );

    \I__3684\ : Span12Mux_s7_h
    port map (
            O => \N__16864\,
            I => \N__16845\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16845\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__16858\,
            I => \N__16845\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__16855\,
            I => \VCCST_EN_c\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__16852\,
            I => \VCCST_EN_c\
        );

    \I__3679\ : Odrv12
    port map (
            O => \N__16845\,
            I => \VCCST_EN_c\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__16838\,
            I => \VCCST_EN_c_cascade_\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__16835\,
            I => \N__16831\
        );

    \I__3676\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16826\
        );

    \I__3675\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16823\
        );

    \I__3674\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16820\
        );

    \I__3673\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16817\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__16826\,
            I => \N__16814\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16809\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__16820\,
            I => \N__16806\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__16817\,
            I => \N__16803\
        );

    \I__3668\ : Span4Mux_v
    port map (
            O => \N__16814\,
            I => \N__16800\
        );

    \I__3667\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16797\
        );

    \I__3666\ : InMux
    port map (
            O => \N__16812\,
            I => \N__16794\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__16809\,
            I => \POWERLED.N_162\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__16806\,
            I => \POWERLED.N_162\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__16803\,
            I => \POWERLED.N_162\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__16800\,
            I => \POWERLED.N_162\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__16797\,
            I => \POWERLED.N_162\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__16794\,
            I => \POWERLED.N_162\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16775\
        );

    \I__3658\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16775\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__16775\,
            I => \POWERLED.N_115\
        );

    \I__3656\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16763\
        );

    \I__3655\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16763\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16763\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__16760\,
            I => \POWERLED.N_92\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__16757\,
            I => \POWERLED.N_120_cascade_\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16750\
        );

    \I__3649\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16747\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__16750\,
            I => \N__16743\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16747\,
            I => \N__16740\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16746\,
            I => \N__16737\
        );

    \I__3645\ : Span4Mux_v
    port map (
            O => \N__16743\,
            I => \N__16732\
        );

    \I__3644\ : Span4Mux_v
    port map (
            O => \N__16740\,
            I => \N__16732\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__16737\,
            I => \N__16729\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__16729\,
            I => \N__16723\
        );

    \I__3640\ : Span4Mux_v
    port map (
            O => \N__16726\,
            I => \N__16720\
        );

    \I__3639\ : Span4Mux_v
    port map (
            O => \N__16723\,
            I => \N__16717\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__16720\,
            I => \POWERLED.N_100\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__16717\,
            I => \POWERLED.N_100\
        );

    \I__3636\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__16709\,
            I => \POWERLED.count_clk_1_sqmuxa_5_0_0\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__16706\,
            I => \POWERLED.N_171_cascade_\
        );

    \I__3633\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16694\
        );

    \I__3632\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16694\
        );

    \I__3631\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16694\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__16694\,
            I => \N__16690\
        );

    \I__3629\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16687\
        );

    \I__3628\ : Span4Mux_h
    port map (
            O => \N__16690\,
            I => \N__16683\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__16687\,
            I => \N__16680\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16677\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__16683\,
            I => \POWERLED.N_163\
        );

    \I__3624\ : Odrv12
    port map (
            O => \N__16680\,
            I => \POWERLED.N_163\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__16677\,
            I => \POWERLED.N_163\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__16670\,
            I => \N__16666\
        );

    \I__3621\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16663\
        );

    \I__3620\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16660\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__16663\,
            I => \N__16655\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__16660\,
            I => \N__16655\
        );

    \I__3617\ : Span4Mux_h
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3616\ : Span4Mux_v
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3615\ : Odrv4
    port map (
            O => \N__16649\,
            I => \POWERLED.count_clk_1_sqmuxa_5_i\
        );

    \I__3614\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16637\
        );

    \I__3613\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16637\
        );

    \I__3612\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16634\
        );

    \I__3611\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16631\
        );

    \I__3610\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16626\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__16637\,
            I => \N__16623\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16634\,
            I => \N__16620\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__16631\,
            I => \N__16617\
        );

    \I__3606\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16614\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16611\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__16626\,
            I => \N__16608\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__16623\,
            I => \N__16599\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__16620\,
            I => \N__16599\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__16617\,
            I => \N__16599\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__16614\,
            I => \N__16599\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16611\,
            I => \N__16596\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__16608\,
            I => \N__16593\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__16599\,
            I => \N__16590\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__16596\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__16593\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__16590\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__16580\,
            I => \N__16576\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__16579\,
            I => \N__16571\
        );

    \I__3590\ : Span4Mux_v
    port map (
            O => \N__16576\,
            I => \N__16567\
        );

    \I__3589\ : InMux
    port map (
            O => \N__16575\,
            I => \N__16562\
        );

    \I__3588\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16562\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16571\,
            I => \N__16557\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16557\
        );

    \I__3585\ : Sp12to4
    port map (
            O => \N__16567\,
            I => \N__16554\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__16562\,
            I => \N__16551\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__16557\,
            I => \N__16548\
        );

    \I__3582\ : Odrv12
    port map (
            O => \N__16554\,
            I => rsmrst_pwrgd_signal
        );

    \I__3581\ : Odrv12
    port map (
            O => \N__16551\,
            I => rsmrst_pwrgd_signal
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__16548\,
            I => rsmrst_pwrgd_signal
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__3578\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3576\ : Span12Mux_v
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__3575\ : Odrv12
    port map (
            O => \N__16529\,
            I => \V33S_OK_c\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__16523\,
            I => \VCCST_CPU_OK_c\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__16520\,
            I => \N__16513\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16519\,
            I => \N__16510\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16505\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16505\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16500\
        );

    \I__3567\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16500\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16510\,
            I => \N__16497\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16492\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__16500\,
            I => \N__16492\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__16497\,
            I => \N__16489\
        );

    \I__3562\ : Span4Mux_s3_v
    port map (
            O => \N__16492\,
            I => \N__16486\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__16489\,
            I => \ALL_SYS_PWRGD.N_194\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__16486\,
            I => \ALL_SYS_PWRGD.N_194\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16478\,
            I => \V5S_OK_c\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__16469\,
            I => \ALL_SYS_PWRGD.m4_0_0_a3_1\
        );

    \I__3554\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__16460\,
            I => \POWERLED.dutycycle_s_2\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16450\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__16456\,
            I => \N__16447\
        );

    \I__3549\ : InMux
    port map (
            O => \N__16455\,
            I => \N__16444\
        );

    \I__3548\ : InMux
    port map (
            O => \N__16454\,
            I => \N__16441\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16453\,
            I => \N__16438\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16450\,
            I => \N__16433\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16430\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__16444\,
            I => \N__16427\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16441\,
            I => \N__16424\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16438\,
            I => \N__16421\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__16437\,
            I => \N__16418\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__16436\,
            I => \N__16414\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__16433\,
            I => \N__16411\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16430\,
            I => \N__16404\
        );

    \I__3537\ : Span12Mux_s1_h
    port map (
            O => \N__16427\,
            I => \N__16404\
        );

    \I__3536\ : Span12Mux_s7_v
    port map (
            O => \N__16424\,
            I => \N__16404\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__16421\,
            I => \N__16401\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16398\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16393\
        );

    \I__3532\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16393\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__16411\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3530\ : Odrv12
    port map (
            O => \N__16404\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__16401\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16398\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__16393\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__16382\,
            I => \POWERLED.N_84_cascade_\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__16379\,
            I => \N__16376\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16372\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16369\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16364\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__16369\,
            I => \N__16364\
        );

    \I__3520\ : Span4Mux_v
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__16361\,
            I => \POWERLED.dutycycle\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16353\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16350\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16347\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16353\,
            I => \N__16342\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16350\,
            I => \N__16342\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__16347\,
            I => \N__16338\
        );

    \I__3512\ : Span4Mux_s2_h
    port map (
            O => \N__16342\,
            I => \N__16335\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16332\
        );

    \I__3510\ : Span12Mux_s3_h
    port map (
            O => \N__16338\,
            I => \N__16329\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__16335\,
            I => \N__16326\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16332\,
            I => \POWERLED.N_119\
        );

    \I__3507\ : Odrv12
    port map (
            O => \N__16329\,
            I => \POWERLED.N_119\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__16326\,
            I => \POWERLED.N_119\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__16319\,
            I => \N__16310\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__16318\,
            I => \N__16306\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__16317\,
            I => \N__16302\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \N__16298\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__16315\,
            I => \N__16293\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__16314\,
            I => \N__16289\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__16313\,
            I => \N__16285\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16266\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16266\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16266\
        );

    \I__3495\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16266\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16266\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16266\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16266\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16266\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16251\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16251\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16251\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16251\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16251\
        );

    \I__3485\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16251\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16251\
        );

    \I__3483\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16248\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__16266\,
            I => \N__16245\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__16251\,
            I => \N__16242\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16248\,
            I => \N__16239\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__16245\,
            I => \N__16236\
        );

    \I__3478\ : Span4Mux_h
    port map (
            O => \N__16242\,
            I => \N__16233\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__16239\,
            I => \POWERLED.N_65_i\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__16236\,
            I => \POWERLED.N_65_i\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__16233\,
            I => \POWERLED.N_65_i\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__16226\,
            I => \N__16220\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16225\,
            I => \N__16216\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16210\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16207\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16202\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16202\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16216\,
            I => \N__16199\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16196\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__16214\,
            I => \N__16192\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__16213\,
            I => \N__16189\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16186\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__16207\,
            I => \N__16183\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16202\,
            I => \N__16180\
        );

    \I__3461\ : Span4Mux_h
    port map (
            O => \N__16199\,
            I => \N__16177\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16196\,
            I => \N__16174\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16167\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16167\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16167\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__16186\,
            I => \N__16160\
        );

    \I__3455\ : Span4Mux_s1_h
    port map (
            O => \N__16183\,
            I => \N__16160\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__16180\,
            I => \N__16160\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__16177\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3452\ : Odrv12
    port map (
            O => \N__16174\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16167\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__16160\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__16151\,
            I => \N__16148\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16143\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16140\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16136\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16143\,
            I => \N__16133\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__16140\,
            I => \N__16130\
        );

    \I__3443\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16127\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__16136\,
            I => \N__16124\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__16133\,
            I => \N__16118\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__16130\,
            I => \N__16115\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16110\
        );

    \I__3438\ : Span12Mux_s9_v
    port map (
            O => \N__16124\,
            I => \N__16110\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16107\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16102\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16102\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__16118\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__16115\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3432\ : Odrv12
    port map (
            O => \N__16110\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__16107\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__16102\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16091\,
            I => \N__16086\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \N__16083\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16080\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__16086\,
            I => \N__16075\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16072\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16069\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16064\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16064\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__16075\,
            I => \N__16060\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16072\,
            I => \N__16057\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__16069\,
            I => \N__16054\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__16064\,
            I => \N__16051\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16063\,
            I => \N__16048\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__16060\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__3415\ : Odrv4
    port map (
            O => \N__16057\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__16054\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__16051\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16048\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__16037\,
            I => \N__16034\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16030\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16027\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16023\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16027\,
            I => \N__16019\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__16026\,
            I => \N__16016\
        );

    \I__3405\ : Span4Mux_h
    port map (
            O => \N__16023\,
            I => \N__16010\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16007\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__16019\,
            I => \N__16004\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16016\,
            I => \N__15995\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16015\,
            I => \N__15995\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16014\,
            I => \N__15995\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16013\,
            I => \N__15995\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__16010\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__16007\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__16004\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__15995\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__15983\,
            I => \POWERLED.N_84\
        );

    \I__3392\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15973\
        );

    \I__3391\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15973\
        );

    \I__3390\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15970\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__15973\,
            I => \N__15967\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__3387\ : Span4Mux_s3_h
    port map (
            O => \N__15967\,
            I => \N__15961\
        );

    \I__3386\ : Span4Mux_s3_h
    port map (
            O => \N__15964\,
            I => \N__15958\
        );

    \I__3385\ : Span4Mux_v
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__15958\,
            I => \POWERLED.N_116\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__15955\,
            I => \POWERLED.N_116\
        );

    \I__3382\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__15947\,
            I => \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_2\
        );

    \I__3380\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__15941\,
            I => \N__15937\
        );

    \I__3378\ : InMux
    port map (
            O => \N__15940\,
            I => \N__15934\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__15937\,
            I => \POWERLED.N_197\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__15934\,
            I => \POWERLED.N_197\
        );

    \I__3375\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15923\
        );

    \I__3374\ : InMux
    port map (
            O => \N__15928\,
            I => \N__15923\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__15920\,
            I => \POWERLED.dutycycle_cnst_1_i_o2_0_a3_2_5\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__15917\,
            I => \POWERLED.N_196_cascade_\
        );

    \I__3370\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15911\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__15911\,
            I => \N__15908\
        );

    \I__3368\ : Span4Mux_s2_h
    port map (
            O => \N__15908\,
            I => \N__15904\
        );

    \I__3367\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15901\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__15904\,
            I => \POWERLED.dutycycle_s_6\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__15901\,
            I => \POWERLED.dutycycle_s_6\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__15896\,
            I => \N__15889\
        );

    \I__3363\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15883\
        );

    \I__3362\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15878\
        );

    \I__3361\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15878\
        );

    \I__3360\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15875\
        );

    \I__3359\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15872\
        );

    \I__3358\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15867\
        );

    \I__3357\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15867\
        );

    \I__3356\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15864\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__15883\,
            I => \N__15859\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__15878\,
            I => \N__15859\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__15875\,
            I => \N__15856\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__15872\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__15867\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__15864\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__15859\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__15856\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__15845\,
            I => \N__15842\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15838\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__15841\,
            I => \N__15835\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__15838\,
            I => \N__15832\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15829\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__15832\,
            I => \N__15826\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__15829\,
            I => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__15826\,
            I => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15818\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__15818\,
            I => \N__15815\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__15812\,
            I => \POWERLED.dutycycle_RNI6NI81Z0Z_5\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__15809\,
            I => \N__15805\
        );

    \I__3334\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15802\
        );

    \I__3333\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15799\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15802\,
            I => \N__15796\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__15799\,
            I => \N__15793\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__15796\,
            I => \N__15790\
        );

    \I__3329\ : Span4Mux_h
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__15790\,
            I => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__15787\,
            I => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__3324\ : Span4Mux_v
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__15773\,
            I => \POWERLED.dutycycle_RNIK4I81Z0Z_6\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15763\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__15769\,
            I => \N__15760\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__15768\,
            I => \N__15757\
        );

    \I__3319\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15753\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__15766\,
            I => \N__15749\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__15763\,
            I => \N__15744\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15741\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15738\
        );

    \I__3314\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15735\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__15753\,
            I => \N__15732\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15723\
        );

    \I__3311\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15723\
        );

    \I__3310\ : InMux
    port map (
            O => \N__15748\,
            I => \N__15723\
        );

    \I__3309\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15723\
        );

    \I__3308\ : Span4Mux_v
    port map (
            O => \N__15744\,
            I => \N__15716\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__15741\,
            I => \N__15716\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__15738\,
            I => \N__15716\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__15735\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__15732\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__15723\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__15716\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__15704\,
            I => \N__15701\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__15701\,
            I => \POWERLED.un1_dutycycle_1_axb_8\
        );

    \I__3298\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__3296\ : Span4Mux_s3_h
    port map (
            O => \N__15692\,
            I => \N__15683\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__15691\,
            I => \N__15680\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15675\
        );

    \I__3293\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15675\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__15688\,
            I => \N__15671\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__15687\,
            I => \N__15668\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15663\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__15683\,
            I => \N__15660\
        );

    \I__3288\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15657\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__15675\,
            I => \N__15654\
        );

    \I__3286\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15649\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15649\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15642\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15642\
        );

    \I__3282\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15642\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__15663\,
            I => \N__15639\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__15660\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__15657\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__15654\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15649\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__15642\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__15639\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__15626\,
            I => \N__15622\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15617\
        );

    \I__3272\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15614\
        );

    \I__3271\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15611\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15608\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15604\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15614\,
            I => \N__15598\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15611\,
            I => \N__15593\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__15608\,
            I => \N__15593\
        );

    \I__3265\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15590\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15604\,
            I => \N__15587\
        );

    \I__3263\ : InMux
    port map (
            O => \N__15603\,
            I => \N__15580\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15580\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15580\
        );

    \I__3260\ : Span4Mux_v
    port map (
            O => \N__15598\,
            I => \N__15575\
        );

    \I__3259\ : Span4Mux_v
    port map (
            O => \N__15593\,
            I => \N__15575\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__15590\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__15587\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15580\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__15575\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__15566\,
            I => \N__15562\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15555\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15552\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15547\
        );

    \I__3250\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15547\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__15559\,
            I => \N__15544\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15541\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15536\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__15552\,
            I => \N__15533\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__15547\,
            I => \N__15530\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15527\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15524\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15540\,
            I => \N__15519\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15519\
        );

    \I__3240\ : Span4Mux_s1_h
    port map (
            O => \N__15536\,
            I => \N__15512\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__15533\,
            I => \N__15512\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__15530\,
            I => \N__15512\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15527\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__15524\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__15519\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__15512\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15497\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3230\ : Odrv12
    port map (
            O => \N__15494\,
            I => \POWERLED.dutycycle_RNIEJ021Z0Z_4\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__15491\,
            I => \POWERLED.N_173_cascade_\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15485\,
            I => \N__15481\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15478\
        );

    \I__3225\ : Span4Mux_s3_h
    port map (
            O => \N__15481\,
            I => \N__15475\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15478\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__15475\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15464\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__15458\,
            I => \POWERLED.func_state_ns_0_i_o2_11_1\
        );

    \I__3217\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15452\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__15452\,
            I => \N__15448\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__15451\,
            I => \N__15445\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__15448\,
            I => \N__15442\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15439\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__15442\,
            I => \POWERLED.dutycycle_RNIFHLJZ0Z_0\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15439\,
            I => \POWERLED.dutycycle_RNIFHLJZ0Z_0\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__3208\ : Span4Mux_v
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__15425\,
            I => \POWERLED.dutycycle_RNI16B71Z0Z_5\
        );

    \I__3206\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15419\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__15419\,
            I => \N__15415\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__3203\ : Span4Mux_v
    port map (
            O => \N__15415\,
            I => \N__15409\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15412\,
            I => \POWERLED.N_126\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__15409\,
            I => \POWERLED.N_126\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__15404\,
            I => \POWERLED.N_168_cascade_\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__15401\,
            I => \POWERLED.un2_slp_s3n_2_0_2_cascade_\
        );

    \I__3198\ : SRMux
    port map (
            O => \N__15398\,
            I => \N__15393\
        );

    \I__3197\ : SRMux
    port map (
            O => \N__15397\,
            I => \N__15390\
        );

    \I__3196\ : SRMux
    port map (
            O => \N__15396\,
            I => \N__15387\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15393\,
            I => \N__15384\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15381\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__15387\,
            I => \N__15378\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__15384\,
            I => \N__15375\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__15381\,
            I => \N__15372\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__15378\,
            I => \N__15369\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__15375\,
            I => \POWERLED.count_clk_RNI95RKLZ0Z_8\
        );

    \I__3188\ : Odrv4
    port map (
            O => \N__15372\,
            I => \POWERLED.count_clk_RNI95RKLZ0Z_8\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__15369\,
            I => \POWERLED.count_clk_RNI95RKLZ0Z_8\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__15362\,
            I => \POWERLED.count_clk_RNI95RKLZ0Z_8_cascade_\
        );

    \I__3185\ : CEMux
    port map (
            O => \N__15359\,
            I => \N__15356\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__15350\,
            I => \POWERLED.N_39_1\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15344\,
            I => \POWERLED.N_167\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15341\,
            I => \bfn_9_11_0_\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \N__15327\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15322\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15317\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15317\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15306\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15306\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15306\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15306\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15306\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15303\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15298\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15298\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__15322\,
            I => \N__15291\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__15317\,
            I => \N__15291\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15306\,
            I => \N__15291\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__15303\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__15298\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__15291\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__15284\,
            I => \N__15280\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15273\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15270\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15279\,
            I => \N__15267\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__15278\,
            I => \N__15263\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15277\,
            I => \N__15258\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15276\,
            I => \N__15255\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__15273\,
            I => \N__15248\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__15270\,
            I => \N__15248\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__15267\,
            I => \N__15248\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15239\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15239\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15239\
        );

    \I__3147\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15239\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15258\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15255\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__15248\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__15239\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__15230\,
            I => \POWERLED.func_state_ns_0_i_o3_5_0_cascade_\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15224\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15224\,
            I => \POWERLED.func_state_ns_0_i_o3_6_0\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15215\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__15220\,
            I => \N__15211\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__15219\,
            I => \N__15208\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__15218\,
            I => \N__15205\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15202\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15199\
        );

    \I__3133\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15194\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15208\,
            I => \N__15191\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15188\
        );

    \I__3130\ : Span4Mux_h
    port map (
            O => \N__15202\,
            I => \N__15183\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__15199\,
            I => \N__15183\
        );

    \I__3128\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15178\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15178\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__15194\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15191\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15188\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__15183\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__15178\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__15164\,
            I => \POWERLED.func_state_ns_0_i_o3_7_0\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__15161\,
            I => \N__15154\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__15160\,
            I => \N__15150\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15159\,
            I => \N__15147\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__15158\,
            I => \N__15140\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15129\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15129\
        );

    \I__3113\ : InMux
    port map (
            O => \N__15153\,
            I => \N__15129\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15129\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15129\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15124\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15124\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15121\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15116\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15116\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__15129\,
            I => \N__15111\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15124\,
            I => \N__15111\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__15121\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__15116\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3101\ : Odrv4
    port map (
            O => \N__15111\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__15104\,
            I => \POWERLED.un1_dutycycle_1_39_0_cascade_\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__15101\,
            I => \N__15098\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15095\,
            I => \N__15092\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__15092\,
            I => \POWERLED.dutycycle_RNI34C41Z0Z_8\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__15089\,
            I => \N__15085\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__15088\,
            I => \N__15082\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15076\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15069\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15069\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15069\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15066\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__15076\,
            I => \N__15063\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15069\,
            I => \N__15060\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15066\,
            I => \N__15057\
        );

    \I__3085\ : Span4Mux_v
    port map (
            O => \N__15063\,
            I => \N__15054\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__15060\,
            I => \N__15051\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__15057\,
            I => \N__15048\
        );

    \I__3082\ : Sp12to4
    port map (
            O => \N__15054\,
            I => \N__15045\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__15051\,
            I => \POWERLED.N_78\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__15048\,
            I => \POWERLED.N_78\
        );

    \I__3079\ : Odrv12
    port map (
            O => \N__15045\,
            I => \POWERLED.N_78\
        );

    \I__3078\ : InMux
    port map (
            O => \N__15038\,
            I => \N__15035\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__15032\,
            I => \N__15028\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15025\
        );

    \I__3074\ : Span4Mux_s0_h
    port map (
            O => \N__15028\,
            I => \N__15022\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15025\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__15022\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15014\,
            I => \N__15010\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15007\
        );

    \I__3068\ : Span4Mux_s3_h
    port map (
            O => \N__15010\,
            I => \N__15004\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__15007\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__15004\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__14999\,
            I => \N__14996\
        );

    \I__3064\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14989\
        );

    \I__3062\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14986\
        );

    \I__3061\ : Span4Mux_s3_h
    port map (
            O => \N__14989\,
            I => \N__14983\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__14986\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__14983\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3058\ : InMux
    port map (
            O => \N__14978\,
            I => \POWERLED.dutycycle_cry_5\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14975\,
            I => \bfn_9_10_0_\
        );

    \I__3056\ : InMux
    port map (
            O => \N__14972\,
            I => \POWERLED.dutycycle_cry_7\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14969\,
            I => \POWERLED.dutycycle_cry_8\
        );

    \I__3054\ : InMux
    port map (
            O => \N__14966\,
            I => \POWERLED.dutycycle_cry_9\
        );

    \I__3053\ : InMux
    port map (
            O => \N__14963\,
            I => \POWERLED.dutycycle_cry_10\
        );

    \I__3052\ : InMux
    port map (
            O => \N__14960\,
            I => \POWERLED.dutycycle_cry_11\
        );

    \I__3051\ : InMux
    port map (
            O => \N__14957\,
            I => \POWERLED.dutycycle_cry_12\
        );

    \I__3050\ : InMux
    port map (
            O => \N__14954\,
            I => \POWERLED.dutycycle_cry_13\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__14951\,
            I => \N__14948\
        );

    \I__3048\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14940\
        );

    \I__3047\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14940\
        );

    \I__3046\ : IoInMux
    port map (
            O => \N__14946\,
            I => \N__14935\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__14945\,
            I => \N__14932\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14940\,
            I => \N__14928\
        );

    \I__3043\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14925\
        );

    \I__3042\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14922\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14919\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14932\,
            I => \N__14913\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14931\,
            I => \N__14913\
        );

    \I__3038\ : Span4Mux_h
    port map (
            O => \N__14928\,
            I => \N__14906\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__14925\,
            I => \N__14906\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__14922\,
            I => \N__14906\
        );

    \I__3035\ : IoSpan4Mux
    port map (
            O => \N__14919\,
            I => \N__14903\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14900\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__14913\,
            I => \N__14897\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__14906\,
            I => \N__14892\
        );

    \I__3031\ : Span4Mux_s1_h
    port map (
            O => \N__14903\,
            I => \N__14887\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__14900\,
            I => \N__14887\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__14897\,
            I => \N__14883\
        );

    \I__3028\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14880\
        );

    \I__3027\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14877\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__14892\,
            I => \N__14873\
        );

    \I__3025\ : Span4Mux_v
    port map (
            O => \N__14887\,
            I => \N__14870\
        );

    \I__3024\ : InMux
    port map (
            O => \N__14886\,
            I => \N__14867\
        );

    \I__3023\ : Sp12to4
    port map (
            O => \N__14883\,
            I => \N__14864\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__14880\,
            I => \N__14859\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__14877\,
            I => \N__14859\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14856\
        );

    \I__3019\ : Span4Mux_v
    port map (
            O => \N__14873\,
            I => \N__14852\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__14870\,
            I => \N__14847\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14847\
        );

    \I__3016\ : Span12Mux_s8_v
    port map (
            O => \N__14864\,
            I => \N__14840\
        );

    \I__3015\ : Span12Mux_s8_h
    port map (
            O => \N__14859\,
            I => \N__14840\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__14856\,
            I => \N__14840\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14837\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__14852\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__14847\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3010\ : Odrv12
    port map (
            O => \N__14840\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__14837\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3008\ : InMux
    port map (
            O => \N__14828\,
            I => \bfn_9_8_0_\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14818\
        );

    \I__3005\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14815\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__14818\,
            I => \N__14812\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__14815\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__3002\ : Odrv12
    port map (
            O => \N__14812\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__3000\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__14798\,
            I => \N__14795\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__14795\,
            I => \POWERLED.dutycycle_s_0\
        );

    \I__2996\ : InMux
    port map (
            O => \N__14792\,
            I => \POWERLED.dutycycle_cry_c_0_THRU_CO\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__14789\,
            I => \N__14786\
        );

    \I__2994\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__2992\ : Span4Mux_h
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__14777\,
            I => \POWERLED.dutycycle_s_1\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14774\,
            I => \POWERLED.dutycycle_cry_0\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14771\,
            I => \POWERLED.dutycycle_cry_1\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14768\,
            I => \POWERLED.dutycycle_cry_2\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14765\,
            I => \POWERLED.dutycycle_cry_3\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14762\,
            I => \POWERLED.dutycycle_cry_4\
        );

    \I__2985\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14754\
        );

    \I__2984\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14751\
        );

    \I__2983\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14748\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__14754\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14751\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__14748\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14741\,
            I => \POWERLED.un1_count_clk_1_cry_6\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14738\,
            I => \bfn_9_7_0_\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14731\
        );

    \I__2976\ : InMux
    port map (
            O => \N__14734\,
            I => \N__14728\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__14731\,
            I => \N__14725\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__14728\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__14725\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__2972\ : InMux
    port map (
            O => \N__14720\,
            I => \POWERLED.un1_count_clk_1_cry_8\
        );

    \I__2971\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14713\
        );

    \I__2970\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14710\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__14713\,
            I => \N__14707\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__14710\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__14707\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__2966\ : InMux
    port map (
            O => \N__14702\,
            I => \POWERLED.un1_count_clk_1_cry_9\
        );

    \I__2965\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14695\
        );

    \I__2964\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14692\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14695\,
            I => \N__14689\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__14692\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__14689\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__2960\ : InMux
    port map (
            O => \N__14684\,
            I => \POWERLED.un1_count_clk_1_cry_10\
        );

    \I__2959\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14677\
        );

    \I__2958\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14674\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__14677\,
            I => \N__14671\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__14674\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__14671\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__2954\ : InMux
    port map (
            O => \N__14666\,
            I => \POWERLED.un1_count_clk_1_cry_11\
        );

    \I__2953\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14659\
        );

    \I__2952\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14656\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__14659\,
            I => \N__14653\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__14656\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__2949\ : Odrv12
    port map (
            O => \N__14653\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__2948\ : InMux
    port map (
            O => \N__14648\,
            I => \POWERLED.un1_count_clk_1_cry_12\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__2946\ : InMux
    port map (
            O => \N__14642\,
            I => \N__14638\
        );

    \I__2945\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14635\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14638\,
            I => \N__14632\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14635\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__14632\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14627\,
            I => \POWERLED.un1_count_clk_1_cry_13\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__14624\,
            I => \POWERLED.dutycycle_1_sqmuxa_i_o6_1_5_cascade_\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__14618\,
            I => \POWERLED.dutycycle_1_sqmuxa_i_o6_1_6\
        );

    \I__2937\ : SRMux
    port map (
            O => \N__14615\,
            I => \N__14611\
        );

    \I__2936\ : SRMux
    port map (
            O => \N__14614\,
            I => \N__14608\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__14611\,
            I => \N__14605\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__14608\,
            I => \N__14601\
        );

    \I__2933\ : Span4Mux_v
    port map (
            O => \N__14605\,
            I => \N__14598\
        );

    \I__2932\ : SRMux
    port map (
            O => \N__14604\,
            I => \N__14595\
        );

    \I__2931\ : Span4Mux_v
    port map (
            O => \N__14601\,
            I => \N__14587\
        );

    \I__2930\ : Span4Mux_s2_v
    port map (
            O => \N__14598\,
            I => \N__14587\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14595\,
            I => \N__14587\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14584\
        );

    \I__2927\ : Sp12to4
    port map (
            O => \N__14587\,
            I => \N__14581\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14578\
        );

    \I__2925\ : Odrv12
    port map (
            O => \N__14581\,
            I => \ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__14578\,
            I => \ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0\
        );

    \I__2923\ : CEMux
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__14570\,
            I => \N__14567\
        );

    \I__2921\ : Odrv12
    port map (
            O => \N__14567\,
            I => \ALL_SYS_PWRGD.N_39_5\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14560\
        );

    \I__2919\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14557\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__14560\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__14557\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14548\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14545\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__14548\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__14545\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14540\,
            I => \POWERLED.un1_count_clk_1_cry_0\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14530\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14530\
        );

    \I__2909\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14527\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__14530\,
            I => \N__14524\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14527\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__14524\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__2905\ : InMux
    port map (
            O => \N__14519\,
            I => \POWERLED.un1_count_clk_1_cry_1\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14511\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14506\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14506\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__14511\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__14506\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14501\,
            I => \POWERLED.un1_count_clk_1_cry_2\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14491\
        );

    \I__2897\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14491\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14496\,
            I => \N__14488\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__14491\,
            I => \N__14485\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14488\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__14485\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14480\,
            I => \POWERLED.un1_count_clk_1_cry_3\
        );

    \I__2891\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14473\
        );

    \I__2890\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14470\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__14473\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__14470\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__2887\ : InMux
    port map (
            O => \N__14465\,
            I => \POWERLED.un1_count_clk_1_cry_4\
        );

    \I__2886\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14457\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14454\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14451\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14457\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14454\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__14451\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14444\,
            I => \POWERLED.un1_count_clk_1_cry_5\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14438\,
            I => \ALL_SYS_PWRGD.un4_count_10\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__14435\,
            I => \ALL_SYS_PWRGD.un4_count_9_cascade_\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__14432\,
            I => \N__14429\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14422\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14422\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14419\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__14422\,
            I => \ALL_SYS_PWRGD.N_1_i\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__14419\,
            I => \ALL_SYS_PWRGD.N_1_i\
        );

    \I__2870\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14410\
        );

    \I__2869\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14407\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__14410\,
            I => \ALL_SYS_PWRGD.countZ0Z_7\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__14407\,
            I => \ALL_SYS_PWRGD.countZ0Z_7\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14398\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14401\,
            I => \N__14395\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14398\,
            I => \ALL_SYS_PWRGD.countZ0Z_6\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__14395\,
            I => \ALL_SYS_PWRGD.countZ0Z_6\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__14390\,
            I => \N__14386\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14383\,
            I => \ALL_SYS_PWRGD.countZ0Z_8\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__14380\,
            I => \ALL_SYS_PWRGD.countZ0Z_8\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14371\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14368\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__14371\,
            I => \ALL_SYS_PWRGD.countZ0Z_4\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__14368\,
            I => \ALL_SYS_PWRGD.countZ0Z_4\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14363\,
            I => \N__14360\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14360\,
            I => \ALL_SYS_PWRGD.un4_count_8\
        );

    \I__2851\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14353\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14350\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14353\,
            I => \ALL_SYS_PWRGD.countZ0Z_14\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__14350\,
            I => \ALL_SYS_PWRGD.countZ0Z_14\
        );

    \I__2847\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14341\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14338\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__14341\,
            I => \ALL_SYS_PWRGD.countZ0Z_13\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14338\,
            I => \ALL_SYS_PWRGD.countZ0Z_13\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__14333\,
            I => \N__14329\
        );

    \I__2842\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14326\
        );

    \I__2841\ : InMux
    port map (
            O => \N__14329\,
            I => \N__14323\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14326\,
            I => \ALL_SYS_PWRGD.countZ0Z_15\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__14323\,
            I => \ALL_SYS_PWRGD.countZ0Z_15\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14314\
        );

    \I__2837\ : InMux
    port map (
            O => \N__14317\,
            I => \N__14311\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__14314\,
            I => \ALL_SYS_PWRGD.countZ0Z_12\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14311\,
            I => \ALL_SYS_PWRGD.countZ0Z_12\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14303\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14303\,
            I => \N__14300\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__14300\,
            I => \ALL_SYS_PWRGD.un4_count_11\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14294\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14294\,
            I => \POWERLED.func_state_ns_0_i_o2_10_1\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14291\,
            I => \N__14288\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14288\,
            I => \POWERLED.func_state_ns_0_i_o2_9_1\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14282\,
            I => \POWERLED.func_state_ns_0_i_o2_8_1\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14276\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__14276\,
            I => \POWERLED.un1_func_state11_2_i_o6_0_2\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__14273\,
            I => \POWERLED.N_100_cascade_\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__14270\,
            I => \N__14267\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__14264\,
            I => \POWERLED.dutycycle_RNI75MGZ0Z_15\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14258\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__14258\,
            I => \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa\
        );

    \I__2817\ : IoInMux
    port map (
            O => \N__14255\,
            I => \N__14251\
        );

    \I__2816\ : IoInMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14244\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14241\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__14247\,
            I => \N__14236\
        );

    \I__2812\ : Span4Mux_s3_v
    port map (
            O => \N__14244\,
            I => \N__14233\
        );

    \I__2811\ : IoSpan4Mux
    port map (
            O => \N__14241\,
            I => \N__14230\
        );

    \I__2810\ : IoInMux
    port map (
            O => \N__14240\,
            I => \N__14227\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14222\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14222\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__14233\,
            I => \N__14219\
        );

    \I__2806\ : Span4Mux_s1_v
    port map (
            O => \N__14230\,
            I => \N__14216\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14213\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__14222\,
            I => \N__14210\
        );

    \I__2803\ : Span4Mux_v
    port map (
            O => \N__14219\,
            I => \N__14207\
        );

    \I__2802\ : Span4Mux_h
    port map (
            O => \N__14216\,
            I => \N__14202\
        );

    \I__2801\ : Span4Mux_s1_v
    port map (
            O => \N__14213\,
            I => \N__14202\
        );

    \I__2800\ : Span12Mux_s8_h
    port map (
            O => \N__14210\,
            I => \N__14199\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__14207\,
            I => \VCCIN_EN_c\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__14202\,
            I => \VCCIN_EN_c\
        );

    \I__2797\ : Odrv12
    port map (
            O => \N__14199\,
            I => \VCCIN_EN_c\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__14192\,
            I => \ALL_SYS_PWRGD.N_44_cascade_\
        );

    \I__2795\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14185\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14182\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14185\,
            I => \ALL_SYS_PWRGD.countZ0Z_5\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__14182\,
            I => \ALL_SYS_PWRGD.countZ0Z_5\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14173\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14170\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14173\,
            I => \ALL_SYS_PWRGD.countZ0Z_3\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__14170\,
            I => \ALL_SYS_PWRGD.countZ0Z_3\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__14165\,
            I => \N__14161\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14155\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__14158\,
            I => \ALL_SYS_PWRGD.countZ0Z_11\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14155\,
            I => \ALL_SYS_PWRGD.countZ0Z_11\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14146\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14143\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14146\,
            I => \ALL_SYS_PWRGD.countZ0Z_2\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__14143\,
            I => \ALL_SYS_PWRGD.countZ0Z_2\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14123\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14134\,
            I => \N__14123\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14133\,
            I => \N__14123\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14120\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14115\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14115\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__14123\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__14120\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14115\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14096\
        );

    \I__2767\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14096\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14106\,
            I => \N__14096\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14093\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14088\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14088\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__14096\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__14093\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__14088\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__14081\,
            I => \N__14077\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14074\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14071\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__14074\,
            I => \ALL_SYS_PWRGD.un1_curr_state10_0\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__14071\,
            I => \ALL_SYS_PWRGD.un1_curr_state10_0\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14066\,
            I => \N__14062\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14065\,
            I => \N__14059\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__14062\,
            I => \ALL_SYS_PWRGD.countZ0Z_9\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14059\,
            I => \ALL_SYS_PWRGD.countZ0Z_9\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14050\
        );

    \I__2749\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14047\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14050\,
            I => \ALL_SYS_PWRGD.countZ0Z_0\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14047\,
            I => \ALL_SYS_PWRGD.countZ0Z_0\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__14042\,
            I => \N__14038\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__14035\,
            I => \ALL_SYS_PWRGD.countZ0Z_1\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__14032\,
            I => \ALL_SYS_PWRGD.countZ0Z_1\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14023\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14020\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14023\,
            I => \ALL_SYS_PWRGD.countZ0Z_10\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14020\,
            I => \ALL_SYS_PWRGD.countZ0Z_10\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14012\,
            I => \POWERLED.dutycycle_RNIE4FLZ0Z_9\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__14003\,
            I => \POWERLED.N_165\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13996\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__13999\,
            I => \N__13993\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2729\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__13990\,
            I => \POWERLED.dutycycle_RNI2V0PZ0Z_10\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__13987\,
            I => \POWERLED.dutycycle_RNI2V0PZ0Z_10\
        );

    \I__2726\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__13979\,
            I => \POWERLED.dutycycle_RNI712I1Z0Z_15\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \POWERLED.un1_dutycycle_1_44_0_cascade_\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__2722\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__13967\,
            I => \POWERLED.dutycycle_RNIF3561Z0Z_9\
        );

    \I__2720\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__13961\,
            I => \POWERLED.dutycycle_RNI53MGZ0Z_14\
        );

    \I__2718\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13955\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__13955\,
            I => \POWERLED.dutycycle_RNI31MGZ0Z_12\
        );

    \I__2716\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13949\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__13949\,
            I => \POWERLED.dutycycle_RNI73C11Z0Z_15\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2713\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__13940\,
            I => \POWERLED.dutycycle_RNI31MG_0Z0Z_12\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \N__13933\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__13936\,
            I => \N__13930\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13922\
        );

    \I__2708\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13922\
        );

    \I__2707\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13922\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__13922\,
            I => \POWERLED.dutycycle_fastZ0Z_6\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__2704\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13913\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__13907\,
            I => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__13904\,
            I => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6_cascade_\
        );

    \I__2699\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__13895\,
            I => \POWERLED.dutycycle_RNIJL1R1Z0Z_6\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__13886\,
            I => \POWERLED.dutycycle_RNIC8C11Z0Z_15\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2692\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__13877\,
            I => \POWERLED.dutycycle_RNIO18NZ0Z_9\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__13874\,
            I => \POWERLED.dutycycle_RNIO18NZ0Z_9_cascade_\
        );

    \I__2689\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__13868\,
            I => \POWERLED.dutycycle_RNIQ09G1Z0Z_10\
        );

    \I__2687\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__13862\,
            I => \POWERLED.dutycycle_RNIB1FLZ0Z_8\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__2684\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__13853\,
            I => \POWERLED.dutycycle_RNI84C11Z0Z_14\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__13850\,
            I => \N__13846\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13843\
        );

    \I__2680\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13840\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__13843\,
            I => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__13840\,
            I => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\
        );

    \I__2677\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__13832\,
            I => \POWERLED.dutycycle_RNIJNBA1Z0Z_6\
        );

    \I__2675\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13825\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__13825\,
            I => \N__13819\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__13822\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__13819\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__2670\ : InMux
    port map (
            O => \N__13814\,
            I => \POWERLED.un1_count_off_1_cry_12\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13807\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__13807\,
            I => \N__13801\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13804\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__13801\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13796\,
            I => \POWERLED.un1_count_off_1_cry_13\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13793\,
            I => \bfn_8_9_0_\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__13790\,
            I => \N__13787\
        );

    \I__2661\ : InMux
    port map (
            O => \N__13787\,
            I => \N__13783\
        );

    \I__2660\ : InMux
    port map (
            O => \N__13786\,
            I => \N__13780\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__13783\,
            I => \N__13777\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__13780\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__13777\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__2656\ : CEMux
    port map (
            O => \N__13772\,
            I => \N__13769\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__13769\,
            I => \N__13766\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__13766\,
            I => \N__13763\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__13763\,
            I => \POWERLED.N_39_0\
        );

    \I__2652\ : SRMux
    port map (
            O => \N__13760\,
            I => \N__13756\
        );

    \I__2651\ : SRMux
    port map (
            O => \N__13759\,
            I => \N__13752\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__13756\,
            I => \N__13749\
        );

    \I__2649\ : SRMux
    port map (
            O => \N__13755\,
            I => \N__13746\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13752\,
            I => \N__13743\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__13749\,
            I => \N__13740\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__13746\,
            I => \N__13737\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__13743\,
            I => \N__13734\
        );

    \I__2644\ : Span4Mux_s3_h
    port map (
            O => \N__13740\,
            I => \N__13731\
        );

    \I__2643\ : Span12Mux_s6_h
    port map (
            O => \N__13737\,
            I => \N__13728\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__13734\,
            I => \POWERLED.func_state_RNI9L40BZ0Z_0\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__13731\,
            I => \POWERLED.func_state_RNI9L40BZ0Z_0\
        );

    \I__2640\ : Odrv12
    port map (
            O => \N__13728\,
            I => \POWERLED.func_state_RNI9L40BZ0Z_0\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__13721\,
            I => \N__13718\
        );

    \I__2638\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13715\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__13715\,
            I => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__13712\,
            I => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6_cascade_\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__13706\,
            I => \POWERLED.dutycycle_RNIQAI81Z0Z_4\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13700\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__13700\,
            I => \POWERLED.dutycycle_RNIOQLJZ0Z_4\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13697\,
            I => \POWERLED.un1_count_off_1_cry_4\
        );

    \I__2630\ : InMux
    port map (
            O => \N__13694\,
            I => \POWERLED.un1_count_off_1_cry_5\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__13691\,
            I => \N__13687\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13684\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13681\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__13684\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__13681\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13676\,
            I => \POWERLED.un1_count_off_1_cry_6\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13669\
        );

    \I__2622\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13666\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13669\,
            I => \N__13663\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__13666\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__13663\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13658\,
            I => \bfn_8_8_0_\
        );

    \I__2617\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13651\
        );

    \I__2616\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13648\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__13651\,
            I => \N__13645\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13648\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__13645\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__2612\ : InMux
    port map (
            O => \N__13640\,
            I => \POWERLED.un1_count_off_1_cry_8\
        );

    \I__2611\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13633\
        );

    \I__2610\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13630\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13633\,
            I => \N__13627\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__13630\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__13627\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__2606\ : InMux
    port map (
            O => \N__13622\,
            I => \POWERLED.un1_count_off_1_cry_9\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__13619\,
            I => \N__13616\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13612\
        );

    \I__2603\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13609\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13612\,
            I => \N__13606\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__13609\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__13606\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13601\,
            I => \POWERLED.un1_count_off_1_cry_10\
        );

    \I__2598\ : InMux
    port map (
            O => \N__13598\,
            I => \N__13594\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13597\,
            I => \N__13591\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__13594\,
            I => \N__13588\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__13591\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__13588\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13583\,
            I => \POWERLED.un1_count_off_1_cry_11\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__13580\,
            I => \POWERLED.dutycycle_1_sqmuxa_i_o6_0_0_cascade_\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__13577\,
            I => \N__13573\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13576\,
            I => \N__13570\
        );

    \I__2589\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13567\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__13570\,
            I => \POWERLED.N_68_i\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13567\,
            I => \POWERLED.N_68_i\
        );

    \I__2586\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13558\
        );

    \I__2585\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13555\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__13558\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__13555\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2582\ : InMux
    port map (
            O => \N__13550\,
            I => \POWERLED.un1_count_off_1_cry_0\
        );

    \I__2581\ : InMux
    port map (
            O => \N__13547\,
            I => \POWERLED.un1_count_off_1_cry_1\
        );

    \I__2580\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13540\
        );

    \I__2579\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13537\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__13540\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__13537\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2576\ : InMux
    port map (
            O => \N__13532\,
            I => \POWERLED.un1_count_off_1_cry_2\
        );

    \I__2575\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13525\
        );

    \I__2574\ : InMux
    port map (
            O => \N__13528\,
            I => \N__13522\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__13525\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__13522\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13517\,
            I => \POWERLED.un1_count_off_1_cry_3\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13514\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_9\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13511\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_10\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13508\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_11\
        );

    \I__2567\ : InMux
    port map (
            O => \N__13505\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_12\
        );

    \I__2566\ : InMux
    port map (
            O => \N__13502\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_13\
        );

    \I__2565\ : InMux
    port map (
            O => \N__13499\,
            I => \bfn_8_5_0_\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13496\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_0\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13493\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_1\
        );

    \I__2562\ : InMux
    port map (
            O => \N__13490\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_2\
        );

    \I__2561\ : InMux
    port map (
            O => \N__13487\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_3\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13484\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_4\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13481\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_5\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13478\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_6\
        );

    \I__2557\ : InMux
    port map (
            O => \N__13475\,
            I => \bfn_8_4_0_\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13472\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_8\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13463\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__2552\ : InMux
    port map (
            O => \N__13460\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__2550\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13451\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__13445\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13442\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2544\ : InMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13433\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2540\ : Span4Mux_h
    port map (
            O => \N__13424\,
            I => \N__13421\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__13421\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13418\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__13415\,
            I => \N__13412\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13405\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13405\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13402\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13405\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__13402\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13392\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13396\,
            I => \N__13389\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13395\,
            I => \N__13386\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13392\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13389\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13386\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__13379\,
            I => \N__13376\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13373\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__2522\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13367\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13367\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13364\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13361\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__13358\,
            I => \N__13355\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13352\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13352\,
            I => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13344\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13339\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13339\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__13344\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13339\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__13334\,
            I => \N__13331\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__13328\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13325\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__13322\,
            I => \N__13319\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13316\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13316\,
            I => \POWERLED.mult1_un47_sum_axb_4\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13313\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13304\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13304\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13301\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__13292\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_5\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13289\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13286\,
            I => \POWERLED.mult1_un47_sum_cry_6\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__13283\,
            I => \POWERLED.mult1_un54_sum_s_8_cascade_\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__13280\,
            I => \N__13276\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__13279\,
            I => \N__13272\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13265\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13275\,
            I => \N__13265\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13265\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13265\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__13262\,
            I => \N__13258\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13253\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13253\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__13250\,
            I => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13247\,
            I => \N__13243\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13240\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13237\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13240\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__13237\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13226\,
            I => \POWERLED.un1_dutycycle_1_i_28\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13217\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13217\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__2470\ : InMux
    port map (
            O => \N__13214\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13211\,
            I => \bfn_7_13_0_\
        );

    \I__2468\ : InMux
    port map (
            O => \N__13208\,
            I => \POWERLED.CO2\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13205\,
            I => \N__13202\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__13202\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__13199\,
            I => \N__13195\
        );

    \I__2464\ : InMux
    port map (
            O => \N__13198\,
            I => \N__13190\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13190\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__13190\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \N__13183\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__13186\,
            I => \N__13179\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13169\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13169\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13169\
        );

    \I__2456\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13169\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__13169\,
            I => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13157\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13157\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13164\,
            I => \N__13157\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__13157\,
            I => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13149\
        );

    \I__2449\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13144\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13144\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13149\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__13144\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__2445\ : IoInMux
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13136\,
            I => \N__13133\
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__13133\,
            I => \VPP_VDDQ_un2_vpp_en_0_i\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__13130\,
            I => \N__13127\
        );

    \I__2441\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13124\,
            I => \POWERLED.un1_dutycycle_1_i_29\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13118\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__13118\,
            I => \N__13114\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13111\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__13114\,
            I => \N__13108\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13105\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__13108\,
            I => \N__13102\
        );

    \I__2433\ : Odrv12
    port map (
            O => \N__13105\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__13102\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13097\,
            I => \bfn_7_12_0_\
        );

    \I__2430\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13091\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__13091\,
            I => \N__13087\
        );

    \I__2428\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13084\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__13087\,
            I => \N__13081\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__13084\,
            I => \N__13078\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__13081\,
            I => \N__13075\
        );

    \I__2424\ : Odrv12
    port map (
            O => \N__13078\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__13075\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2422\ : InMux
    port map (
            O => \N__13070\,
            I => \POWERLED.un1_dutycycle_1_cry_8\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13064\,
            I => \N__13060\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13057\
        );

    \I__2418\ : Span4Mux_h
    port map (
            O => \N__13060\,
            I => \N__13052\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__13057\,
            I => \N__13052\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__13052\,
            I => \N__13049\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__13049\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13046\,
            I => \POWERLED.un1_dutycycle_1_cry_9\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13040\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__13040\,
            I => \N__13036\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13033\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__13036\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13033\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13028\,
            I => \POWERLED.un1_dutycycle_1_cry_10\
        );

    \I__2407\ : InMux
    port map (
            O => \N__13025\,
            I => \N__13021\
        );

    \I__2406\ : InMux
    port map (
            O => \N__13024\,
            I => \N__13018\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__13021\,
            I => \N__13015\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__13018\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__13015\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13010\,
            I => \POWERLED.un1_dutycycle_1_cry_11\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13007\,
            I => \POWERLED.un1_dutycycle_1_cry_12\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13004\,
            I => \POWERLED.un1_dutycycle_1_cry_13\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13001\,
            I => \POWERLED.un1_dutycycle_1_cry_14\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12994\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12991\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__12994\,
            I => \N__12986\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__12991\,
            I => \N__12986\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__12986\,
            I => \POWERLED.un1_dutycycle_1_axb_0\
        );

    \I__2393\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12980\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__12980\,
            I => \POWERLED.un1_dutycycle_1_axb_1\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__2390\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12970\
        );

    \I__2389\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12967\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__12970\,
            I => \N__12964\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__12967\,
            I => \N__12959\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__12964\,
            I => \N__12959\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__12959\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__2384\ : InMux
    port map (
            O => \N__12956\,
            I => \POWERLED.un1_dutycycle_1_cry_0\
        );

    \I__2383\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12950\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__12950\,
            I => \N__12946\
        );

    \I__2381\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12943\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__12946\,
            I => \N__12940\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__12943\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__12940\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__2377\ : InMux
    port map (
            O => \N__12935\,
            I => \POWERLED.un1_dutycycle_1_cry_1\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__12932\,
            I => \N__12929\
        );

    \I__2375\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12925\
        );

    \I__2374\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12922\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__12925\,
            I => \N__12919\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__12922\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__12919\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12914\,
            I => \POWERLED.un1_dutycycle_1_cry_2\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12904\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12907\,
            I => \N__12901\
        );

    \I__2366\ : Span4Mux_v
    port map (
            O => \N__12904\,
            I => \N__12898\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__12901\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__12898\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__2363\ : InMux
    port map (
            O => \N__12893\,
            I => \POWERLED.un1_dutycycle_1_cry_3\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12890\,
            I => \N__12886\
        );

    \I__2361\ : InMux
    port map (
            O => \N__12889\,
            I => \N__12883\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12886\,
            I => \N__12878\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__12883\,
            I => \N__12878\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__12878\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__2357\ : InMux
    port map (
            O => \N__12875\,
            I => \POWERLED.un1_dutycycle_1_cry_4\
        );

    \I__2356\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12868\
        );

    \I__2355\ : InMux
    port map (
            O => \N__12871\,
            I => \N__12865\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__12868\,
            I => \N__12860\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__12865\,
            I => \N__12860\
        );

    \I__2352\ : Odrv12
    port map (
            O => \N__12860\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12857\,
            I => \POWERLED.un1_dutycycle_1_cry_5\
        );

    \I__2350\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12850\
        );

    \I__2349\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12847\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__12850\,
            I => \N__12842\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12842\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__12839\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__2344\ : InMux
    port map (
            O => \N__12836\,
            I => \POWERLED.un1_dutycycle_1_cry_6\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__12830\,
            I => \N__12826\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__12829\,
            I => \N__12823\
        );

    \I__2340\ : Span4Mux_s2_h
    port map (
            O => \N__12826\,
            I => \N__12819\
        );

    \I__2339\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12814\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12814\
        );

    \I__2337\ : Span4Mux_h
    port map (
            O => \N__12819\,
            I => \N__12809\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__12814\,
            I => \N__12806\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12803\
        );

    \I__2334\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12800\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__12809\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__12806\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__12803\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__12800\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__12791\,
            I => \N__12787\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12784\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12781\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12784\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__12781\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__2324\ : InMux
    port map (
            O => \N__12776\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__2323\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__12767\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__12764\,
            I => \N__12760\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__12763\,
            I => \N__12756\
        );

    \I__2318\ : InMux
    port map (
            O => \N__12760\,
            I => \N__12749\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12749\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12749\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__12749\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__12740\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12737\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__12734\,
            I => \N__12731\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__12725\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12722\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \N__12712\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__12718\,
            I => \N__12708\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__12717\,
            I => \N__12705\
        );

    \I__2302\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12702\
        );

    \I__2301\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12697\
        );

    \I__2300\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12697\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12694\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12708\,
            I => \N__12689\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12689\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__12702\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__12697\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12694\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__12689\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__12680\,
            I => \POWERLED.mult1_un110_sum_s_8_cascade_\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12671\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__12671\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__2288\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__2286\ : Span4Mux_s2_h
    port map (
            O => \N__12662\,
            I => \N__12659\
        );

    \I__2285\ : Span4Mux_h
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__12656\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12650\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__12650\,
            I => \N__12647\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__12647\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12641\,
            I => \POWERLED.mult1_un117_sum_axb_7_l_fx\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12635\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12635\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12628\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12625\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12628\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12625\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__2272\ : InMux
    port map (
            O => \N__12620\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12614\,
            I => \N__12611\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__12611\,
            I => \N__12608\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__12608\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12605\,
            I => \N__12602\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12602\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12599\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__12596\,
            I => \N__12593\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12590\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12590\,
            I => \N__12587\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__12587\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__12584\,
            I => \N__12581\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12581\,
            I => \N__12578\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12578\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__2257\ : InMux
    port map (
            O => \N__12575\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12569\,
            I => \N__12566\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__12566\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12563\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__12560\,
            I => \N__12557\
        );

    \I__2251\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12554\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__12554\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12551\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12545\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__2246\ : InMux
    port map (
            O => \N__12542\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__12539\,
            I => \N__12534\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12530\
        );

    \I__2243\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12525\
        );

    \I__2242\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12525\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12522\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__12530\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__12525\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__12522\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12509\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12509\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12506\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__2233\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__12500\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__12497\,
            I => \N__12493\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__12496\,
            I => \N__12489\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12482\
        );

    \I__2228\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12482\
        );

    \I__2227\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12482\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__12482\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12479\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__12470\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__2221\ : InMux
    port map (
            O => \N__12467\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12461\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__2217\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12452\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__12452\,
            I => \POWERLED.mult1_un117_sum_axb_4_l_fx\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12445\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12442\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__12445\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12442\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12433\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12430\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__12433\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12430\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__12425\,
            I => \N__12421\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12418\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12415\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12418\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12415\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12406\
        );

    \I__2201\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12403\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__12406\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12403\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12395\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12395\,
            I => \RSMRST_PWRGD.un4_count_10\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12392\,
            I => \N__12388\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12391\,
            I => \N__12385\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__12388\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__12385\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12376\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12373\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12376\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12373\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__12368\,
            I => \N__12364\
        );

    \I__2187\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12361\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12358\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12361\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__12358\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12349\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12346\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12349\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__12346\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12338\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__12338\,
            I => \RSMRST_PWRGD.un4_count_9\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12324\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12324\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12333\,
            I => \N__12324\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12319\
        );

    \I__2173\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12319\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12324\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12319\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__12314\,
            I => \N__12307\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__12313\,
            I => \N__12304\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12299\
        );

    \I__2167\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12299\
        );

    \I__2166\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12292\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12292\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12292\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12299\,
            I => \N__12289\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12292\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__12289\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__2159\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12277\
        );

    \I__2158\ : InMux
    port map (
            O => \N__12280\,
            I => \N__12274\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__12277\,
            I => \N__12271\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__12274\,
            I => \RSMRST_PWRGD.N_51_i\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__12271\,
            I => \RSMRST_PWRGD.N_51_i\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12262\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12259\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12262\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__12259\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12250\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12247\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12250\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12247\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__12242\,
            I => \N__12238\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12235\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12232\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12235\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12232\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__2141\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12223\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12220\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__12223\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12220\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__2137\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__12209\,
            I => \RSMRST_PWRGD.un4_count_11\
        );

    \I__2134\ : SRMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12203\,
            I => \N__12200\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__12200\,
            I => \N__12196\
        );

    \I__2131\ : SRMux
    port map (
            O => \N__12199\,
            I => \N__12193\
        );

    \I__2130\ : Span4Mux_s2_v
    port map (
            O => \N__12196\,
            I => \N__12186\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12193\,
            I => \N__12186\
        );

    \I__2128\ : SRMux
    port map (
            O => \N__12192\,
            I => \N__12183\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12180\
        );

    \I__2126\ : Sp12to4
    port map (
            O => \N__12186\,
            I => \N__12177\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__12183\,
            I => \N__12174\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__12180\,
            I => \N__12171\
        );

    \I__2123\ : Odrv12
    port map (
            O => \N__12177\,
            I => \RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0\
        );

    \I__2122\ : Odrv12
    port map (
            O => \N__12174\,
            I => \RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__12171\,
            I => \RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0\
        );

    \I__2120\ : CEMux
    port map (
            O => \N__12164\,
            I => \N__12161\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12161\,
            I => \N__12158\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__12158\,
            I => \RSMRST_PWRGD.N_39_3\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12152\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__12152\,
            I => \N__12147\
        );

    \I__2115\ : IoInMux
    port map (
            O => \N__12151\,
            I => \N__12144\
        );

    \I__2114\ : IoInMux
    port map (
            O => \N__12150\,
            I => \N__12141\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__12147\,
            I => \N__12138\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12135\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12141\,
            I => \N__12132\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__12138\,
            I => \N__12129\
        );

    \I__2109\ : IoSpan4Mux
    port map (
            O => \N__12135\,
            I => \N__12126\
        );

    \I__2108\ : Span12Mux_s8_h
    port map (
            O => \N__12132\,
            I => \N__12123\
        );

    \I__2107\ : IoSpan4Mux
    port map (
            O => \N__12129\,
            I => \N__12118\
        );

    \I__2106\ : IoSpan4Mux
    port map (
            O => \N__12126\,
            I => \N__12118\
        );

    \I__2105\ : Odrv12
    port map (
            O => \N__12123\,
            I => \V5A_EN_c\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__12118\,
            I => \V5A_EN_c\
        );

    \I__2103\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__12110\,
            I => \N__12107\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__12101\,
            I => \V5A_OK_c\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__2095\ : Sp12to4
    port map (
            O => \N__12089\,
            I => \N__12086\
        );

    \I__2094\ : Span12Mux_v
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__2093\ : Odrv12
    port map (
            O => \N__12083\,
            I => \V33A_OK_c\
        );

    \I__2092\ : IoInMux
    port map (
            O => \N__12080\,
            I => \N__12077\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__2090\ : IoSpan4Mux
    port map (
            O => \N__12074\,
            I => \N__12070\
        );

    \I__2089\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12067\
        );

    \I__2088\ : Span4Mux_s1_h
    port map (
            O => \N__12070\,
            I => \N__12064\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__12067\,
            I => \N__12061\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__12064\,
            I => \N__12056\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__12061\,
            I => \N__12056\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__2083\ : Span4Mux_h
    port map (
            O => \N__12053\,
            I => \N__12050\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__12050\,
            I => \V1P8A_OK_c\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12044\,
            I => \N__12041\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__12041\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__2078\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12035\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__12035\,
            I => \N__12032\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__12032\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12029\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__12026\,
            I => \N__12021\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12025\,
            I => \N__12018\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12024\,
            I => \N__12013\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12013\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12018\,
            I => \N__12009\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__12013\,
            I => \N__12005\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12012\,
            I => \N__12002\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__12009\,
            I => \N__11999\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12008\,
            I => \N__11996\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__12005\,
            I => \N__11991\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12002\,
            I => \N__11991\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__11999\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__11996\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__11991\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__2060\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11980\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11977\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__11980\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__11977\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__2056\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11968\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__11968\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__11965\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__11960\,
            I => \N__11956\
        );

    \I__2051\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11953\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11950\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__11953\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__11950\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__2047\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11941\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11938\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__11941\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11938\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__11933\,
            I => \RSMRST_PWRGD.un4_count_8_cascade_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__11927\,
            I => \RSMRST_PWRGD.N_1_i\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__11924\,
            I => \RSMRST_PWRGD.N_1_i_cascade_\
        );

    \I__2039\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__11918\,
            I => \RSMRST_PWRGD.N_85\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__11915\,
            I => \RSMRST_PWRGD.N_85_cascade_\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__11912\,
            I => \N__11908\
        );

    \I__2035\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11902\
        );

    \I__2034\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11899\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11894\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11906\,
            I => \N__11894\
        );

    \I__2031\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11891\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__11902\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__11899\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__11894\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__11891\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2026\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11871\
        );

    \I__2025\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11871\
        );

    \I__2024\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11866\
        );

    \I__2023\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11866\
        );

    \I__2022\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11861\
        );

    \I__2021\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11861\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11858\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__11871\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__11866\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__11861\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__11858\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__11849\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__11846\,
            I => \N__11843\
        );

    \I__2013\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11840\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__11840\,
            I => \N__11837\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__11837\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__2010\ : InMux
    port map (
            O => \N__11834\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__2009\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__11825\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11822\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__11819\,
            I => \N__11816\
        );

    \I__2004\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11813\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__11810\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__2001\ : InMux
    port map (
            O => \N__11807\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__2000\ : InMux
    port map (
            O => \N__11804\,
            I => \N__11801\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__11801\,
            I => \N__11798\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__11798\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__1997\ : InMux
    port map (
            O => \N__11795\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__1996\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11789\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__11786\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11783\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__1991\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__11774\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__1989\ : InMux
    port map (
            O => \N__11771\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__1988\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__11765\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__1986\ : InMux
    port map (
            O => \N__11762\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1984\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__11753\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11750\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__1981\ : InMux
    port map (
            O => \N__11747\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__11744\,
            I => \N__11739\
        );

    \I__1979\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11735\
        );

    \I__1978\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11730\
        );

    \I__1977\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11730\
        );

    \I__1976\ : InMux
    port map (
            O => \N__11738\,
            I => \N__11727\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__11735\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11730\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__11727\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__11720\,
            I => \POWERLED.mult1_un68_sum_s_8_cascade_\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__11717\,
            I => \N__11713\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__11716\,
            I => \N__11709\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11702\
        );

    \I__1968\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11702\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11702\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__11702\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__11699\,
            I => \N__11695\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__11698\,
            I => \N__11691\
        );

    \I__1963\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11684\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11684\
        );

    \I__1961\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11684\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__11684\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__1959\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11678\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__11678\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__11675\,
            I => \N__11671\
        );

    \I__1956\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11668\
        );

    \I__1955\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11665\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__11668\,
            I => \N__11660\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__11665\,
            I => \N__11660\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__11657\,
            I => \VPP_VDDQ.N_32_i\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__11648\,
            I => \POWERLED.count_off_0_sqmuxa\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11639\
        );

    \I__1945\ : Span4Mux_s2_h
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__11633\,
            I => \POWERLED.un1_count_2_8\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__11630\,
            I => \POWERLED.func_state_RNI9L40BZ0Z_0_cascade_\
        );

    \I__1941\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__1939\ : Odrv12
    port map (
            O => \N__11621\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11614\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__11617\,
            I => \N__11610\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11614\,
            I => \N__11605\
        );

    \I__1935\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11600\
        );

    \I__1934\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11600\
        );

    \I__1933\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11597\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11594\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__11605\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__11600\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11597\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11594\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11582\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__1925\ : Odrv12
    port map (
            O => \N__11579\,
            I => \POWERLED.un1_count_2_7\
        );

    \I__1924\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__11573\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__11564\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__1919\ : InMux
    port map (
            O => \N__11561\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11555\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__11555\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11552\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11543\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__11543\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__11534\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11531\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11525\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11525\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__1905\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__11516\,
            I => \N__11513\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__11513\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__1902\ : InMux
    port map (
            O => \N__11510\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11501\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__11492\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__1895\ : InMux
    port map (
            O => \N__11489\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__1894\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__11483\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__11480\,
            I => \N__11476\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__11479\,
            I => \N__11472\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11465\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11465\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11465\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11465\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11459\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11459\,
            I => \N__11456\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__11456\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__1883\ : InMux
    port map (
            O => \N__11453\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__11450\,
            I => \N__11447\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11444\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11441\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11434\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__11437\,
            I => \N__11430\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11434\,
            I => \N__11427\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11422\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11422\
        );

    \I__1873\ : Span4Mux_s3_h
    port map (
            O => \N__11427\,
            I => \N__11415\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__11422\,
            I => \N__11415\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11421\,
            I => \N__11412\
        );

    \I__1870\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11409\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__11415\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__11412\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__11409\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__11402\,
            I => \N__11398\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__11401\,
            I => \N__11394\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11387\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11387\
        );

    \I__1862\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11387\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__11384\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__11372\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__11363\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11360\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11357\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11354\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11351\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11348\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11345\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1845\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__11333\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11330\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__11327\,
            I => \POWERLED.mult1_un96_sum_s_8_cascade_\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11320\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11317\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__11320\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__11317\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11308\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11308\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11305\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11300\,
            I => \N__11296\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__11293\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11290\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11281\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11281\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__11278\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11269\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11266\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11269\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11266\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__1819\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11257\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11254\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__11257\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11254\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11239\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11236\
        );

    \I__1811\ : Span4Mux_h
    port map (
            O => \N__11239\,
            I => \N__11233\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11236\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__11233\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11224\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11221\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__11224\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11221\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__11216\,
            I => \VPP_VDDQ.un6_count_11_cascade_\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11210\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__11210\,
            I => \VPP_VDDQ.un6_count_8\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11203\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11200\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__11203\,
            I => \N__11197\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11200\,
            I => \N__11194\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__11197\,
            I => \N__11189\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__11194\,
            I => \N__11189\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__11189\,
            I => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11186\,
            I => \N__11182\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11185\,
            I => \N__11179\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__11182\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__11179\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11170\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11167\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11170\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11167\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11162\,
            I => \N__11158\
        );

    \I__1785\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11152\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11155\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11152\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11143\
        );

    \I__1780\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11140\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11143\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11140\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__11132\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11125\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11128\,
            I => \N__11122\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__11125\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__11122\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11113\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11113\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__11110\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__11105\,
            I => \N__11101\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11098\
        );

    \I__1765\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11095\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11098\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11095\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11086\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11086\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__11083\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__11075\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__1756\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__1754\ : Span4Mux_s2_h
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__11060\,
            I => \POWERLED.un1_count_2_10\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11057\,
            I => \bfn_6_5_0_\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11054\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__11045\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11042\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__11036\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11033\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11026\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__11029\,
            I => \N__11022\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__11026\,
            I => \N__11017\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11012\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11012\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11021\,
            I => \N__11009\
        );

    \I__1736\ : InMux
    port map (
            O => \N__11020\,
            I => \N__11006\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__11017\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11012\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11009\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__11006\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__10997\,
            I => \N__10994\
        );

    \I__1730\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10991\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__10991\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__1728\ : InMux
    port map (
            O => \N__10988\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__1727\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__10982\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__10979\,
            I => \N__10975\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__10978\,
            I => \N__10971\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10964\
        );

    \I__1722\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10964\
        );

    \I__1721\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10964\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__10964\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__1719\ : InMux
    port map (
            O => \N__10961\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1717\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10952\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__10952\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10949\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__1714\ : InMux
    port map (
            O => \N__10946\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__1713\ : InMux
    port map (
            O => \N__10943\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__1712\ : InMux
    port map (
            O => \N__10940\,
            I => \bfn_6_4_0_\
        );

    \I__1711\ : InMux
    port map (
            O => \N__10937\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__1710\ : InMux
    port map (
            O => \N__10934\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__1709\ : InMux
    port map (
            O => \N__10931\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__1708\ : InMux
    port map (
            O => \N__10928\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10925\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10922\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__10919\,
            I => \VPP_VDDQ.G_110_0_cascade_\
        );

    \I__1704\ : SRMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10908\
        );

    \I__1702\ : SRMux
    port map (
            O => \N__10912\,
            I => \N__10905\
        );

    \I__1701\ : SRMux
    port map (
            O => \N__10911\,
            I => \N__10901\
        );

    \I__1700\ : Span4Mux_h
    port map (
            O => \N__10908\,
            I => \N__10896\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10896\
        );

    \I__1698\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10893\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__10901\,
            I => \N__10890\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__10896\,
            I => \N__10887\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10884\
        );

    \I__1694\ : Odrv12
    port map (
            O => \N__10890\,
            I => \VPP_VDDQ.curr_state_RNIQINR7Z0Z_0\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__10887\,
            I => \VPP_VDDQ.curr_state_RNIQINR7Z0Z_0\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__10884\,
            I => \VPP_VDDQ.curr_state_RNIQINR7Z0Z_0\
        );

    \I__1691\ : InMux
    port map (
            O => \N__10877\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__1690\ : InMux
    port map (
            O => \N__10874\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__1689\ : InMux
    port map (
            O => \N__10871\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__1688\ : InMux
    port map (
            O => \N__10868\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10865\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__10856\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10853\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__10850\,
            I => \N__10847\
        );

    \I__1681\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__10841\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10838\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__1677\ : InMux
    port map (
            O => \N__10835\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__1676\ : CEMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__10826\,
            I => \VPP_VDDQ.N_39_2\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__1671\ : Odrv12
    port map (
            O => \N__10817\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__1670\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__10808\,
            I => \POWERLED.un1_count_2_14\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__10805\,
            I => \N__10801\
        );

    \I__1666\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10795\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10795\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__10800\,
            I => \N__10792\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10787\
        );

    \I__1662\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10784\
        );

    \I__1661\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10781\
        );

    \I__1660\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10778\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__10787\,
            I => \N__10773\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10773\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__10781\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__10778\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__10773\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1653\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__1651\ : Odrv12
    port map (
            O => \N__10757\,
            I => \POWERLED.un1_count_2_13\
        );

    \I__1650\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10751\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__10751\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10748\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10745\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__1646\ : InMux
    port map (
            O => \N__10742\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__1645\ : InMux
    port map (
            O => \N__10739\,
            I => \bfn_5_9_0_\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__10724\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__1639\ : InMux
    port map (
            O => \N__10721\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__1638\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10715\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__10712\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__1635\ : InMux
    port map (
            O => \N__10709\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1633\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__10697\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__1630\ : InMux
    port map (
            O => \N__10694\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10691\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10688\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__1627\ : InMux
    port map (
            O => \N__10685\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10682\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__1625\ : InMux
    port map (
            O => \N__10679\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10676\,
            I => \bfn_5_8_0_\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10673\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10670\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__1621\ : InMux
    port map (
            O => \N__10667\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10658\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10655\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__10649\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10646\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__1613\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10639\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__10642\,
            I => \N__10635\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__10639\,
            I => \N__10631\
        );

    \I__1610\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10626\
        );

    \I__1609\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10626\
        );

    \I__1608\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10623\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__10631\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10626\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10623\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__10610\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10607\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__10601\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__10598\,
            I => \N__10594\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__10597\,
            I => \N__10590\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10583\
        );

    \I__1595\ : InMux
    port map (
            O => \N__10593\,
            I => \N__10583\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10583\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__10583\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10580\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10571\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__10571\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__1588\ : InMux
    port map (
            O => \N__10568\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10565\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10562\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10555\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10552\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__10555\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__10552\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10543\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__10543\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__10540\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__10535\,
            I => \N__10531\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10528\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10525\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10528\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__10525\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1572\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10516\
        );

    \I__1571\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10513\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__10516\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__10513\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10505\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__10502\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10495\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__10495\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10492\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10483\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10480\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10483\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__10480\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__10475\,
            I => \N__10471\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10468\
        );

    \I__1555\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10465\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__10468\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__10465\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1552\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10456\
        );

    \I__1551\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10456\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__10453\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__10442\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10435\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10432\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10435\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__10432\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10423\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10420\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10423\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10420\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__10415\,
            I => \N__10411\
        );

    \I__1536\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10408\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10405\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10408\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10405\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10396\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10393\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10396\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__10393\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__10382\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10375\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10372\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__10375\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10372\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10363\
        );

    \I__1520\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10360\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__10363\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__10360\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__10355\,
            I => \N__10351\
        );

    \I__1516\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10348\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10345\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10348\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10345\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10336\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10333\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10336\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10333\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1506\ : Odrv12
    port map (
            O => \N__10322\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10315\
        );

    \I__1504\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10312\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__10315\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10312\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10303\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10300\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10303\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10300\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__10295\,
            I => \N__10291\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10288\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10285\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__10288\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10285\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10276\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10273\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__10276\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10273\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__10262\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10259\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1482\ : Span4Mux_s2_v
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__10247\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10244\,
            I => \bfn_5_3_0_\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10238\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__10238\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__10235\,
            I => \N__10231\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10226\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10223\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10218\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10218\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10226\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10223\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10218\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10206\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10201\
        );

    \I__1467\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10201\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10206\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10201\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__10196\,
            I => \N__10192\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10189\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10186\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10189\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10186\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10176\
        );

    \I__1458\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10171\
        );

    \I__1457\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10171\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10176\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10171\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10163\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10157\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__1450\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10148\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10148\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__1447\ : Span4Mux_h
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__10142\,
            I => \N__10132\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10123\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10123\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10123\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10123\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10116\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10116\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10116\
        );

    \I__1438\ : Span4Mux_v
    port map (
            O => \N__10132\,
            I => \N__10113\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__10123\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10116\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__10113\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10101\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10096\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10104\,
            I => \N__10096\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10101\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10096\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10091\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__10088\,
            I => \N__10083\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10080\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10075\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10075\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__10080\,
            I => \N__10071\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10075\,
            I => \N__10068\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10065\
        );

    \I__1421\ : Span4Mux_s3_h
    port map (
            O => \N__10071\,
            I => \N__10062\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__10068\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__10065\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__10062\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__10055\,
            I => \POWERLED.mult1_un145_sum_s_8_cascade_\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__1414\ : Span4Mux_s3_h
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__10043\,
            I => \POWERLED.un1_count_2_3\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__1410\ : Span4Mux_s3_h
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__10031\,
            I => \POWERLED.un1_count_2_15\
        );

    \I__1408\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10024\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10020\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10017\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10014\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__10011\
        );

    \I__1403\ : Span4Mux_s3_h
    port map (
            O => \N__10017\,
            I => \N__10008\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__10014\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__10011\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__10008\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__10001\,
            I => \N__9997\
        );

    \I__1398\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9994\
        );

    \I__1397\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9986\
        );

    \I__1395\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9981\
        );

    \I__1394\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9981\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9978\
        );

    \I__1392\ : Span4Mux_s3_h
    port map (
            O => \N__9986\,
            I => \N__9975\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__9981\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__9978\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__9975\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1388\ : SRMux
    port map (
            O => \N__9968\,
            I => \N__9964\
        );

    \I__1387\ : SRMux
    port map (
            O => \N__9967\,
            I => \N__9961\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__9964\,
            I => \N__9955\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9952\
        );

    \I__1384\ : SRMux
    port map (
            O => \N__9960\,
            I => \N__9949\
        );

    \I__1383\ : SRMux
    port map (
            O => \N__9959\,
            I => \N__9946\
        );

    \I__1382\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9943\
        );

    \I__1381\ : Span4Mux_h
    port map (
            O => \N__9955\,
            I => \N__9938\
        );

    \I__1380\ : Span4Mux_s2_v
    port map (
            O => \N__9952\,
            I => \N__9938\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__9949\,
            I => \N__9931\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__9946\,
            I => \N__9931\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__9943\,
            I => \N__9931\
        );

    \I__1376\ : Odrv4
    port map (
            O => \N__9938\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__9931\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1374\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__9923\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1371\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__9914\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__1369\ : InMux
    port map (
            O => \N__9911\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__9908\,
            I => \POWERLED.mult1_un138_sum_s_8_cascade_\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1366\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__9896\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__1363\ : InMux
    port map (
            O => \N__9893\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__1361\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9884\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__1359\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9878\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__9875\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9872\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__1355\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__9866\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__9863\,
            I => \N__9860\
        );

    \I__1352\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__9854\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9851\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__1348\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__9845\,
            I => \N__9841\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__9844\,
            I => \N__9837\
        );

    \I__1345\ : Span4Mux_s3_h
    port map (
            O => \N__9841\,
            I => \N__9833\
        );

    \I__1344\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9828\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9828\
        );

    \I__1342\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9825\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__9833\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__9828\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__9825\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9812\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__9812\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9803\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__9803\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__1332\ : InMux
    port map (
            O => \N__9800\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__1331\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__9794\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__9791\,
            I => \N__9787\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__9790\,
            I => \N__9783\
        );

    \I__1327\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9776\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9786\,
            I => \N__9776\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9776\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__9776\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__1323\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__9770\,
            I => \N__9767\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__9767\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9764\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__9755\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__1316\ : InMux
    port map (
            O => \N__9752\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9749\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__9746\,
            I => \N__9743\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__9740\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9737\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9731\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9731\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9728\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__1307\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9721\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__9724\,
            I => \N__9717\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__9721\,
            I => \N__9712\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9707\
        );

    \I__1303\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9707\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9704\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9701\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__9712\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9707\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__9704\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__9701\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__1295\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__9686\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9683\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__9677\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__9674\,
            I => \N__9670\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__9673\,
            I => \N__9666\
        );

    \I__1288\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9659\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9659\
        );

    \I__1286\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9659\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__9659\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9656\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__9653\,
            I => \POWERLED.mult1_un82_sum_s_8_cascade_\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__9650\,
            I => \N__9646\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__9649\,
            I => \N__9642\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9635\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9635\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9635\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9635\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__9629\,
            I => \N__9626\
        );

    \I__1274\ : Span4Mux_s3_h
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__9623\,
            I => \POWERLED.un1_count_2_11\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9617\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9614\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9611\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9608\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9605\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9602\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__1264\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9590\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9590\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__9590\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__1260\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9578\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9578\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__9578\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__9575\,
            I => \N__9571\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9566\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9566\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9566\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__1253\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9557\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9557\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9554\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9551\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9548\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9545\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9542\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9539\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__1244\ : InMux
    port map (
            O => \N__9536\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9533\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9530\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9527\,
            I => \bfn_4_6_0_\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9524\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9521\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9518\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9515\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__1236\ : InMux
    port map (
            O => \N__9512\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__1235\ : InMux
    port map (
            O => \N__9509\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9506\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9503\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9500\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9497\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9494\,
            I => \bfn_4_5_0_\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9491\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9488\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9485\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__1226\ : InMux
    port map (
            O => \N__9482\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__9479\,
            I => \N__9474\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9471\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9466\
        );

    \I__1222\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9466\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9471\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__9466\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1219\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__9458\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9455\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__1216\ : InMux
    port map (
            O => \N__9452\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__1215\ : InMux
    port map (
            O => \N__9449\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9446\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9443\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9440\,
            I => \bfn_4_4_0_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9437\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9434\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9431\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9428\,
            I => \bfn_2_16_0_\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__9425\,
            I => \N__9421\
        );

    \I__1206\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9417\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9413\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9410\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9407\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9404\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__9413\,
            I => \N__9401\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__9410\,
            I => \N__9396\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__9407\,
            I => \N__9396\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9404\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1197\ : Odrv12
    port map (
            O => \N__9401\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__9396\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1195\ : CEMux
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__9386\,
            I => \N__9383\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__9383\,
            I => \POWERLED.N_39_6\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9375\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9370\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9370\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9375\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9370\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9362\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9359\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9351\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9346\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9346\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9351\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9346\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9338\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9335\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9328\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9324\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9328\,
            I => \N__9321\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9317\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9324\,
            I => \N__9312\
        );

    \I__1171\ : Span4Mux_s1_h
    port map (
            O => \N__9321\,
            I => \N__9312\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9309\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9317\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__9312\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__9309\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9302\,
            I => \bfn_2_15_0_\
        );

    \I__1165\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__9296\,
            I => \N__9292\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9289\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__9292\,
            I => \N__9282\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9289\,
            I => \N__9282\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9288\,
            I => \N__9279\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9276\
        );

    \I__1158\ : Span4Mux_s1_h
    port map (
            O => \N__9282\,
            I => \N__9273\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__9279\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9276\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__9273\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9266\,
            I => \POWERLED.un1_count_1_cry_9\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9259\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9254\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9259\,
            I => \N__9251\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9248\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9245\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__9254\,
            I => \N__9240\
        );

    \I__1147\ : Span4Mux_s1_h
    port map (
            O => \N__9251\,
            I => \N__9240\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9248\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9245\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__9240\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9233\,
            I => \POWERLED.un1_count_1_cry_10\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9226\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9221\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9226\,
            I => \N__9218\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9215\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9212\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9207\
        );

    \I__1136\ : Span4Mux_s1_h
    port map (
            O => \N__9218\,
            I => \N__9207\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__9215\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9212\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__9207\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9200\,
            I => \POWERLED.un1_count_1_cry_11\
        );

    \I__1131\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9193\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9189\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9185\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9182\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9179\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9176\
        );

    \I__1125\ : Span4Mux_s2_h
    port map (
            O => \N__9185\,
            I => \N__9173\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9182\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__9179\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__9176\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__9173\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9164\,
            I => \POWERLED.un1_count_1_cry_12\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9157\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9152\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__9157\,
            I => \N__9149\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9146\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9143\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9152\,
            I => \N__9138\
        );

    \I__1113\ : Span4Mux_s1_h
    port map (
            O => \N__9149\,
            I => \N__9138\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9146\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9143\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__9138\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9131\,
            I => \POWERLED.un1_count_1_cry_13\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9125\,
            I => \N__9120\
        );

    \I__1106\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9116\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9113\
        );

    \I__1104\ : Span4Mux_h
    port map (
            O => \N__9120\,
            I => \N__9110\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9107\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__9116\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9113\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__9110\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9107\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1098\ : IoInMux
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__1096\ : Span4Mux_s3_v
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__9089\,
            I => \PWRBTN_LED_c\
        );

    \I__1094\ : CEMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__9077\,
            I => \POWERLED.pwm_out_RNOZ0\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9070\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9066\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9070\,
            I => \N__9063\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9059\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9054\
        );

    \I__1085\ : Span4Mux_s1_h
    port map (
            O => \N__9063\,
            I => \N__9054\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9051\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__9059\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__9054\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9051\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9044\,
            I => \POWERLED.un1_count_1_cry_1\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9037\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9033\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__9037\,
            I => \N__9030\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9026\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__9033\,
            I => \N__9021\
        );

    \I__1074\ : Span4Mux_s1_h
    port map (
            O => \N__9030\,
            I => \N__9021\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9018\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__9026\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__9021\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9018\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9011\,
            I => \POWERLED.un1_count_1_cry_2\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9008\,
            I => \N__9004\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9000\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9004\,
            I => \N__8997\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8993\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8988\
        );

    \I__1063\ : Span4Mux_s1_h
    port map (
            O => \N__8997\,
            I => \N__8988\
        );

    \I__1062\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8985\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__8993\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__8988\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__8985\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1058\ : InMux
    port map (
            O => \N__8978\,
            I => \POWERLED.un1_count_1_cry_3\
        );

    \I__1057\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8971\
        );

    \I__1056\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8966\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__8971\,
            I => \N__8963\
        );

    \I__1054\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8960\
        );

    \I__1053\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8957\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8952\
        );

    \I__1051\ : Span4Mux_s2_h
    port map (
            O => \N__8963\,
            I => \N__8952\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__8960\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__8957\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__8952\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1047\ : InMux
    port map (
            O => \N__8945\,
            I => \POWERLED.un1_count_1_cry_4\
        );

    \I__1046\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8938\
        );

    \I__1045\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8933\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8938\,
            I => \N__8930\
        );

    \I__1043\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8927\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8924\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__8933\,
            I => \N__8919\
        );

    \I__1040\ : Span4Mux_s1_h
    port map (
            O => \N__8930\,
            I => \N__8919\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__8927\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__8924\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__8919\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1036\ : InMux
    port map (
            O => \N__8912\,
            I => \POWERLED.un1_count_1_cry_5\
        );

    \I__1035\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8904\
        );

    \I__1034\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8901\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__8907\,
            I => \N__8897\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8904\,
            I => \N__8892\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__8901\,
            I => \N__8892\
        );

    \I__1030\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8889\
        );

    \I__1029\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8886\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__8892\,
            I => \N__8883\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__8889\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__8886\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__8883\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8876\,
            I => \POWERLED.un1_count_1_cry_6\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8869\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__8869\,
            I => \N__8862\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__8866\,
            I => \N__8858\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8855\
        );

    \I__1018\ : Span4Mux_s2_h
    port map (
            O => \N__8862\,
            I => \N__8852\
        );

    \I__1017\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8849\
        );

    \I__1016\ : Span4Mux_s1_h
    port map (
            O => \N__8858\,
            I => \N__8846\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__8855\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__8852\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__8849\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__8846\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1011\ : InMux
    port map (
            O => \N__8837\,
            I => \POWERLED.un1_count_1_cry_7\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__8834\,
            I => \N__8830\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__8833\,
            I => \N__8826\
        );

    \I__1008\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8819\
        );

    \I__1007\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8819\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8819\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__8819\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__1004\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__8813\,
            I => \POWERLED.g0_0_4\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__8810\,
            I => \POWERLED.g0_0_7_cascade_\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__1000\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__8801\,
            I => \POWERLED.un1_countlt6_0\
        );

    \I__998\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__8795\,
            I => \POWERLED.g0_0_5\
        );

    \I__996\ : IoInMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__994\ : Span4Mux_s1_v
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__8780\,
            I => \tmp_RNIRH3P\
        );

    \I__991\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8773\
        );

    \I__990\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8770\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__8773\,
            I => \POWERLED.un1_count_2_cry_15_THRU_CO\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__8770\,
            I => \POWERLED.un1_count_2_cry_15_THRU_CO\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__8765\,
            I => \tmp_RNIRH3P_cascade_\
        );

    \I__986\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__8759\,
            I => \POWERLED.un1_count_0\
        );

    \I__984\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8750\
        );

    \I__983\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8750\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8750\,
            I => \COUNTER.tmp_i\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__8747\,
            I => \N__8743\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__8746\,
            I => \N__8739\
        );

    \I__979\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8732\
        );

    \I__978\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8732\
        );

    \I__977\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8732\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__8732\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__8729\,
            I => \POWERLED.mult1_un159_sum_s_7_cascade_\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__973\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__8720\,
            I => \POWERLED.un1_count_2_1\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__970\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8711\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__968\ : InMux
    port map (
            O => \N__8708\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__967\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8702\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__965\ : InMux
    port map (
            O => \N__8699\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__963\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__8690\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__961\ : InMux
    port map (
            O => \N__8687\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__960\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__8681\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__958\ : InMux
    port map (
            O => \N__8678\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__956\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__8669\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__954\ : InMux
    port map (
            O => \N__8666\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__953\ : InMux
    port map (
            O => \N__8663\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__952\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8656\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__8659\,
            I => \N__8652\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__8656\,
            I => \N__8648\
        );

    \I__949\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8643\
        );

    \I__948\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8643\
        );

    \I__947\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8640\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__8648\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__8643\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__8640\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__8633\,
            I => \POWERLED.mult1_un152_sum_s_8_cascade_\
        );

    \I__942\ : InMux
    port map (
            O => \N__8630\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__940\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8621\,
            I => \POWERLED.un1_count_2_0\
        );

    \I__938\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8615\,
            I => \POWERLED.un1_count_2_5\
        );

    \I__936\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__8606\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__932\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8597\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__930\ : InMux
    port map (
            O => \N__8594\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__928\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__8585\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__926\ : InMux
    port map (
            O => \N__8582\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__925\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__8576\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__923\ : InMux
    port map (
            O => \N__8573\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__922\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__8567\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__920\ : InMux
    port map (
            O => \N__8564\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__918\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__8555\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__916\ : InMux
    port map (
            O => \N__8552\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__915\ : InMux
    port map (
            O => \N__8549\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__8546\,
            I => \N__8542\
        );

    \I__913\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8537\
        );

    \I__912\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8530\
        );

    \I__911\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8530\
        );

    \I__910\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8530\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8537\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8530\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__907\ : InMux
    port map (
            O => \N__8525\,
            I => \bfn_2_8_0_\
        );

    \I__906\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8518\
        );

    \I__905\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__8518\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8515\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__902\ : CEMux
    port map (
            O => \N__8510\,
            I => \N__8507\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__900\ : Span4Mux_v
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__8501\,
            I => \PCH_PWRGD.N_39_4\
        );

    \I__898\ : SRMux
    port map (
            O => \N__8498\,
            I => \N__8494\
        );

    \I__897\ : SRMux
    port map (
            O => \N__8497\,
            I => \N__8490\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8487\
        );

    \I__895\ : SRMux
    port map (
            O => \N__8493\,
            I => \N__8484\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8481\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__8487\,
            I => \N__8476\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8476\
        );

    \I__891\ : Odrv12
    port map (
            O => \N__8481\,
            I => \PCH_PWRGD.curr_state_RNICTB05Z0Z_0\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__8476\,
            I => \PCH_PWRGD.curr_state_RNICTB05Z0Z_0\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__8471\,
            I => \N__8467\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \N__8463\
        );

    \I__887\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8456\
        );

    \I__886\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8456\
        );

    \I__885\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8456\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8456\,
            I => \G_386\
        );

    \I__883\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8449\
        );

    \I__882\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8446\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8449\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8446\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__879\ : InMux
    port map (
            O => \N__8441\,
            I => \PCH_PWRGD.un1_count_1_cry_5\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__8438\,
            I => \N__8434\
        );

    \I__877\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8431\
        );

    \I__876\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8431\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__8428\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__873\ : InMux
    port map (
            O => \N__8423\,
            I => \PCH_PWRGD.un1_count_1_cry_6\
        );

    \I__872\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8416\
        );

    \I__871\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8413\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8416\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__8413\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__868\ : InMux
    port map (
            O => \N__8408\,
            I => \bfn_2_7_0_\
        );

    \I__867\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8401\
        );

    \I__866\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8398\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__8401\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8398\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__863\ : InMux
    port map (
            O => \N__8393\,
            I => \PCH_PWRGD.un1_count_1_cry_8\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__8390\,
            I => \N__8386\
        );

    \I__861\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8383\
        );

    \I__860\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8380\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8383\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8380\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__857\ : InMux
    port map (
            O => \N__8375\,
            I => \PCH_PWRGD.un1_count_1_cry_9\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__8372\,
            I => \N__8368\
        );

    \I__855\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8365\
        );

    \I__854\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8362\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__8365\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8362\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__851\ : InMux
    port map (
            O => \N__8357\,
            I => \PCH_PWRGD.un1_count_1_cry_10\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__8354\,
            I => \N__8350\
        );

    \I__849\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8347\
        );

    \I__848\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8344\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__8347\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8344\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__845\ : InMux
    port map (
            O => \N__8339\,
            I => \PCH_PWRGD.un1_count_1_cry_11\
        );

    \I__844\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8332\
        );

    \I__843\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8329\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8332\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8329\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__840\ : InMux
    port map (
            O => \N__8324\,
            I => \PCH_PWRGD.un1_count_1_cry_12\
        );

    \I__839\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8317\
        );

    \I__838\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8314\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8317\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8314\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__835\ : InMux
    port map (
            O => \N__8309\,
            I => \PCH_PWRGD.un1_count_1_cry_13\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__8306\,
            I => \PCH_PWRGD.N_3_i_cascade_\
        );

    \I__833\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8296\
        );

    \I__832\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8296\
        );

    \I__831\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8293\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8296\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8293\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__828\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8285\,
            I => \PCH_PWRGD.un1_curr_state_0_sqmuxa_0\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__8282\,
            I => \N__8277\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8281\,
            I => \N__8274\
        );

    \I__824\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8265\
        );

    \I__823\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8265\
        );

    \I__822\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8265\
        );

    \I__821\ : InMux
    port map (
            O => \N__8273\,
            I => \N__8260\
        );

    \I__820\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8260\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8265\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8260\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__817\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8249\
        );

    \I__816\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8249\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__814\ : IoSpan4Mux
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__8243\,
            I => \VR_READY_VCCIN_c\
        );

    \I__812\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8229\
        );

    \I__811\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8229\
        );

    \I__810\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8229\
        );

    \I__809\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8224\
        );

    \I__808\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8224\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8229\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8224\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__805\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8215\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__8218\,
            I => \N__8212\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__802\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__8209\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8206\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__799\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8197\
        );

    \I__798\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8194\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8197\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8194\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__795\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8185\
        );

    \I__794\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8182\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8185\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8182\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__791\ : InMux
    port map (
            O => \N__8177\,
            I => \PCH_PWRGD.un1_count_1_cry_0\
        );

    \I__790\ : InMux
    port map (
            O => \N__8174\,
            I => \N__8170\
        );

    \I__789\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8170\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__8167\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__786\ : InMux
    port map (
            O => \N__8162\,
            I => \PCH_PWRGD.un1_count_1_cry_1\
        );

    \I__785\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8155\
        );

    \I__784\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8152\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8155\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__8152\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__781\ : InMux
    port map (
            O => \N__8147\,
            I => \PCH_PWRGD.un1_count_1_cry_2\
        );

    \I__780\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8140\
        );

    \I__779\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__8140\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8137\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__776\ : InMux
    port map (
            O => \N__8132\,
            I => \PCH_PWRGD.un1_count_1_cry_3\
        );

    \I__775\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8125\
        );

    \I__774\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8122\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8125\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8122\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__771\ : InMux
    port map (
            O => \N__8117\,
            I => \PCH_PWRGD.un1_count_1_cry_4\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \POWERLED.un1_countlto15_4_cascade_\
        );

    \I__769\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__8108\,
            I => \POWERLED.un1_countlto15_7\
        );

    \I__767\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8102\,
            I => \POWERLED.count_RNIOVT24Z0Z_11\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__8099\,
            I => \POWERLED.count_RNIOVT24Z0Z_11_cascade_\
        );

    \I__764\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8093\,
            I => \POWERLED.un1_countlt6\
        );

    \I__762\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__760\ : Span4Mux_s3_v
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__8081\,
            I => \VPP_OK_c\
        );

    \I__758\ : IoInMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__8072\,
            I => \VDDQ_EN_c\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__8069\,
            I => \PCH_PWRGD.curr_state_RNICTB05Z0Z_0_cascade_\
        );

    \I__754\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8057\
        );

    \I__753\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8057\
        );

    \I__752\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8057\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8057\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__750\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8051\,
            I => \POWERLED.count_i_13\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__747\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8042\,
            I => \POWERLED.count_i_14\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__744\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__8033\,
            I => \POWERLED.count_i_15\
        );

    \I__742\ : InMux
    port map (
            O => \N__8030\,
            I => \bfn_1_12_0_\
        );

    \I__741\ : IoInMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8024\,
            I => \VCCST_EN_c_i\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__8021\,
            I => \POWERLED.un1_countlto15_5_cascade_\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__737\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__8009\,
            I => \POWERLED.count_i_5\
        );

    \I__734\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8003\,
            I => \POWERLED.un1_count_2_6\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__731\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7994\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__7994\,
            I => \POWERLED.count_i_6\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__728\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__7982\,
            I => \POWERLED.count_i_7\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__724\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7973\,
            I => \POWERLED.count_i_8\
        );

    \I__722\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__7964\,
            I => \POWERLED.un1_count_2_9\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__718\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__7955\,
            I => \POWERLED.count_i_9\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__715\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__7946\,
            I => \POWERLED.count_i_10\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__712\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__7937\,
            I => \POWERLED.count_i_11\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__709\ : InMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__7925\,
            I => \POWERLED.un1_count_2_12\
        );

    \I__706\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__7919\,
            I => \POWERLED.count_i_12\
        );

    \I__704\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__7913\,
            I => \POWERLED.count_i_0_0\
        );

    \I__702\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__7907\,
            I => \POWERLED.count_i_1\
        );

    \I__700\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__7901\,
            I => \POWERLED.un1_count_2_2\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__697\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__7892\,
            I => \POWERLED.count_i_2\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__694\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__7883\,
            I => \POWERLED.count_i_3\
        );

    \I__692\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__7877\,
            I => \POWERLED.un1_count_2_4\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__689\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__7868\,
            I => \POWERLED.count_i_4\
        );

    \I__687\ : IoInMux
    port map (
            O => \N__7865\,
            I => \N__7862\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7859\
        );

    \I__685\ : Span4Mux_s3_h
    port map (
            O => \N__7859\,
            I => \N__7856\
        );

    \I__684\ : Span4Mux_h
    port map (
            O => \N__7856\,
            I => \N__7852\
        );

    \I__683\ : IoInMux
    port map (
            O => \N__7855\,
            I => \N__7849\
        );

    \I__682\ : Span4Mux_h
    port map (
            O => \N__7852\,
            I => \N__7846\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7849\,
            I => \N__7843\
        );

    \I__680\ : Sp12to4
    port map (
            O => \N__7846\,
            I => \N__7840\
        );

    \I__679\ : Span4Mux_s0_h
    port map (
            O => \N__7843\,
            I => \N__7837\
        );

    \I__678\ : Odrv12
    port map (
            O => \N__7840\,
            I => \PCH_PWROK_c\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__7837\,
            I => \PCH_PWROK_c\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__7832\,
            I => \PCH_PWRGD.un4_count_9_cascade_\
        );

    \I__675\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__7826\,
            I => \PCH_PWRGD.un4_count_11\
        );

    \I__673\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__7820\,
            I => \PCH_PWRGD.un4_count_8\
        );

    \I__671\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__7814\,
            I => \PCH_PWRGD.un4_count_10\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.dutycycle_cry_6\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.dutycycle_cry_14\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_1_cry_8\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.un4_counter_7\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_2_cry_7\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_2_cry_15\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_1_cry_7\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_1_cry_15\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_off_1_cry_7\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_off_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_1_cry_7\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALL_SYS_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_5_0_\
        );

    \COUNTER.tmp_RNIRH3P_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8792\,
            GLOBALBUFFEROUTPUT => \N_39_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PCH_PWRGD.pch_pwrok_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8240\,
            in1 => \N__8064\,
            in2 => \_gnd_net_\,
            in3 => \N__8280\,
            lcout => \PCH_PWROK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18188\,
            ce => \N__17664\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000110010"
        )
    port map (
            in0 => \N__8066\,
            in1 => \N__8239\,
            in2 => \N__8282\,
            in3 => \N__8303\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18188\,
            ce => \N__17664\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100000001000"
        )
    port map (
            in0 => \N__8065\,
            in1 => \N__8238\,
            in2 => \N__8281\,
            in3 => \N__8302\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18188\,
            ce => \N__17664\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIESHJ_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8452\,
            in1 => \N__8173\,
            in2 => \N__8390\,
            in3 => \N__8188\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7829\,
            in1 => \N__7817\,
            in2 => \N__7832\,
            in3 => \N__7823\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI7J2B_3_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8128\,
            in1 => \N__8143\,
            in2 => \N__8438\,
            in3 => \N__8158\,
            lcout => \PCH_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8320\,
            in1 => \N__8335\,
            in2 => \N__8354\,
            in3 => \N__8521\,
            lcout => \PCH_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIN5IJ_0_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8404\,
            in1 => \N__8200\,
            in2 => \N__8372\,
            in3 => \N__8419\,
            lcout => \PCH_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10643\,
            lcout => \POWERLED.un1_count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8660\,
            lcout => \POWERLED.un1_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11438\,
            lcout => \POWERLED.un1_count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12833\,
            lcout => \POWERLED.un1_count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16455\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9848\,
            lcout => \POWERLED.un1_count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_0_c_inv_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7916\,
            in2 => \N__8627\,
            in3 => \N__10000\,
            lcout => \POWERLED.count_i_0_0\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \POWERLED.un1_count_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_1_c_inv_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7910\,
            in2 => \N__8726\,
            in3 => \N__10028\,
            lcout => \POWERLED.count_i_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_0\,
            carryout => \POWERLED.un1_count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_2_c_inv_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7904\,
            in2 => \N__7898\,
            in3 => \N__9074\,
            lcout => \POWERLED.count_i_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_1\,
            carryout => \POWERLED.un1_count_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_3_c_inv_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10052\,
            in2 => \N__7889\,
            in3 => \N__9041\,
            lcout => \POWERLED.count_i_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_2\,
            carryout => \POWERLED.un1_count_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_4_c_inv_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7880\,
            in2 => \N__7874\,
            in3 => \N__9008\,
            lcout => \POWERLED.count_i_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_3\,
            carryout => \POWERLED.un1_count_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_5_c_inv_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8618\,
            in2 => \N__8018\,
            in3 => \N__8975\,
            lcout => \POWERLED.count_i_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_4\,
            carryout => \POWERLED.un1_count_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_6_c_inv_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8006\,
            in2 => \N__8000\,
            in3 => \N__8942\,
            lcout => \POWERLED.count_i_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_5\,
            carryout => \POWERLED.un1_count_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_7_c_inv_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11585\,
            in2 => \N__7991\,
            in3 => \N__8908\,
            lcout => \POWERLED.count_i_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_6\,
            carryout => \POWERLED.un1_count_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_8_c_inv_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11645\,
            in2 => \N__7979\,
            in3 => \N__8872\,
            lcout => \POWERLED.count_i_8\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \POWERLED.un1_count_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_9_c_inv_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7970\,
            in2 => \N__7961\,
            in3 => \N__9332\,
            lcout => \POWERLED.count_i_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_8\,
            carryout => \POWERLED.un1_count_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_10_c_inv_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11072\,
            in2 => \N__7952\,
            in3 => \N__9295\,
            lcout => \POWERLED.count_i_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_9\,
            carryout => \POWERLED.un1_count_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_11_c_inv_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9632\,
            in2 => \N__7943\,
            in3 => \N__9263\,
            lcout => \POWERLED.count_i_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_10\,
            carryout => \POWERLED.un1_count_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_12_c_inv_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7922\,
            in2 => \N__7934\,
            in3 => \N__9230\,
            lcout => \POWERLED.count_i_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_11\,
            carryout => \POWERLED.un1_count_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_13_c_inv_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8054\,
            in2 => \N__10766\,
            in3 => \N__9197\,
            lcout => \POWERLED.count_i_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_12\,
            carryout => \POWERLED.un1_count_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_14_c_inv_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9161\,
            in1 => \N__10814\,
            in2 => \N__8048\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_13\,
            carryout => \POWERLED.un1_count_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_15_c_inv_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9424\,
            in1 => \N__10040\,
            in2 => \N__8039\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_15\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_14\,
            carryout => \POWERLED.un1_count_2_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8030\,
            lcout => \POWERLED.un1_count_2_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_1_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8873\,
            in1 => \N__9262\,
            in2 => \_gnd_net_\,
            in3 => \N__9229\,
            lcout => \POWERLED.g0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_RNIS4LI_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16882\,
            lcout => \VCCST_EN_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__9123\,
            in1 => \N__8105\,
            in2 => \_gnd_net_\,
            in3 => \N__8777\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18206\,
            ce => \N__17657\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNID4E61_7_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9320\,
            in1 => \N__8861\,
            in2 => \N__8907\,
            in3 => \N__9287\,
            lcout => OPEN,
            ltout => \POWERLED.un1_countlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI6IPJ2_5_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__8936\,
            in1 => \N__8969\,
            in2 => \N__8021\,
            in3 => \N__8096\,
            lcout => \POWERLED.un1_countlto15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_RNIBHMO_15_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9155\,
            in1 => \N__9420\,
            in2 => \_gnd_net_\,
            in3 => \N__9188\,
            lcout => OPEN,
            ltout => \POWERLED.un1_countlto15_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIOVT24_11_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9257\,
            in1 => \N__9224\,
            in2 => \N__8114\,
            in3 => \N__8111\,
            lcout => \POWERLED.count_RNIOVT24Z0Z_11\,
            ltout => \POWERLED.count_RNIOVT24Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI75RB5_0_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9119\,
            in2 => \N__8099\,
            in3 => \N__17948\,
            lcout => \POWERLED.curr_state_RNI75RB5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICO6R_2_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8996\,
            in1 => \N__9029\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => \POWERLED.un1_countlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8090\,
            lcout => \VDDQ_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_RNO_0_15_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9958\,
            in2 => \_gnd_net_\,
            in3 => \N__17957\,
            lcout => \POWERLED.N_39_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNICTB05_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8288\,
            in2 => \_gnd_net_\,
            in3 => \N__17950\,
            lcout => \PCH_PWRGD.curr_state_RNICTB05Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNICTB05Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNO_0_15_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__17951\,
            in1 => \_gnd_net_\,
            in2 => \N__8069\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_39_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_sys_pwrok_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14239\,
            lcout => \PCH_PWRGD.N_3_i\,
            ltout => \PCH_PWRGD.N_3_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIHB874_0_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__8273\,
            in1 => \N__8236\,
            in2 => \N__8306\,
            in3 => \N__8301\,
            lcout => \PCH_PWRGD.un1_curr_state_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIMQRI1_0_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__8272\,
            in1 => \N__8254\,
            in2 => \N__14247\,
            in3 => \N__8237\,
            lcout => \PCH_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18064\,
            in1 => \N__8201\,
            in2 => \N__8218\,
            in3 => \N__8219\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_0\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18005\,
            in1 => \N__8189\,
            in2 => \_gnd_net_\,
            in3 => \N__8177\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_0\,
            carryout => \PCH_PWRGD.un1_count_1_cry_1\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18065\,
            in1 => \N__8174\,
            in2 => \_gnd_net_\,
            in3 => \N__8162\,
            lcout => \PCH_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_1\,
            carryout => \PCH_PWRGD.un1_count_1_cry_2\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_3_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18006\,
            in1 => \N__8159\,
            in2 => \_gnd_net_\,
            in3 => \N__8147\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_2\,
            carryout => \PCH_PWRGD.un1_count_1_cry_3\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_4_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18066\,
            in1 => \N__8144\,
            in2 => \_gnd_net_\,
            in3 => \N__8132\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_3\,
            carryout => \PCH_PWRGD.un1_count_1_cry_4\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_5_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18007\,
            in1 => \N__8129\,
            in2 => \_gnd_net_\,
            in3 => \N__8117\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_4\,
            carryout => \PCH_PWRGD.un1_count_1_cry_5\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_6_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18067\,
            in1 => \N__8453\,
            in2 => \_gnd_net_\,
            in3 => \N__8441\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_5\,
            carryout => \PCH_PWRGD.un1_count_1_cry_6\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_7_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18008\,
            in1 => \N__8437\,
            in2 => \_gnd_net_\,
            in3 => \N__8423\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_6\,
            carryout => \PCH_PWRGD.un1_count_1_cry_7\,
            clk => \N__18189\,
            ce => 'H',
            sr => \N__8493\
        );

    \PCH_PWRGD.count_8_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18059\,
            in1 => \N__8420\,
            in2 => \_gnd_net_\,
            in3 => \N__8408\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_8\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.count_9_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18000\,
            in1 => \N__8405\,
            in2 => \_gnd_net_\,
            in3 => \N__8393\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_8\,
            carryout => \PCH_PWRGD.un1_count_1_cry_9\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.count_10_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__8389\,
            in2 => \_gnd_net_\,
            in3 => \N__8375\,
            lcout => \PCH_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_9\,
            carryout => \PCH_PWRGD.un1_count_1_cry_10\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.count_11_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17998\,
            in1 => \N__8371\,
            in2 => \_gnd_net_\,
            in3 => \N__8357\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_10\,
            carryout => \PCH_PWRGD.un1_count_1_cry_11\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.count_12_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18057\,
            in1 => \N__8353\,
            in2 => \_gnd_net_\,
            in3 => \N__8339\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_11\,
            carryout => \PCH_PWRGD.un1_count_1_cry_12\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.count_13_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17999\,
            in1 => \N__8336\,
            in2 => \_gnd_net_\,
            in3 => \N__8324\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_12\,
            carryout => \PCH_PWRGD.un1_count_1_cry_13\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.count_14_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18058\,
            in1 => \N__8321\,
            in2 => \_gnd_net_\,
            in3 => \N__8309\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_13\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14\,
            clk => \N__18194\,
            ce => 'H',
            sr => \N__8497\
        );

    \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14918\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_14\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_15_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8522\,
            in2 => \_gnd_net_\,
            in3 => \N__8525\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18196\,
            ce => \N__8510\,
            sr => \N__8498\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16146\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12668\,
            in2 => \N__8470\,
            in3 => \N__8540\,
            lcout => \G_386\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8466\,
            in2 => \N__8603\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8541\,
            in2 => \N__8591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8579\,
            in2 => \N__8546\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8570\,
            in2 => \N__8471\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8561\,
            in3 => \N__8630\,
            lcout => \POWERLED.un1_count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16215\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8612\,
            in2 => \N__8833\,
            in3 => \N__8594\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8829\,
            in2 => \N__8717\,
            in3 => \N__8582\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8705\,
            in2 => \N__8659\,
            in3 => \N__8573\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8655\,
            in2 => \N__8696\,
            in3 => \N__8564\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8545\,
            in1 => \N__8684\,
            in2 => \N__8834\,
            in3 => \N__8552\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8675\,
            in3 => \N__8549\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => \POWERLED.mult1_un159_sum_s_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8729\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16454\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10823\,
            in2 => \N__8746\,
            in3 => \N__8708\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8742\,
            in2 => \N__9905\,
            in3 => \N__8699\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9881\,
            in2 => \N__10088\,
            in3 => \N__8687\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10086\,
            in2 => \N__9863\,
            in3 => \N__8678\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8651\,
            in1 => \N__9809\,
            in2 => \N__8747\,
            in3 => \N__8666\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9773\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => \POWERLED.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8633\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_2_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__8941\,
            in1 => \N__8798\,
            in2 => \N__8807\,
            in3 => \N__8974\,
            lcout => OPEN,
            ltout => \POWERLED.g0_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8816\,
            in1 => \N__9299\,
            in2 => \N__8810\,
            in3 => \N__8909\,
            lcout => \POWERLED.un1_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_4_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9007\,
            in1 => \N__9040\,
            in2 => \_gnd_net_\,
            in3 => \N__9073\,
            lcout => \POWERLED.un1_countlt6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9196\,
            in1 => \N__9160\,
            in2 => \N__9425\,
            in3 => \N__9331\,
            lcout => \POWERLED.g0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_RNIRH3P_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8755\,
            in2 => \_gnd_net_\,
            in3 => \N__10153\,
            lcout => \tmp_RNIRH3P\,
            ltout => \tmp_RNIRH3P_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__9128\,
            in1 => \N__8776\,
            in2 => \N__8765\,
            in3 => \N__8762\,
            lcout => \POWERLED.pwm_out_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8756\,
            in2 => \_gnd_net_\,
            in3 => \N__10154\,
            lcout => \COUNTER.tmp_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10087\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9124\,
            lcout => \PWRBTN_LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18205\,
            ce => \N__9086\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_1_cry_1_c_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10027\,
            in2 => \N__10001\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \POWERLED.un1_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18016\,
            in1 => \N__9069\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_1\,
            carryout => \POWERLED.un1_count_1_cry_2\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_3_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17964\,
            in1 => \N__9036\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_2\,
            carryout => \POWERLED.un1_count_1_cry_3\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_4_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18017\,
            in1 => \N__9003\,
            in2 => \_gnd_net_\,
            in3 => \N__8978\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_3\,
            carryout => \POWERLED.un1_count_1_cry_4\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_5_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17965\,
            in1 => \N__8970\,
            in2 => \_gnd_net_\,
            in3 => \N__8945\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_4\,
            carryout => \POWERLED.un1_count_1_cry_5\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_6_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18018\,
            in1 => \N__8937\,
            in2 => \_gnd_net_\,
            in3 => \N__8912\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_5\,
            carryout => \POWERLED.un1_count_1_cry_6\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_7_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17966\,
            in1 => \N__8900\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_6\,
            carryout => \POWERLED.un1_count_1_cry_7\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_8_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18019\,
            in1 => \N__8865\,
            in2 => \_gnd_net_\,
            in3 => \N__8837\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_7\,
            carryout => \POWERLED.un1_count_1_cry_8\,
            clk => \N__18207\,
            ce => 'H',
            sr => \N__9959\
        );

    \POWERLED.count_9_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17963\,
            in1 => \N__9327\,
            in2 => \_gnd_net_\,
            in3 => \N__9302\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \POWERLED.un1_count_1_cry_9\,
            clk => \N__18208\,
            ce => 'H',
            sr => \N__9967\
        );

    \POWERLED.count_10_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18013\,
            in1 => \N__9288\,
            in2 => \_gnd_net_\,
            in3 => \N__9266\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_9\,
            carryout => \POWERLED.un1_count_1_cry_10\,
            clk => \N__18208\,
            ce => 'H',
            sr => \N__9967\
        );

    \POWERLED.count_11_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17961\,
            in1 => \N__9258\,
            in2 => \_gnd_net_\,
            in3 => \N__9233\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_10\,
            carryout => \POWERLED.un1_count_1_cry_11\,
            clk => \N__18208\,
            ce => 'H',
            sr => \N__9967\
        );

    \POWERLED.count_12_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18014\,
            in1 => \N__9225\,
            in2 => \_gnd_net_\,
            in3 => \N__9200\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_11\,
            carryout => \POWERLED.un1_count_1_cry_12\,
            clk => \N__18208\,
            ce => 'H',
            sr => \N__9967\
        );

    \POWERLED.count_13_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17962\,
            in1 => \N__9192\,
            in2 => \_gnd_net_\,
            in3 => \N__9164\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_12\,
            carryout => \POWERLED.un1_count_1_cry_13\,
            clk => \N__18208\,
            ce => 'H',
            sr => \N__9967\
        );

    \POWERLED.count_14_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18015\,
            in1 => \N__9156\,
            in2 => \_gnd_net_\,
            in3 => \N__9131\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_13\,
            carryout => \POWERLED.un1_count_1_cry_14\,
            clk => \N__18208\,
            ce => 'H',
            sr => \N__9967\
        );

    \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14947\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_14\,
            carryout => \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__14951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryout => \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_15_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9416\,
            in2 => \_gnd_net_\,
            in3 => \N__9428\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18209\,
            ce => \N__9389\,
            sr => \N__9960\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9354\,
            in1 => \N__9378\,
            in2 => \N__9479\,
            in3 => \N__10229\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9379\,
            in1 => \N__9365\,
            in2 => \_gnd_net_\,
            in3 => \N__10138\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9341\,
            in1 => \N__9355\,
            in2 => \_gnd_net_\,
            in3 => \N__10139\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10230\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10141\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9461\,
            in1 => \N__9477\,
            in2 => \_gnd_net_\,
            in3 => \N__10140\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10181\,
            in2 => \N__10235\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9380\,
            in2 => \_gnd_net_\,
            in3 => \N__9359\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9356\,
            in2 => \_gnd_net_\,
            in3 => \N__9335\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9478\,
            in2 => \_gnd_net_\,
            in3 => \N__9455\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10106\,
            in2 => \_gnd_net_\,
            in3 => \N__9452\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10211\,
            in2 => \_gnd_net_\,
            in3 => \N__9449\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10195\,
            in2 => \_gnd_net_\,
            in3 => \N__9446\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__18173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10400\,
            in2 => \_gnd_net_\,
            in3 => \N__9443\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__18173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10427\,
            in2 => \_gnd_net_\,
            in3 => \N__9440\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_4_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10439\,
            in2 => \_gnd_net_\,
            in3 => \N__9437\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10414\,
            in2 => \_gnd_net_\,
            in3 => \N__9434\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10520\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10547\,
            in2 => \_gnd_net_\,
            in3 => \N__9506\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10559\,
            in2 => \_gnd_net_\,
            in3 => \N__9503\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10534\,
            in2 => \_gnd_net_\,
            in3 => \N__9500\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10460\,
            in2 => \_gnd_net_\,
            in3 => \N__9497\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__18176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10487\,
            in2 => \_gnd_net_\,
            in3 => \N__9494\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10499\,
            in2 => \_gnd_net_\,
            in3 => \N__9491\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10474\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10280\,
            in2 => \_gnd_net_\,
            in3 => \N__9485\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10307\,
            in2 => \_gnd_net_\,
            in3 => \N__9482\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10319\,
            in2 => \_gnd_net_\,
            in3 => \N__9536\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10294\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10340\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__18177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10367\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10379\,
            in2 => \_gnd_net_\,
            in3 => \N__9524\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10354\,
            in2 => \_gnd_net_\,
            in3 => \N__9521\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9563\,
            in2 => \_gnd_net_\,
            in3 => \N__9518\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9587\,
            in3 => \N__9515\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9599\,
            in3 => \N__9512\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9574\,
            in2 => \_gnd_net_\,
            in3 => \N__9509\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9595\,
            in1 => \N__9583\,
            in2 => \N__9575\,
            in3 => \N__9562\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13094\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9620\,
            in2 => \N__9649\,
            in3 => \N__9554\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9645\,
            in2 => \N__10736\,
            in3 => \N__9551\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10718\,
            in2 => \N__10805\,
            in3 => \N__9548\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10804\,
            in2 => \N__10706\,
            in3 => \N__9545\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10634\,
            in1 => \N__10862\,
            in2 => \N__9650\,
            in3 => \N__9542\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10850\,
            in3 => \N__9539\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => \POWERLED.mult1_un82_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9653\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10800\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11030\,
            lcout => \POWERLED.un1_count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13067\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12953\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11381\,
            in2 => \N__11401\,
            in3 => \N__9614\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11397\,
            in2 => \N__11342\,
            in3 => \N__9611\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11540\,
            in2 => \N__11437\,
            in3 => \N__9608\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11433\,
            in2 => \N__11522\,
            in3 => \N__9605\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9716\,
            in1 => \N__11498\,
            in2 => \N__11402\,
            in3 => \N__9602\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11462\,
            in2 => \_gnd_net_\,
            in3 => \N__9752\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9715\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12977\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11627\,
            in2 => \N__9673\,
            in3 => \N__9749\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9669\,
            in2 => \N__9746\,
            in3 => \N__9737\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9734\,
            in2 => \N__9724\,
            in3 => \N__9728\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9720\,
            in2 => \N__9692\,
            in3 => \N__9683\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9836\,
            in1 => \N__9680\,
            in2 => \N__9674\,
            in3 => \N__9656\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9920\,
            in3 => \N__9911\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => \POWERLED.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9908\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12997\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10754\,
            in2 => \N__9790\,
            in3 => \N__9893\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9786\,
            in2 => \N__9890\,
            in3 => \N__9872\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9869\,
            in2 => \N__9844\,
            in3 => \N__9851\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9840\,
            in2 => \N__9818\,
            in3 => \N__9800\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10074\,
            in1 => \N__9797\,
            in2 => \N__9791\,
            in3 => \N__9764\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9761\,
            in3 => \N__10091\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => \POWERLED.mult1_un145_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10055\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12025\,
            lcout => \POWERLED.un1_count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__9993\,
            in1 => \_gnd_net_\,
            in2 => \N__18068\,
            in3 => \N__10023\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18203\,
            ce => 'H',
            sr => \N__9968\
        );

    \POWERLED.count_0_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18009\,
            in2 => \_gnd_net_\,
            in3 => \N__9992\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18203\,
            ce => 'H',
            sr => \N__9968\
        );

    \COUNTER.un4_counter_0_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9926\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10166\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10388\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10508\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10448\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10268\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10328\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10256\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER.un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_THRU_LUT4_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10244\,
            lcout => \COUNTER.un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__10241\,
            in1 => \N__10210\,
            in2 => \_gnd_net_\,
            in3 => \N__10136\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10137\,
            in1 => \N__10180\,
            in2 => \_gnd_net_\,
            in3 => \N__10234\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__10209\,
            in1 => \N__10104\,
            in2 => \N__10196\,
            in3 => \N__10179\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__10105\,
            in1 => \N__10160\,
            in2 => \_gnd_net_\,
            in3 => \N__10135\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10558\,
            in1 => \N__10546\,
            in2 => \N__10535\,
            in3 => \N__10519\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10498\,
            in1 => \N__10486\,
            in2 => \N__10475\,
            in3 => \N__10459\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10438\,
            in1 => \N__10426\,
            in2 => \N__10415\,
            in3 => \N__10399\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10378\,
            in1 => \N__10366\,
            in2 => \N__10355\,
            in3 => \N__10339\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10318\,
            in1 => \N__10306\,
            in2 => \N__10295\,
            in3 => \N__10279\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13121\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12047\,
            in2 => \N__10597\,
            in3 => \N__10259\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10593\,
            in2 => \N__10664\,
            in3 => \N__10655\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10652\,
            in2 => \N__10642\,
            in3 => \N__10646\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10638\,
            in2 => \N__10616\,
            in3 => \N__10607\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11021\,
            in1 => \N__10604\,
            in2 => \N__10598\,
            in3 => \N__10580\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10577\,
            in3 => \N__10568\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11020\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18036\,
            in1 => \N__11174\,
            in2 => \N__11675\,
            in3 => \N__11674\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17980\,
            in1 => \N__11104\,
            in2 => \_gnd_net_\,
            in3 => \N__10565\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_2_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18037\,
            in1 => \N__11090\,
            in2 => \_gnd_net_\,
            in3 => \N__10562\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_3_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17981\,
            in1 => \N__11285\,
            in2 => \_gnd_net_\,
            in3 => \N__10691\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_4_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18038\,
            in1 => \N__11312\,
            in2 => \_gnd_net_\,
            in3 => \N__10688\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_5_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17982\,
            in1 => \N__11324\,
            in2 => \_gnd_net_\,
            in3 => \N__10685\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_6_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18039\,
            in1 => \N__11117\,
            in2 => \_gnd_net_\,
            in3 => \N__10682\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_7_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17983\,
            in1 => \N__11299\,
            in2 => \_gnd_net_\,
            in3 => \N__10679\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__18181\,
            ce => 'H',
            sr => \N__10911\
        );

    \VPP_VDDQ.count_8_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18031\,
            in1 => \N__11186\,
            in2 => \_gnd_net_\,
            in3 => \N__10676\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.count_9_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17976\,
            in1 => \N__11147\,
            in2 => \_gnd_net_\,
            in3 => \N__10673\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.count_10_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18028\,
            in1 => \N__11129\,
            in2 => \_gnd_net_\,
            in3 => \N__10670\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.count_11_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17974\,
            in1 => \N__11161\,
            in2 => \_gnd_net_\,
            in3 => \N__10667\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.count_12_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18029\,
            in1 => \N__11228\,
            in2 => \_gnd_net_\,
            in3 => \N__10748\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.count_13_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17975\,
            in1 => \N__11261\,
            in2 => \_gnd_net_\,
            in3 => \N__10745\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.count_14_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18030\,
            in1 => \N__11273\,
            in2 => \_gnd_net_\,
            in3 => \N__10742\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__18185\,
            ce => 'H',
            sr => \N__10916\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14896\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11242\,
            in2 => \_gnd_net_\,
            in3 => \N__10739\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18190\,
            ce => \N__10832\,
            sr => \N__10912\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13063\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11369\,
            in2 => \N__11716\,
            in3 => \N__10721\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11712\,
            in2 => \N__11570\,
            in3 => \N__10709\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11558\,
            in2 => \N__11744\,
            in3 => \N__10694\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11742\,
            in2 => \N__11780\,
            in3 => \N__10853\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10790\,
            in1 => \N__11768\,
            in2 => \N__11717\,
            in3 => \N__10838\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11759\,
            in3 => \N__10835\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10904\,
            in2 => \_gnd_net_\,
            in3 => \N__17958\,
            lcout => \VPP_VDDQ.N_39_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12998\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11743\,
            lcout => \POWERLED.un1_count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10791\,
            lcout => \POWERLED.un1_count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12973\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNII0FM2_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__11906\,
            in1 => \N__11877\,
            in2 => \N__18395\,
            in3 => \N__17946\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.G_110_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIQINR7_0_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__11878\,
            in1 => \N__11907\,
            in2 => \N__10919\,
            in3 => \N__11206\,
            lcout => \VPP_VDDQ.curr_state_RNIQINR7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11881\,
            in2 => \_gnd_net_\,
            in3 => \N__18406\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18201\,
            ce => \N__17651\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100001100"
        )
    port map (
            in0 => \N__11207\,
            in1 => \N__11911\,
            in2 => \N__18410\,
            in3 => \N__11882\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18201\,
            ce => \N__17651\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18060\,
            in1 => \N__12367\,
            in2 => \N__12284\,
            in3 => \N__12280\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_1_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18001\,
            in1 => \N__12380\,
            in2 => \_gnd_net_\,
            in3 => \N__10877\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_2_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18061\,
            in1 => \N__12392\,
            in2 => \_gnd_net_\,
            in3 => \N__10874\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_3_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18002\,
            in1 => \N__11945\,
            in2 => \_gnd_net_\,
            in3 => \N__10871\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_4_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18062\,
            in1 => \N__12410\,
            in2 => \_gnd_net_\,
            in3 => \N__10868\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_5_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18003\,
            in1 => \N__12437\,
            in2 => \_gnd_net_\,
            in3 => \N__10865\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_6_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18063\,
            in1 => \N__12449\,
            in2 => \_gnd_net_\,
            in3 => \N__10946\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_7_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18004\,
            in1 => \N__11972\,
            in2 => \_gnd_net_\,
            in3 => \N__10943\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__18166\,
            ce => 'H',
            sr => \N__12192\
        );

    \RSMRST_PWRGD.count_8_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18051\,
            in1 => \N__11984\,
            in2 => \_gnd_net_\,
            in3 => \N__10940\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.count_9_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17993\,
            in1 => \N__11959\,
            in2 => \_gnd_net_\,
            in3 => \N__10937\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.count_10_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18048\,
            in1 => \N__12424\,
            in2 => \_gnd_net_\,
            in3 => \N__10934\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.count_11_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17991\,
            in1 => \N__12227\,
            in2 => \_gnd_net_\,
            in3 => \N__10931\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.count_12_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18049\,
            in1 => \N__12353\,
            in2 => \_gnd_net_\,
            in3 => \N__10928\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.count_13_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17992\,
            in1 => \N__12254\,
            in2 => \_gnd_net_\,
            in3 => \N__10925\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.count_14_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18050\,
            in1 => \N__12266\,
            in2 => \_gnd_net_\,
            in3 => \N__10922\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__18171\,
            ce => 'H',
            sr => \N__12199\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14886\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12241\,
            in2 => \_gnd_net_\,
            in3 => \N__11057\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18174\,
            ce => \N__12164\,
            sr => \N__12206\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12853\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12038\,
            in2 => \N__10978\,
            in3 => \N__11054\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10974\,
            in2 => \N__11051\,
            in3 => \N__11042\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11039\,
            in2 => \N__11029\,
            in3 => \N__11033\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11025\,
            in2 => \N__10997\,
            in3 => \N__10988\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12533\,
            in1 => \N__10985\,
            in2 => \N__10979\,
            in3 => \N__10961\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10958\,
            in3 => \N__10949\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => \POWERLED.mult1_un96_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11327\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11323\,
            in1 => \N__11311\,
            in2 => \N__11300\,
            in3 => \N__11284\,
            lcout => \VPP_VDDQ.un6_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11272\,
            in1 => \N__11260\,
            in2 => \N__11249\,
            in3 => \N__11227\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11078\,
            in1 => \N__11135\,
            in2 => \N__11216\,
            in3 => \N__11213\,
            lcout => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11185\,
            in1 => \N__11173\,
            in2 => \N__11162\,
            in3 => \N__11146\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11128\,
            in1 => \N__11116\,
            in2 => \N__11105\,
            in3 => \N__11089\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12538\,
            lcout => \POWERLED.un1_count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12911\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12653\,
            in2 => \N__12677\,
            in3 => \N__11360\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12631\,
            in2 => \N__12458\,
            in3 => \N__11357\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12605\,
            in2 => \N__12719\,
            in3 => \N__11354\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12715\,
            in2 => \N__12584\,
            in3 => \N__11351\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11609\,
            in1 => \N__12644\,
            in2 => \N__12791\,
            in3 => \N__11348\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12746\,
            in3 => \N__11345\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11608\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11576\,
            in2 => \N__11479\,
            in3 => \N__11330\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11475\,
            in2 => \N__11549\,
            in3 => \N__11531\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11528\,
            in2 => \N__11617\,
            in3 => \N__11510\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11613\,
            in2 => \N__11507\,
            in3 => \N__11489\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11421\,
            in1 => \N__11486\,
            in2 => \N__11480\,
            in3 => \N__11453\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11450\,
            in3 => \N__11441\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11420\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12928\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13043\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12716\,
            lcout => \POWERLED.un1_count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9L40B_0_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11654\,
            in2 => \_gnd_net_\,
            in3 => \N__17952\,
            lcout => \POWERLED.func_state_RNI9L40BZ0Z_0\,
            ltout => \POWERLED.func_state_RNI9L40BZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_esr_RNO_0_15_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__17953\,
            in1 => \_gnd_net_\,
            in2 => \N__11630\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12949\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11618\,
            lcout => \POWERLED.un1_count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12907\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13039\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11681\,
            in2 => \N__11698\,
            in3 => \N__11561\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11694\,
            in2 => \N__11846\,
            in3 => \N__11552\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11831\,
            in2 => \N__12026\,
            in3 => \N__11771\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12024\,
            in2 => \N__11819\,
            in3 => \N__11762\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11738\,
            in1 => \N__11804\,
            in2 => \N__11699\,
            in3 => \N__11750\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11792\,
            in2 => \_gnd_net_\,
            in3 => \N__11747\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => \POWERLED.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11720\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12012\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNINEBT1_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__11876\,
            in1 => \N__11905\,
            in2 => \_gnd_net_\,
            in3 => \N__18382\,
            lcout => \VPP_VDDQ.N_32_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIE317A_0_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__15079\,
            in1 => \N__16753\,
            in2 => \_gnd_net_\,
            in3 => \N__16693\,
            lcout => \POWERLED.count_off_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111010011001"
        )
    port map (
            in0 => \N__11879\,
            in1 => \N__13152\,
            in2 => \N__11912\,
            in3 => \N__17960\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001111000010"
        )
    port map (
            in0 => \N__13153\,
            in1 => \N__11880\,
            in2 => \N__11849\,
            in3 => \N__18405\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13025\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13205\,
            in2 => \N__13279\,
            in3 => \N__11834\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13275\,
            in2 => \N__13223\,
            in3 => \N__11822\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13411\,
            in2 => \N__13469\,
            in3 => \N__11807\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13448\,
            in2 => \N__13415\,
            in3 => \N__11795\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12008\,
            in1 => \N__13430\,
            in2 => \N__13280\,
            in3 => \N__11783\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13370\,
            in2 => \_gnd_net_\,
            in3 => \N__12029\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__13395\,
            in1 => \N__13396\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16574\,
            in1 => \N__12333\,
            in2 => \_gnd_net_\,
            in3 => \N__12310\,
            lcout => \RSMRSTn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18165\,
            ce => \N__17662\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100010000"
        )
    port map (
            in0 => \N__12334\,
            in1 => \N__11930\,
            in2 => \N__12313\,
            in3 => \N__16575\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18165\,
            ce => \N__17662\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__12335\,
            in1 => \_gnd_net_\,
            in2 => \N__12314\,
            in3 => \N__11921\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18165\,
            ce => \N__17662\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIF1MK1_3_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11983\,
            in1 => \N__11971\,
            in2 => \N__11960\,
            in3 => \N__11944\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un4_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIR8OP4_10_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12215\,
            in1 => \N__12398\,
            in2 => \N__11933\,
            in3 => \N__12341\,
            lcout => \RSMRST_PWRGD.N_1_i\,
            ltout => \RSMRST_PWRGD.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_0_o2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__12312\,
            in1 => \_gnd_net_\,
            in2 => \N__11924\,
            in3 => \N__16570\,
            lcout => \RSMRST_PWRGD.N_85\,
            ltout => \RSMRST_PWRGD.N_85_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNI6HIT6_0_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__12332\,
            in1 => \_gnd_net_\,
            in2 => \N__11915\,
            in3 => \N__17949\,
            lcout => \RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIKOU91_10_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12448\,
            in1 => \N__12436\,
            in2 => \N__12425\,
            in3 => \N__12409\,
            lcout => \RSMRST_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIAEU91_12_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__12391\,
            in1 => \N__12379\,
            in2 => \N__12368\,
            in3 => \N__12352\,
            lcout => \RSMRST_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIGMMA1_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011100"
        )
    port map (
            in0 => \N__12331\,
            in1 => \N__12311\,
            in2 => \N__16579\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_51_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNIE05H_15_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12265\,
            in1 => \N__12253\,
            in2 => \N__12242\,
            in3 => \N__12226\,
            lcout => \RSMRST_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12191\,
            in2 => \_gnd_net_\,
            in3 => \N__17959\,
            lcout => \RSMRST_PWRGD.N_39_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12155\,
            in1 => \N__12113\,
            in2 => \N__12098\,
            in3 => \N__12073\,
            lcout => rsmrst_pwrgd_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13090\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13117\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12871\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12464\,
            in2 => \N__12496\,
            in3 => \N__12563\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12492\,
            in2 => \N__12560\,
            in3 => \N__12551\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12548\,
            in2 => \N__12539\,
            in3 => \N__12542\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12537\,
            in2 => \N__12515\,
            in3 => \N__12506\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12813\,
            in1 => \N__12503\,
            in2 => \N__12497\,
            in3 => \N__12479\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12476\,
            in3 => \N__12467\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12854\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_4_l_fx_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12632\,
            in2 => \N__12717\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12890\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12872\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12812\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_7_l_fx_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__12790\,
            in1 => \_gnd_net_\,
            in2 => \N__12718\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12889\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12638\,
            in2 => \N__12763\,
            in3 => \N__12620\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12759\,
            in2 => \N__12617\,
            in3 => \N__12599\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12822\,
            in2 => \N__12596\,
            in3 => \N__12575\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12572\,
            in2 => \N__12829\,
            in3 => \N__12776\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12711\,
            in1 => \N__12773\,
            in2 => \N__12764\,
            in3 => \N__12737\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12734\,
            in3 => \N__12722\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => \POWERLED.mult1_un110_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12680\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__17399\,
            in1 => \N__15080\,
            in2 => \N__14807\,
            in3 => \N__16702\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18184\,
            ce => \N__17652\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFHLJ_0_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16121\,
            in2 => \N__16213\,
            in3 => \N__15560\,
            lcout => \POWERLED.un1_dutycycle_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__17400\,
            in1 => \N__15081\,
            in2 => \N__14789\,
            in3 => \N__16703\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18184\,
            ce => \N__17652\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFHLJ_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16122\,
            in2 => \N__16214\,
            in3 => \N__15561\,
            lcout => \POWERLED.dutycycle_RNIFHLJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16195\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__16701\,
            in1 => \N__14009\,
            in2 => \N__15088\,
            in3 => \N__16754\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18184\,
            ce => \N__17652\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVL3D_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16123\,
            in2 => \N__15626\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \POWERLED.un1_dutycycle_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12983\,
            in2 => \_gnd_net_\,
            in3 => \N__12956\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_0\,
            carryout => \POWERLED.un1_dutycycle_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15434\,
            in2 => \N__15451\,
            in3 => \N__12935\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_1\,
            carryout => \POWERLED.un1_dutycycle_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15782\,
            in2 => \N__15809\,
            in3 => \N__12914\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_2\,
            carryout => \POWERLED.un1_dutycycle_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13709\,
            in2 => \N__13721\,
            in3 => \N__12893\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_3\,
            carryout => \POWERLED.un1_dutycycle_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13703\,
            in2 => \N__15503\,
            in3 => \N__12875\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_4\,
            carryout => \POWERLED.un1_dutycycle_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15821\,
            in2 => \N__15845\,
            in3 => \N__12857\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_5\,
            carryout => \POWERLED.un1_dutycycle_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13835\,
            in2 => \N__13850\,
            in3 => \N__12836\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_6\,
            carryout => \POWERLED.un1_dutycycle_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13901\,
            in2 => \N__13919\,
            in3 => \N__13097\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \POWERLED.un1_dutycycle_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13865\,
            in2 => \N__15101\,
            in3 => \N__13070\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_8\,
            carryout => \POWERLED.un1_dutycycle_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14015\,
            in2 => \N__13973\,
            in3 => \N__13046\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_9\,
            carryout => \POWERLED.un1_dutycycle_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13871\,
            in2 => \N__13883\,
            in3 => \N__13028\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_10\,
            carryout => \POWERLED.un1_dutycycle_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13982\,
            in2 => \N__13999\,
            in3 => \N__13010\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_11\,
            carryout => \POWERLED.un1_dutycycle_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13952\,
            in2 => \N__13946\,
            in3 => \N__13007\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_12\,
            carryout => \POWERLED.un1_dutycycle_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13958\,
            in2 => \N__13859\,
            in3 => \N__13004\,
            lcout => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_13\,
            carryout => \POWERLED.un1_dutycycle_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13964\,
            in2 => \N__13892\,
            in3 => \N__13001\,
            lcout => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_14\,
            carryout => \POWERLED.un1_dutycycle_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15221\,
            in2 => \N__14270\,
            in3 => \N__13211\,
            lcout => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13208\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100101"
        )
    port map (
            in0 => \N__13182\,
            in1 => \_gnd_net_\,
            in2 => \N__13199\,
            in3 => \N__13165\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13246\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13186\,
            in3 => \N__13164\,
            lcout => \POWERLED.mult1_un47_sum_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13178\,
            lcout => \POWERLED.un1_dutycycle_1_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__13198\,
            in1 => \_gnd_net_\,
            in2 => \N__13187\,
            in3 => \N__13166\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIO3TP_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__18355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13154\,
            lcout => \VPP_VDDQ_un2_vpp_en_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13262\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13130\,
            in3 => \N__13325\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13322\,
            in3 => \N__13313\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14931\,
            in2 => \N__13310\,
            in3 => \N__13301\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13298\,
            in2 => \N__14945\,
            in3 => \N__13289\,
            lcout => \POWERLED.mult1_un47_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_5\,
            carryout => \POWERLED.mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13358\,
            in3 => \N__13286\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => \POWERLED.mult1_un54_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13283\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13261\,
            lcout => \POWERLED.un1_dutycycle_1_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13247\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13232\,
            in3 => \N__13214\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13348\,
            in2 => \N__13334\,
            in3 => \N__13460\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14938\,
            in2 => \N__13457\,
            in3 => \N__13442\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14939\,
            in2 => \N__13439\,
            in3 => \N__13418\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13410\,
            in1 => \N__13397\,
            in2 => \N__13379\,
            in3 => \N__13364\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13361\,
            lcout => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__13347\,
            in1 => \N__13349\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_0_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__16519\,
            in1 => \N__14132\,
            in2 => \_gnd_net_\,
            in3 => \N__14105\,
            lcout => \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18052\,
            in1 => \N__14054\,
            in2 => \N__14081\,
            in3 => \N__14080\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_0\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17994\,
            in1 => \N__14041\,
            in2 => \_gnd_net_\,
            in3 => \N__13496\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_0\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_1\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_2_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18053\,
            in1 => \N__14150\,
            in2 => \_gnd_net_\,
            in3 => \N__13493\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_1\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_2\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17995\,
            in1 => \N__14177\,
            in2 => \_gnd_net_\,
            in3 => \N__13490\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_2\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_3\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_4_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18054\,
            in1 => \N__14375\,
            in2 => \_gnd_net_\,
            in3 => \N__13487\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_3\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_4\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_5_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17996\,
            in1 => \N__14189\,
            in2 => \_gnd_net_\,
            in3 => \N__13484\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_4\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_5\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_6_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18055\,
            in1 => \N__14402\,
            in2 => \_gnd_net_\,
            in3 => \N__13481\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_5\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_6\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_7_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17997\,
            in1 => \N__14414\,
            in2 => \_gnd_net_\,
            in3 => \N__13478\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_6\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_7\,
            clk => \N__18167\,
            ce => 'H',
            sr => \N__14604\
        );

    \ALL_SYS_PWRGD.count_8_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18047\,
            in1 => \N__14389\,
            in2 => \_gnd_net_\,
            in3 => \N__13475\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_8\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.count_9_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17990\,
            in1 => \N__14066\,
            in2 => \_gnd_net_\,
            in3 => \N__13472\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_8\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_9\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.count_10_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18044\,
            in1 => \N__14027\,
            in2 => \_gnd_net_\,
            in3 => \N__13514\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_9\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_10\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.count_11_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17988\,
            in1 => \N__14164\,
            in2 => \_gnd_net_\,
            in3 => \N__13511\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_10\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_11\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.count_12_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18045\,
            in1 => \N__14318\,
            in2 => \_gnd_net_\,
            in3 => \N__13508\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_11\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_12\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.count_13_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17989\,
            in1 => \N__14345\,
            in2 => \_gnd_net_\,
            in3 => \N__13505\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_12\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_13\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.count_14_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18046\,
            in1 => \N__14357\,
            in2 => \_gnd_net_\,
            in3 => \N__13502\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_13\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_14\,
            clk => \N__18172\,
            ce => 'H',
            sr => \N__14615\
        );

    \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14855\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_14\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_15_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14332\,
            in2 => \_gnd_net_\,
            in3 => \N__13499\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18175\,
            ce => \N__14573\,
            sr => \N__14614\
        );

    \POWERLED.count_off_esr_RNI7VF31_15_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13811\,
            in1 => \N__13829\,
            in2 => \N__13790\,
            in3 => \N__13598\,
            lcout => \POWERLED.func_state_ns_0_i_o2_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI092U_10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13637\,
            in1 => \N__13655\,
            in2 => \N__13619\,
            in3 => \N__13673\,
            lcout => \POWERLED.func_state_ns_0_i_o2_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINOP11_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__14498\,
            in1 => \N__14514\,
            in2 => \_gnd_net_\,
            in3 => \N__14536\,
            lcout => \POWERLED.un1_func_state11_2_i_o6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIR2P11_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13528\,
            in1 => \N__13543\,
            in2 => \N__13691\,
            in3 => \N__13561\,
            lcout => \POWERLED.func_state_ns_0_i_o2_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIFHLP9_8_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16341\,
            in1 => \N__17019\,
            in2 => \N__15089\,
            in3 => \N__15418\,
            lcout => \POWERLED.N_68_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIU9HM_4_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14460\,
            in2 => \_gnd_net_\,
            in3 => \N__14497\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_sqmuxa_i_o6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIO5BO1_2_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__14757\,
            in1 => \N__14515\,
            in2 => \N__13580\,
            in3 => \N__14537\,
            lcout => \POWERLED.N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18024\,
            in1 => \N__15484\,
            in2 => \N__13577\,
            in3 => \N__13576\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \POWERLED.un1_count_off_1_cry_0\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17970\,
            in1 => \N__13562\,
            in2 => \_gnd_net_\,
            in3 => \N__13550\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_0\,
            carryout => \POWERLED.un1_count_off_1_cry_1\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18025\,
            in1 => \N__15013\,
            in2 => \_gnd_net_\,
            in3 => \N__13547\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_1\,
            carryout => \POWERLED.un1_count_off_1_cry_2\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_3_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17971\,
            in1 => \N__13544\,
            in2 => \_gnd_net_\,
            in3 => \N__13532\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_2\,
            carryout => \POWERLED.un1_count_off_1_cry_3\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18026\,
            in1 => \N__13529\,
            in2 => \_gnd_net_\,
            in3 => \N__13517\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_3\,
            carryout => \POWERLED.un1_count_off_1_cry_4\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17972\,
            in1 => \N__15031\,
            in2 => \_gnd_net_\,
            in3 => \N__13697\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_4\,
            carryout => \POWERLED.un1_count_off_1_cry_5\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_6_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18027\,
            in1 => \N__14992\,
            in2 => \_gnd_net_\,
            in3 => \N__13694\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_5\,
            carryout => \POWERLED.un1_count_off_1_cry_6\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_7_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17973\,
            in1 => \N__13690\,
            in2 => \_gnd_net_\,
            in3 => \N__13676\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_6\,
            carryout => \POWERLED.un1_count_off_1_cry_7\,
            clk => \N__18178\,
            ce => 'H',
            sr => \N__13759\
        );

    \POWERLED.count_off_8_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18023\,
            in1 => \N__13672\,
            in2 => \_gnd_net_\,
            in3 => \N__13658\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \POWERLED.un1_count_off_1_cry_8\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.count_off_9_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17969\,
            in1 => \N__13654\,
            in2 => \_gnd_net_\,
            in3 => \N__13640\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_8\,
            carryout => \POWERLED.un1_count_off_1_cry_9\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.count_off_10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18020\,
            in1 => \N__13636\,
            in2 => \_gnd_net_\,
            in3 => \N__13622\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_9\,
            carryout => \POWERLED.un1_count_off_1_cry_10\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.count_off_11_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17967\,
            in1 => \N__13615\,
            in2 => \_gnd_net_\,
            in3 => \N__13601\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_10\,
            carryout => \POWERLED.un1_count_off_1_cry_11\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.count_off_12_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18021\,
            in1 => \N__13597\,
            in2 => \_gnd_net_\,
            in3 => \N__13583\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_11\,
            carryout => \POWERLED.un1_count_off_1_cry_12\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.count_off_13_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17968\,
            in1 => \N__13828\,
            in2 => \_gnd_net_\,
            in3 => \N__13814\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_12\,
            carryout => \POWERLED.un1_count_off_1_cry_13\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.count_off_14_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18022\,
            in1 => \N__13810\,
            in2 => \_gnd_net_\,
            in3 => \N__13796\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_13\,
            carryout => \POWERLED.un1_count_off_1_cry_14\,
            clk => \N__18182\,
            ce => 'H',
            sr => \N__13760\
        );

    \POWERLED.un1_count_off_1_cry_14_c_THRU_CRY_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14895\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_14\,
            carryout => \POWERLED.un1_count_off_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_esr_15_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13786\,
            in2 => \_gnd_net_\,
            in3 => \N__13793\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18186\,
            ce => \N__13772\,
            sr => \N__13755\
        );

    \POWERLED.dutycycle_fast_RNI2GSK_6_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15602\,
            in2 => \N__13936\,
            in3 => \N__16453\,
            lcout => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\,
            ltout => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQAI81_4_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15601\,
            in1 => \N__15667\,
            in2 => \N__13712\,
            in3 => \N__15539\,
            lcout => \POWERLED.dutycycle_RNIQAI81Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOQLJ_4_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__15540\,
            in1 => \_gnd_net_\,
            in2 => \N__15687\,
            in3 => \N__15603\,
            lcout => \POWERLED.dutycycle_RNIOQLJZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_6_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__17405\,
            in1 => \N__16834\,
            in2 => \N__17107\,
            in3 => \N__15907\,
            lcout => \POWERLED.dutycycle_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18191\,
            ce => \N__17653\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIBPSK_6_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15886\,
            in2 => \N__13937\,
            in3 => \N__16089\,
            lcout => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNILMLM_6_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15666\,
            in2 => \N__15769\,
            in3 => \N__13929\,
            lcout => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\,
            ltout => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJL1R1_6_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13904\,
            in3 => \N__15707\,
            lcout => \POWERLED.dutycycle_RNIJL1R1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIC8C11_15_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__15266\,
            in1 => \N__15336\,
            in2 => \N__15218\,
            in3 => \N__15276\,
            lcout => \POWERLED.dutycycle_RNIC8C11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO18N_9_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15325\,
            in2 => \N__15766\,
            in3 => \N__15888\,
            lcout => \POWERLED.dutycycle_RNIO18NZ0Z_9\,
            ltout => \POWERLED.dutycycle_RNIO18NZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQ09G1_10_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15261\,
            in1 => \N__15748\,
            in2 => \N__13874\,
            in3 => \N__17236\,
            lcout => \POWERLED.dutycycle_RNIQ09G1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIB1FL_8_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15674\,
            in2 => \N__17257\,
            in3 => \N__17181\,
            lcout => \POWERLED.dutycycle_RNIB1FLZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI84C11_14_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__15326\,
            in1 => \N__15143\,
            in2 => \N__15278\,
            in3 => \N__15335\,
            lcout => \POWERLED.dutycycle_RNI84C11Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2V0P_10_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__15752\,
            in1 => \_gnd_net_\,
            in2 => \N__17258\,
            in3 => \N__15262\,
            lcout => \POWERLED.dutycycle_RNI2V0PZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJNBA1_6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__13849\,
            in1 => \N__15747\,
            in2 => \N__15688\,
            in3 => \N__16033\,
            lcout => \POWERLED.dutycycle_RNIJNBA1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE4FL_9_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15887\,
            in2 => \N__15158\,
            in3 => \N__17182\,
            lcout => \POWERLED.dutycycle_RNIE4FLZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_0_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18573\,
            in1 => \N__16874\,
            in2 => \_gnd_net_\,
            in3 => \N__16629\,
            lcout => \POWERLED.N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI712I1_15_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__14000\,
            in1 => \N__15197\,
            in2 => \N__15159\,
            in3 => \N__17261\,
            lcout => \POWERLED.dutycycle_RNI712I1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1VLG_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15330\,
            in2 => \_gnd_net_\,
            in3 => \N__15770\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIF3561_9_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__15157\,
            in1 => \N__17193\,
            in2 => \N__13976\,
            in3 => \N__15895\,
            lcout => \POWERLED.dutycycle_RNIF3561Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI53MG_14_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15279\,
            in2 => \_gnd_net_\,
            in3 => \N__15333\,
            lcout => \POWERLED.dutycycle_RNI53MGZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31MG_12_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15332\,
            in1 => \_gnd_net_\,
            in2 => \N__15161\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI31MGZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI73C11_15_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__15198\,
            in1 => \N__15334\,
            in2 => \N__17269\,
            in3 => \N__15153\,
            lcout => \POWERLED.dutycycle_RNI73C11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31MG_0_12_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__15331\,
            in1 => \_gnd_net_\,
            in2 => \N__15160\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI31MG_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI75MG_15_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15284\,
            in3 => \N__15214\,
            lcout => \POWERLED.dutycycle_RNI75MGZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_0_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__14108\,
            in1 => \N__14428\,
            in2 => \N__14138\,
            in3 => \N__14261\,
            lcout => \ALL_SYS_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18168\,
            ce => \N__17663\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__16517\,
            in1 => \N__14133\,
            in2 => \_gnd_net_\,
            in3 => \N__14106\,
            lcout => \VCCIN_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18168\,
            ce => \N__17663\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_1_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100100010"
        )
    port map (
            in0 => \N__16518\,
            in1 => \N__14107\,
            in2 => \N__14432\,
            in3 => \N__14134\,
            lcout => \ALL_SYS_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18168\,
            ce => \N__17663\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNI10LN5_0_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__14103\,
            in1 => \N__14131\,
            in2 => \N__16520\,
            in3 => \N__14427\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNISHOG6_0_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14192\,
            in3 => \N__17947\,
            lcout => \ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14188\,
            in1 => \N__14176\,
            in2 => \N__14165\,
            in3 => \N__14149\,
            lcout => \ALL_SYS_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNI6P052_0_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__14130\,
            in1 => \N__14104\,
            in2 => \_gnd_net_\,
            in3 => \N__16516\,
            lcout => \ALL_SYS_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__14065\,
            in1 => \N__14053\,
            in2 => \N__14042\,
            in3 => \N__14026\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14306\,
            in1 => \N__14441\,
            in2 => \N__14435\,
            in3 => \N__14363\,
            lcout => \ALL_SYS_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14413\,
            in1 => \N__14401\,
            in2 => \N__14390\,
            in3 => \N__14374\,
            lcout => \ALL_SYS_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14356\,
            in1 => \N__14344\,
            in2 => \N__14333\,
            in3 => \N__14317\,
            lcout => \ALL_SYS_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_RNI34841_15_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__14563\,
            in1 => \N__14681\,
            in2 => \N__14825\,
            in3 => \N__14735\,
            lcout => \POWERLED.dutycycle_1_sqmuxa_i_o6_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIRB454_10_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14297\,
            in1 => \N__14291\,
            in2 => \N__15470\,
            in3 => \N__14285\,
            lcout => \POWERLED.N_100\,
            ltout => \POWERLED.N_100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJHFT5_6_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__14758\,
            in1 => \N__14279\,
            in2 => \N__14273\,
            in3 => \N__14461\,
            lcout => \POWERLED.N_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIK90F_10_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14663\,
            in1 => \N__14699\,
            in2 => \N__14645\,
            in3 => \N__14717\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_sqmuxa_i_o6_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIHJP92_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14476\,
            in1 => \N__14551\,
            in2 => \N__14624\,
            in3 => \N__14621\,
            lcout => \POWERLED.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14594\,
            in2 => \_gnd_net_\,
            in3 => \N__17956\,
            lcout => \ALL_SYS_PWRGD.N_39_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18040\,
            in1 => \N__14564\,
            in2 => \N__16670\,
            in3 => \N__16669\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \POWERLED.un1_count_clk_1_cry_0\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17984\,
            in1 => \N__14552\,
            in2 => \_gnd_net_\,
            in3 => \N__14540\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_0\,
            carryout => \POWERLED.un1_count_clk_1_cry_1\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18041\,
            in1 => \N__14535\,
            in2 => \_gnd_net_\,
            in3 => \N__14519\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_1\,
            carryout => \POWERLED.un1_count_clk_1_cry_2\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17985\,
            in1 => \N__14516\,
            in2 => \_gnd_net_\,
            in3 => \N__14501\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_2\,
            carryout => \POWERLED.un1_count_clk_1_cry_3\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_4_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18042\,
            in1 => \N__14496\,
            in2 => \_gnd_net_\,
            in3 => \N__14480\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_3\,
            carryout => \POWERLED.un1_count_clk_1_cry_4\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_5_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17986\,
            in1 => \N__14477\,
            in2 => \_gnd_net_\,
            in3 => \N__14465\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_4\,
            carryout => \POWERLED.un1_count_clk_1_cry_5\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18043\,
            in1 => \N__14462\,
            in2 => \_gnd_net_\,
            in3 => \N__14444\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_5\,
            carryout => \POWERLED.un1_count_clk_1_cry_6\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_7_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17987\,
            in1 => \N__14759\,
            in2 => \_gnd_net_\,
            in3 => \N__14741\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_6\,
            carryout => \POWERLED.un1_count_clk_1_cry_7\,
            clk => \N__18179\,
            ce => 'H',
            sr => \N__15398\
        );

    \POWERLED.count_clk_8_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18035\,
            in1 => \N__17009\,
            in2 => \_gnd_net_\,
            in3 => \N__14738\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \POWERLED.un1_count_clk_1_cry_8\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.count_clk_9_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17979\,
            in1 => \N__14734\,
            in2 => \_gnd_net_\,
            in3 => \N__14720\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_8\,
            carryout => \POWERLED.un1_count_clk_1_cry_9\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.count_clk_10_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18032\,
            in1 => \N__14716\,
            in2 => \_gnd_net_\,
            in3 => \N__14702\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_9\,
            carryout => \POWERLED.un1_count_clk_1_cry_10\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.count_clk_11_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17977\,
            in1 => \N__14698\,
            in2 => \_gnd_net_\,
            in3 => \N__14684\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_10\,
            carryout => \POWERLED.un1_count_clk_1_cry_11\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.count_clk_12_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18033\,
            in1 => \N__14680\,
            in2 => \_gnd_net_\,
            in3 => \N__14666\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_11\,
            carryout => \POWERLED.un1_count_clk_1_cry_12\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.count_clk_13_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17978\,
            in1 => \N__14662\,
            in2 => \_gnd_net_\,
            in3 => \N__14648\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_12\,
            carryout => \POWERLED.un1_count_clk_1_cry_13\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.count_clk_14_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18034\,
            in1 => \N__14641\,
            in2 => \_gnd_net_\,
            in3 => \N__14627\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_13\,
            carryout => \POWERLED.un1_count_clk_1_cry_14\,
            clk => \N__18183\,
            ce => 'H',
            sr => \N__15397\
        );

    \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14876\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_14\,
            carryout => \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_15_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14821\,
            in2 => \_gnd_net_\,
            in3 => \N__14828\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18187\,
            ce => \N__15359\,
            sr => \N__15396\
        );

    \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16375\,
            in2 => \N__16379\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \POWERLED.dutycycle_cry_c_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16284\,
            in2 => \N__16151\,
            in3 => \N__14792\,
            lcout => \POWERLED.dutycycle_s_0\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_c_0_THRU_CO\,
            carryout => \POWERLED.dutycycle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16225\,
            in2 => \N__16313\,
            in3 => \N__14774\,
            lcout => \POWERLED.dutycycle_s_1\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_0\,
            carryout => \POWERLED.dutycycle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_1_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16288\,
            in2 => \N__16456\,
            in3 => \N__14771\,
            lcout => \POWERLED.dutycycle_s_2\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_1\,
            carryout => \POWERLED.dutycycle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17410\,
            in1 => \N__15607\,
            in2 => \N__16314\,
            in3 => \N__14768\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_2\,
            carryout => \POWERLED.dutycycle_cry_3\,
            clk => \N__18192\,
            ce => \N__17658\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17411\,
            in1 => \N__16292\,
            in2 => \N__15559\,
            in3 => \N__14765\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_3\,
            carryout => \POWERLED.dutycycle_cry_4\,
            clk => \N__18192\,
            ce => \N__17658\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_RNI937G9_4_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16091\,
            in2 => \N__16315\,
            in3 => \N__14762\,
            lcout => \POWERLED.dutycycle_s_5\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_4\,
            carryout => \POWERLED.dutycycle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_RNIB57G9_5_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16296\,
            in2 => \N__16037\,
            in3 => \N__14978\,
            lcout => \POWERLED.dutycycle_s_6\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_5\,
            carryout => \POWERLED.dutycycle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17403\,
            in1 => \N__16297\,
            in2 => \N__15691\,
            in3 => \N__14975\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \POWERLED.dutycycle_cry_7\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17409\,
            in1 => \N__17183\,
            in2 => \N__16316\,
            in3 => \N__14972\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_7\,
            carryout => \POWERLED.dutycycle_cry_8\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_9_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17404\,
            in1 => \N__16301\,
            in2 => \N__15896\,
            in3 => \N__14969\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_8\,
            carryout => \POWERLED.dutycycle_cry_9\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17406\,
            in1 => \N__15756\,
            in2 => \N__16317\,
            in3 => \N__14966\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_9\,
            carryout => \POWERLED.dutycycle_cry_10\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17401\,
            in1 => \N__16305\,
            in2 => \N__17259\,
            in3 => \N__14963\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_10\,
            carryout => \POWERLED.dutycycle_cry_11\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17407\,
            in1 => \N__15144\,
            in2 => \N__16318\,
            in3 => \N__14960\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_11\,
            carryout => \POWERLED.dutycycle_cry_12\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17402\,
            in1 => \N__16309\,
            in2 => \N__15338\,
            in3 => \N__14957\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_12\,
            carryout => \POWERLED.dutycycle_cry_13\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__17408\,
            in1 => \N__15277\,
            in2 => \N__16319\,
            in3 => \N__14954\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_13\,
            carryout => \POWERLED.dutycycle_cry_14\,
            clk => \N__18195\,
            ce => \N__17656\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000100010010"
        )
    port map (
            in0 => \N__16283\,
            in1 => \N__17398\,
            in2 => \N__15220\,
            in3 => \N__15341\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18197\,
            ce => \N__17654\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNINVIV_4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15337\,
            in1 => \N__15558\,
            in2 => \N__17270\,
            in3 => \N__15283\,
            lcout => \POWERLED.func_state_ns_0_i_o3_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1MPT_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__15146\,
            in1 => \N__16457\,
            in2 => \N__15625\,
            in3 => \N__15767\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_ns_0_i_o3_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIUTDP2_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15167\,
            in2 => \N__15230\,
            in3 => \N__15227\,
            lcout => \POWERLED.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI681S_15_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15894\,
            in1 => \N__15689\,
            in2 => \N__15219\,
            in3 => \N__17192\,
            lcout => \POWERLED.func_state_ns_0_i_o3_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO2TE_9_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15145\,
            in2 => \_gnd_net_\,
            in3 => \N__15893\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_39_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI34C41_8_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__17268\,
            in1 => \N__15690\,
            in2 => \N__15104\,
            in3 => \N__17191\,
            lcout => \POWERLED.dutycycle_RNI34C41Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9K371_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__18563\,
            in1 => \N__18506\,
            in2 => \N__16952\,
            in3 => \N__16642\,
            lcout => \POWERLED.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIP0P11_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__15038\,
            in1 => \N__15017\,
            in2 => \N__14999\,
            in3 => \N__15488\,
            lcout => \POWERLED.func_state_ns_0_i_o2_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI16B71_5_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__15455\,
            in1 => \N__16063\,
            in2 => \N__16436\,
            in3 => \N__16219\,
            lcout => \POWERLED.dutycycle_RNI16B71Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__17392\,
            in1 => \N__16829\,
            in2 => \N__17108\,
            in3 => \N__17291\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18193\,
            ce => \N__17660\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIVCSK_5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16417\,
            in2 => \N__16226\,
            in3 => \N__17131\,
            lcout => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNINT777_1_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__18339\,
            in1 => \N__16644\,
            in2 => \N__17020\,
            in3 => \N__15422\,
            lcout => OPEN,
            ltout => \POWERLED.N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9LUBC_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__17033\,
            in1 => \N__18341\,
            in2 => \N__15404\,
            in3 => \N__16356\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI95RKL_8_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__17083\,
            in1 => \N__15347\,
            in2 => \N__15401\,
            in3 => \N__17954\,
            lcout => \POWERLED.count_clk_RNI95RKLZ0Z_8\,
            ltout => \POWERLED.count_clk_RNI95RKLZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_RNO_0_15_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__17955\,
            in1 => \_gnd_net_\,
            in2 => \N__15362\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_39_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI1J0G7_8_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__18340\,
            in1 => \N__15978\,
            in2 => \N__17021\,
            in3 => \N__15944\,
            lcout => \POWERLED.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNI8MSK_5_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15565\,
            in2 => \N__17135\,
            in3 => \N__17195\,
            lcout => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4I7Q_0_5_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16223\,
            in1 => \N__16139\,
            in2 => \N__16026\,
            in3 => \N__16079\,
            lcout => \POWERLED.dutycycle_cnst_1_i_o2_0_a3_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__17391\,
            in1 => \N__16830\,
            in2 => \N__17100\,
            in3 => \N__15914\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18198\,
            ce => \N__17659\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6NI81_5_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16015\,
            in1 => \N__15892\,
            in2 => \N__15841\,
            in3 => \N__16078\,
            lcout => \POWERLED.dutycycle_RNI6NI81Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIK4I81_6_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__15808\,
            in1 => \N__16014\,
            in2 => \N__16437\,
            in3 => \N__15620\,
            lcout => \POWERLED.dutycycle_RNIK4I81Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIUUB41_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__16013\,
            in1 => \N__15686\,
            in2 => \N__15768\,
            in3 => \N__17201\,
            lcout => \POWERLED.un1_dutycycle_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEJ021_4_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__15698\,
            in1 => \N__15621\,
            in2 => \N__15566\,
            in3 => \N__17114\,
            lcout => \POWERLED.dutycycle_RNIEJ021Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9HME_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16630\,
            lcout => OPEN,
            ltout => \POWERLED.N_173_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI22MP5_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111001"
        )
    port map (
            in0 => \N__18583\,
            in1 => \N__16928\,
            in2 => \N__15491\,
            in3 => \N__15940\,
            lcout => \POWERLED.N_84\,
            ltout => \POWERLED.N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNID041B_8_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110101"
        )
    port map (
            in0 => \N__18501\,
            in1 => \N__16357\,
            in2 => \N__16382\,
            in3 => \N__15950\,
            lcout => \POWERLED.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNILK689_8_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15980\,
            in1 => \N__16970\,
            in2 => \N__18278\,
            in3 => \N__16358\,
            lcout => \POWERLED.N_65_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4I7Q_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__16224\,
            in1 => \N__16147\,
            in2 => \N__16090\,
            in3 => \N__16022\,
            lcout => \POWERLED.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIN6N36_1_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15986\,
            in2 => \_gnd_net_\,
            in3 => \N__18502\,
            lcout => \POWERLED.un1_dutycycle_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI56JJ2_8_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18259\,
            in1 => \N__17010\,
            in2 => \N__16939\,
            in3 => \N__15979\,
            lcout => \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIAA8L4_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__15928\,
            in1 => \N__16780\,
            in2 => \N__18258\,
            in3 => \N__16770\,
            lcout => \POWERLED.N_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8QI11_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15929\,
            in2 => \_gnd_net_\,
            in3 => \N__18238\,
            lcout => OPEN,
            ltout => \POWERLED.N_196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8CGP4_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__18335\,
            in1 => \N__16645\,
            in2 => \N__15917\,
            in3 => \N__16772\,
            lcout => \POWERLED.N_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDSEE1_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__16646\,
            in1 => \N__18239\,
            in2 => \N__16881\,
            in3 => \N__18580\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2GLJ3_5_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16781\,
            in2 => \_gnd_net_\,
            in3 => \N__16771\,
            lcout => \POWERLED.N_120\,
            ltout => \POWERLED.N_120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIA3PQ4_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__16924\,
            in1 => \N__18334\,
            in2 => \N__16757\,
            in3 => \N__18243\,
            lcout => \POWERLED.N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIP49M5_1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__16869\,
            in1 => \N__17044\,
            in2 => \_gnd_net_\,
            in3 => \N__16746\,
            lcout => OPEN,
            ltout => \POWERLED.N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOG1PG_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__16812\,
            in2 => \N__16706\,
            in3 => \N__16686\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2KFU_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__18564\,
            in1 => \N__18510\,
            in2 => \_gnd_net_\,
            in3 => \N__16643\,
            lcout => \POWERLED.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16583\,
            in1 => \N__16475\,
            in2 => \N__16541\,
            in3 => \N__16526\,
            lcout => \ALL_SYS_PWRGD.N_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16481\,
            lcout => \ALL_SYS_PWRGD.m4_0_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__17396\,
            in1 => \N__17057\,
            in2 => \N__18511\,
            in3 => \N__16466\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18199\,
            ce => \N__17661\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_5_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__17090\,
            in1 => \N__17397\,
            in2 => \N__16835\,
            in3 => \N__17287\,
            lcout => \POWERLED.dutycycle_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18199\,
            ce => \N__17661\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM0TE_8_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17260\,
            in3 => \N__17184\,
            lcout => \POWERLED.un1_dutycycle_1_34_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIMOAE_5_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17194\,
            in3 => \N__17130\,
            lcout => \POWERLED.un1_dutycycle_1_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un45_slp_s3n_0_a6_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__16964\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18342\,
            lcout => \POWERLED.un45_slp_s3n\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_2_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__18584\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16963\,
            lcout => \POWERLED.N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI4PO32_8_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__18262\,
            in1 => \N__16870\,
            in2 => \N__17051\,
            in3 => \N__17012\,
            lcout => \POWERLED.un2_slp_s3n_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIABCI1_8_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__17011\,
            in1 => \N__18311\,
            in2 => \N__16962\,
            in3 => \N__18261\,
            lcout => \POWERLED.dutycycle_1_sqmuxa_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_RNIS4LI_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18497\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16953\,
            lcout => \VCCST_EN_c\,
            ltout => \VCCST_EN_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_0_0_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__18581\,
            in1 => \N__18254\,
            in2 => \N__16838\,
            in3 => \N__16813\,
            lcout => \POWERLED.func_state_ns_0_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_RNITA4N_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__18582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18496\,
            lcout => slp_s4n_signal_i_0,
            ltout => \slp_s4n_signal_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a3_0_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18437\,
            in3 => \N__18427\,
            lcout => \VPP_VDDQ.N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__18333\,
            in1 => \N__18284\,
            in2 => \N__18263\,
            in3 => \N__18277\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18204\,
            ce => \N__17655\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
