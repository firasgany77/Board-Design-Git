-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 14 2022 10:43:49

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : in std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : in std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__39838\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15747\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \b2v_inst36.countZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst36.count_2_10\ : std_logic;
signal \b2v_inst36.count_rst_9\ : std_logic;
signal \b2v_inst36.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_5_cascade_\ : std_logic;
signal \b2v_inst36.count_2_5\ : std_logic;
signal \b2v_inst36.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst36.count_2_4\ : std_logic;
signal \b2v_inst36.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst36.count_2_11\ : std_logic;
signal \b2v_inst36.count_2_6\ : std_logic;
signal \b2v_inst36.count_rst_6\ : std_logic;
signal \b2v_inst36.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_8_cascade_\ : std_logic;
signal \b2v_inst36.count_2_8\ : std_logic;
signal \b2v_inst36.count_rst_4\ : std_logic;
signal \b2v_inst36.count_rst_3\ : std_logic;
signal \b2v_inst36.count_rst_13\ : std_logic;
signal \b2v_inst36.count_rst_13_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_1\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_0_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_2\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_7\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_12_cascade_\ : std_logic;
signal \b2v_inst36.N_1_i_cascade_\ : std_logic;
signal \b2v_inst36.count_2_0\ : std_logic;
signal \b2v_inst36.count_rst_14\ : std_logic;
signal \b2v_inst36.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.count_2_1\ : std_logic;
signal \b2v_inst16.count_rst_0_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst16.count_4_11\ : std_logic;
signal \b2v_inst16.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst16.count_4_4\ : std_logic;
signal \b2v_inst16.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst16.count_4_3\ : std_logic;
signal \b2v_inst16.count_4_i_a3_9_0\ : std_logic;
signal \b2v_inst16.count_4_i_a3_8_0_cascade_\ : std_logic;
signal \b2v_inst16.count_4_i_a3_10_0\ : std_logic;
signal \b2v_inst16.N_414_cascade_\ : std_logic;
signal \b2v_inst16.N_416_cascade_\ : std_logic;
signal \b2v_inst16.count_rst_8\ : std_logic;
signal \b2v_inst16.count_RNIE4RF_2Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst16.count_rst_5_cascade_\ : std_logic;
signal \b2v_inst16.N_414\ : std_logic;
signal \b2v_inst16.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst16.count_4_0\ : std_logic;
signal \b2v_inst16.countZ0Z_1\ : std_logic;
signal \b2v_inst16.count_4_i_a3_7_0\ : std_logic;
signal \b2v_inst16.count_RNIE4RF_2Z0Z_1\ : std_logic;
signal \b2v_inst16.count_4_1\ : std_logic;
signal \b2v_inst16.countZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst16.count_4_7\ : std_logic;
signal \b2v_inst16.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst16.count_4_5\ : std_logic;
signal \b2v_inst16.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst16.count_4_8\ : std_logic;
signal \b2v_inst16.count_rst_12\ : std_logic;
signal \b2v_inst16.curr_state_7_0_1_cascade_\ : std_logic;
signal vddq_ok : std_logic;
signal \b2v_inst16.N_208_0_cascade_\ : std_logic;
signal \b2v_inst16.curr_state_RNIBO6I1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst16.curr_state_2_1\ : std_logic;
signal \b2v_inst16.curr_state_2_0\ : std_logic;
signal \b2v_inst11.count_0_7\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \b2v_inst11.un1_count_cry_1_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_cry_2_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_cry_5\ : std_logic;
signal \b2v_inst11.count_1_7\ : std_logic;
signal \b2v_inst11.un1_count_cry_6\ : std_logic;
signal \b2v_inst11.un1_count_cry_7\ : std_logic;
signal \b2v_inst11.un1_count_cry_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \b2v_inst11.un1_count_cry_9\ : std_logic;
signal \b2v_inst11.un1_count_cry_10\ : std_logic;
signal \b2v_inst11.un1_count_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_12\ : std_logic;
signal \b2v_inst11.un1_count_cry_13\ : std_logic;
signal \b2v_inst11.un1_count_cry_14\ : std_logic;
signal \b2v_inst11.count_1_5\ : std_logic;
signal \b2v_inst11.count_0_5\ : std_logic;
signal \b2v_inst11.count_1_14\ : std_logic;
signal \b2v_inst11.count_0_14\ : std_logic;
signal \b2v_inst11.count_1_6\ : std_logic;
signal \b2v_inst11.count_0_6\ : std_logic;
signal \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\ : std_logic;
signal \b2v_inst11.count_0_15\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_0\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_1\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_2\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_3\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_4\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_5\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_6\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_7\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_8\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_9\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_10\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_11\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_12\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_13\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_cry_14\ : std_logic;
signal \b2v_inst11.un85_clk_100khz0\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \b2v_inst36.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_12\ : std_logic;
signal \b2v_inst36.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_3\ : std_logic;
signal \b2v_inst36.count_rst_11\ : std_logic;
signal \b2v_inst36.count_2_2\ : std_logic;
signal \b2v_inst36.count_2_3\ : std_logic;
signal \b2v_inst36.count_2_7\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_1\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_2\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst36.countZ0Z_3\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_4\ : std_logic;
signal \b2v_inst36.count_rst_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_5\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_6\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_5_c_RNIE2FZ0Z8\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst36.countZ0Z_7\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_8\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_8\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \b2v_inst36.countZ0Z_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst36.countZ0Z_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst36.count_2_12\ : std_logic;
signal \b2v_inst36.count_rst_2\ : std_logic;
signal \b2v_inst36.countZ0Z_12\ : std_logic;
signal \b2v_inst36.count_rst_5\ : std_logic;
signal \b2v_inst36.countZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst36.count_2_9\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_6\ : std_logic;
signal \b2v_inst36.countZ0Z_14\ : std_logic;
signal \b2v_inst36.countZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_0\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_10\ : std_logic;
signal \b2v_inst36.count_2_13\ : std_logic;
signal \b2v_inst36.count_rst_1\ : std_logic;
signal \b2v_inst36.countZ0Z_13\ : std_logic;
signal \b2v_inst36.count_rst_0\ : std_logic;
signal \b2v_inst36.count_2_14\ : std_logic;
signal \b2v_inst36.curr_state_RNINSDSZ0Z_0\ : std_logic;
signal \b2v_inst36.count_rst\ : std_logic;
signal \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.count_2_15\ : std_logic;
signal \b2v_inst36.countZ0Z_15\ : std_logic;
signal \b2v_inst16.count_en_cascade_\ : std_logic;
signal \b2v_inst16.un4_count_1_axb_1\ : std_logic;
signal \b2v_inst16.countZ0Z_0\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \b2v_inst16.countZ0Z_2\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_1\ : std_logic;
signal \b2v_inst16.countZ0Z_3\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2\ : std_logic;
signal \b2v_inst16.countZ0Z_4\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3\ : std_logic;
signal \b2v_inst16.countZ0Z_5\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4\ : std_logic;
signal \b2v_inst16.countZ0Z_6\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_5\ : std_logic;
signal \b2v_inst16.countZ0Z_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_9\ : std_logic;
signal \b2v_inst16.countZ0Z_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_12\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_13\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_14\ : std_logic;
signal \b2v_inst16.countZ0Z_12\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst16.countZ0Z_8\ : std_logic;
signal \b2v_inst16.count_rst_13\ : std_logic;
signal \b2v_inst16.count_rst_14_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_9\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst16.countZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst16.N_416\ : std_logic;
signal \b2v_inst16.count_4_9\ : std_logic;
signal \b2v_inst16.count_4_10\ : std_logic;
signal \b2v_inst16.count_rst\ : std_logic;
signal \b2v_inst16.countZ0Z_10\ : std_logic;
signal \b2v_inst16.count_rst_1\ : std_logic;
signal \b2v_inst16.count_4_12\ : std_logic;
signal \b2v_inst11.curr_state_3_0_cascade_\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJZ0Z62\ : std_logic;
signal \b2v_inst11.curr_state_4_0\ : std_logic;
signal \b2v_inst11.count_0_0\ : std_logic;
signal \b2v_inst11.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_1_1_cascade_\ : std_logic;
signal \CONSTANT_ONE_NET_cascade_\ : std_logic;
signal \b2v_inst11.N_5852_i\ : std_logic;
signal \b2v_inst11.countZ0Z_1\ : std_logic;
signal \b2v_inst11.count_0_1\ : std_logic;
signal \b2v_inst11.count_0_8\ : std_logic;
signal \b2v_inst11.count_1_8\ : std_logic;
signal \b2v_inst11.count_1_9\ : std_logic;
signal \b2v_inst11.count_0_9\ : std_logic;
signal \b2v_inst11.count_1_10\ : std_logic;
signal \b2v_inst11.count_0_10\ : std_logic;
signal \b2v_inst11.count_1_11\ : std_logic;
signal \b2v_inst11.count_0_11\ : std_logic;
signal \b2v_inst11.count_1_2\ : std_logic;
signal \b2v_inst11.count_0_2\ : std_logic;
signal \b2v_inst11.count_1_12\ : std_logic;
signal \b2v_inst11.count_0_12\ : std_logic;
signal \b2v_inst11.count_1_3\ : std_logic;
signal \b2v_inst11.count_0_3\ : std_logic;
signal \b2v_inst11.count_1_13\ : std_logic;
signal \b2v_inst11.count_0_13\ : std_logic;
signal \b2v_inst11.count_1_4\ : std_logic;
signal \b2v_inst11.count_0_4\ : std_logic;
signal \b2v_inst11.countZ0Z_2\ : std_logic;
signal \b2v_inst11.countZ0Z_3\ : std_logic;
signal \b2v_inst11.countZ0Z_4\ : std_logic;
signal \b2v_inst11.countZ0Z_7\ : std_logic;
signal \b2v_inst11.countZ0Z_6\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlt6_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_5\ : std_logic;
signal \b2v_inst11.countZ0Z_10\ : std_logic;
signal \b2v_inst11.countZ0Z_12\ : std_logic;
signal \b2v_inst11.countZ0Z_11\ : std_logic;
signal \b2v_inst11.countZ0Z_13\ : std_logic;
signal \b2v_inst11.countZ0Z_14\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_15\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_3\ : std_logic;
signal \b2v_inst11.countZ0Z_8\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_9\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_8\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.curr_state_3_i_m2_0_rep1_1\ : std_logic;
signal \b2v_inst11.N_5853_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \b2v_inst11.N_5854_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_0\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_1\ : std_logic;
signal \b2v_inst11.N_5855_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_1\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_2\ : std_logic;
signal \b2v_inst11.N_5856_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_2\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_3\ : std_logic;
signal \b2v_inst11.N_5857_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_3\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_4\ : std_logic;
signal \b2v_inst11.N_5858_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_4\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_5\ : std_logic;
signal \b2v_inst11.N_5859_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_5\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_6\ : std_logic;
signal \b2v_inst11.N_5860_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_6\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_7\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_8\ : std_logic;
signal \b2v_inst11.N_5861_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0_7\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \b2v_inst11.N_5862_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_8\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_9\ : std_logic;
signal \b2v_inst11.N_5863_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_9\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_10\ : std_logic;
signal \b2v_inst11.N_5864_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_10\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_11\ : std_logic;
signal \b2v_inst11.N_5865_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_11\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_12\ : std_logic;
signal \b2v_inst11.N_5866_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_12\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_13\ : std_logic;
signal \b2v_inst11.N_5867_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_13\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1_cry_14\ : std_logic;
signal \b2v_inst11.un85_clk_100khz1\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i_0_8\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_1_cascade_\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_1_cascade_\ : std_logic;
signal \b2v_inst200.count_RNIZ0Z_1\ : std_logic;
signal \b2v_inst200.countZ0Z_16\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_0\ : std_logic;
signal \b2v_inst200.count_3_1\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_3_cascade_\ : std_logic;
signal \b2v_inst200.count_3_3\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_2\ : std_logic;
signal \b2v_inst200.count_3_13\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_5\ : std_logic;
signal \b2v_inst200.count_3_12\ : std_logic;
signal \b2v_inst200.count_3_9\ : std_logic;
signal \b2v_inst200.countZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_4\ : std_logic;
signal \b2v_inst200.count_3_5\ : std_logic;
signal \b2v_inst16.countZ0Z_15\ : std_logic;
signal \b2v_inst16.count_rst_4\ : std_logic;
signal \b2v_inst16.count_4_15\ : std_logic;
signal \b2v_inst16.countZ0Z_13\ : std_logic;
signal \b2v_inst16.count_rst_2\ : std_logic;
signal \b2v_inst16.count_4_13\ : std_logic;
signal \b2v_inst16.countZ0Z_14\ : std_logic;
signal \b2v_inst16.count_rst_3\ : std_logic;
signal \b2v_inst16.count_4_14\ : std_logic;
signal \b2v_inst16.count_rst_7\ : std_logic;
signal \b2v_inst16.count_4_2\ : std_logic;
signal \b2v_inst16.count_rst_11\ : std_logic;
signal \b2v_inst16.count_4_6\ : std_logic;
signal \b2v_inst16.count_en\ : std_logic;
signal \b2v_inst16.N_3037_i\ : std_logic;
signal \b2v_inst36.curr_state_0_1\ : std_logic;
signal \b2v_inst36.curr_state_7_1_cascade_\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst36.N_1_i\ : std_logic;
signal \b2v_inst36.curr_state_0_0\ : std_logic;
signal \b2v_inst36.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.count_0_sqmuxa\ : std_logic;
signal \b2v_inst11.count_off_0_11\ : std_logic;
signal \b2v_inst11.count_off_0_10\ : std_logic;
signal \b2v_inst11.count_off_0_12\ : std_logic;
signal \b2v_inst11.count_off_0_3\ : std_logic;
signal \b2v_inst11.count_off_0_14\ : std_logic;
signal \b2v_inst11.count_offZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst11.count_off_0_13\ : std_logic;
signal \b2v_inst11.g0_i_o3_0\ : std_logic;
signal \b2v_inst11.un85_clk_100khz1_THRU_CO\ : std_logic;
signal \b2v_inst11.un85_clk_100khz0_THRU_CO\ : std_logic;
signal \b2v_inst11.N_6_cascade_\ : std_logic;
signal \b2v_inst11.g0_0_0_rep1_1\ : std_logic;
signal \b2v_inst11.pwm_outZ0\ : std_logic;
signal \b2v_inst11.g0_i_a3_0_1\ : std_logic;
signal \b2v_inst11.N_6\ : std_logic;
signal pwrbtn_led : std_logic;
signal \b2v_inst200.count_enZ0\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgd_en_cascade_\ : std_logic;
signal vpp_en : std_logic;
signal \b2v_inst16.curr_state_RNIBO6I1Z0Z_0\ : std_logic;
signal \b2v_inst16.N_268\ : std_logic;
signal \b2v_inst16.N_268_cascade_\ : std_logic;
signal \b2v_inst16.N_26\ : std_logic;
signal \b2v_inst11.countZ0Z_0\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i\ : std_logic;
signal \b2v_inst11.count_1_0\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_0\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2848\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_s_6\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i_0_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i_0_8\ : std_logic;
signal \b2v_inst16.N_208_0\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgd_en\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgdZ0\ : std_logic;
signal \b2v_inst200.count_1_0_cascade_\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_1\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \b2v_inst200.countZ0Z_2\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_3\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst200.countZ0Z_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_5\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_5_cZ0\ : std_logic;
signal \b2v_inst200.countZ0Z_7\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst200.countZ0Z_11\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst200.countZ0Z_12\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst200.countZ0Z_14\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_16\ : std_logic;
signal \b2v_inst200.count_1_16\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_15\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16\ : std_logic;
signal \b2v_inst200.countZ0Z_17\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\ : std_logic;
signal \b2v_inst200.count_0_17\ : std_logic;
signal \b2v_inst200.N_56_cascade_\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst200.m6_i_0_cascade_\ : std_logic;
signal \b2v_inst200.N_58_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \N_411\ : std_logic;
signal \N_411_cascade_\ : std_logic;
signal \b2v_inst200.m6_i_0\ : std_logic;
signal \b2v_inst200.curr_state_3_0\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_13\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12\ : std_logic;
signal \b2v_inst11.count_offZ0Z_14\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13\ : std_logic;
signal \b2v_inst11.count_offZ0Z_15\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14\ : std_logic;
signal \b2v_inst11.count_offZ0Z_12\ : std_logic;
signal \b2v_inst11.count_offZ0Z_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_10\ : std_logic;
signal \b2v_inst11.count_offZ0Z_9\ : std_logic;
signal \b2v_inst200.curr_state_i_2_cascade_\ : std_logic;
signal \b2v_inst200.i4_mux\ : std_logic;
signal \b2v_inst200.N_2989_i\ : std_logic;
signal \b2v_inst200.N_205_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_2\ : std_logic;
signal \b2v_inst200.HDA_SDO_ATP_0\ : std_logic;
signal \b2v_inst200.N_205\ : std_logic;
signal \b2v_inst200.curr_state_i_2\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \b2v_inst200.N_282\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst200.curr_state_3_1\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_1\ : std_logic;
signal \b2v_inst20.counter_1_cry_2\ : std_logic;
signal \b2v_inst20.counter_1_cry_3\ : std_logic;
signal \b2v_inst20.counter_1_cry_4\ : std_logic;
signal \b2v_inst20.counter_1_cry_5\ : std_logic;
signal \b2v_inst20.counter_1_cry_6\ : std_logic;
signal \b2v_inst20.counterZ0Z_8\ : std_logic;
signal \b2v_inst20.counter_1_cry_7\ : std_logic;
signal \b2v_inst20.counter_1_cry_8\ : std_logic;
signal \b2v_inst20.counterZ0Z_9\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_10\ : std_logic;
signal \b2v_inst20.counter_1_cry_9\ : std_logic;
signal \b2v_inst20.counterZ0Z_11\ : std_logic;
signal \b2v_inst20.counter_1_cry_10\ : std_logic;
signal \b2v_inst20.counter_1_cry_11\ : std_logic;
signal \b2v_inst20.counter_1_cry_12\ : std_logic;
signal \b2v_inst20.counter_1_cry_13\ : std_logic;
signal \b2v_inst20.counter_1_cry_14\ : std_logic;
signal \b2v_inst20.counter_1_cry_15\ : std_logic;
signal \b2v_inst20.counter_1_cry_16\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_17\ : std_logic;
signal \b2v_inst20.counter_1_cry_18\ : std_logic;
signal \b2v_inst20.counterZ0Z_20\ : std_logic;
signal \b2v_inst20.counter_1_cry_19\ : std_logic;
signal \b2v_inst20.counterZ0Z_21\ : std_logic;
signal \b2v_inst20.counter_1_cry_20\ : std_logic;
signal \b2v_inst20.counterZ0Z_22\ : std_logic;
signal \b2v_inst20.counter_1_cry_21\ : std_logic;
signal \b2v_inst20.counterZ0Z_23\ : std_logic;
signal \b2v_inst20.counter_1_cry_22\ : std_logic;
signal \b2v_inst20.counter_1_cry_23\ : std_logic;
signal \b2v_inst20.counter_1_cry_24\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_25\ : std_logic;
signal \b2v_inst20.counter_1_cry_26\ : std_logic;
signal \b2v_inst20.counterZ0Z_28\ : std_logic;
signal \b2v_inst20.counter_1_cry_27\ : std_logic;
signal \b2v_inst20.counterZ0Z_29\ : std_logic;
signal \b2v_inst20.counter_1_cry_28\ : std_logic;
signal \b2v_inst20.counterZ0Z_30\ : std_logic;
signal \b2v_inst20.counter_1_cry_29\ : std_logic;
signal \b2v_inst20.counter_1_cry_30\ : std_logic;
signal \b2v_inst20.counterZ0Z_31\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i_0_8\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i_0_8\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_15\ : std_logic;
signal \b2v_inst200.un2_count_1_axb_8\ : std_logic;
signal \b2v_inst200.count_3_15\ : std_logic;
signal \b2v_inst200.countZ0Z_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71\ : std_logic;
signal \b2v_inst200.count_1_8\ : std_logic;
signal \b2v_inst200.count_3_8\ : std_logic;
signal \b2v_inst200.countZ0Z_10\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_14\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_6\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_7_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_13\ : std_logic;
signal \b2v_inst200.count_RNI5RUP8Z0Z_8\ : std_logic;
signal \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_0\ : std_logic;
signal \b2v_inst200.count_3_0\ : std_logic;
signal \b2v_inst200.count_1_11\ : std_logic;
signal \b2v_inst200.count_3_11\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\ : std_logic;
signal \b2v_inst200.count_3_14\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\ : std_logic;
signal \b2v_inst200.count_3_2\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\ : std_logic;
signal \b2v_inst200.count_3_4\ : std_logic;
signal \b2v_inst200.count_1_6\ : std_logic;
signal \b2v_inst200.count_3_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\ : std_logic;
signal \b2v_inst200.count_3_7\ : std_logic;
signal \b2v_inst200.count_1_10\ : std_logic;
signal \b2v_inst200.count_3_10\ : std_logic;
signal \b2v_inst200.count_en_g\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_0\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst5.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst5.count_rst_6\ : std_logic;
signal \b2v_inst5.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_8_cascade_\ : std_logic;
signal \b2v_inst5.count_1_8\ : std_logic;
signal \b2v_inst5.count_rst_10\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst5.countZ0Z_4\ : std_logic;
signal \b2v_inst5.count_1_4\ : std_logic;
signal \b2v_inst11.count_off_0_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\ : std_logic;
signal \b2v_inst11.count_off_0_0\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_1\ : std_logic;
signal \b2v_inst11.count_off_0_1\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_offZ0Z_1\ : std_logic;
signal \b2v_inst11.count_offZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_offZ0Z_2\ : std_logic;
signal \b2v_inst20.counterZ0Z_7\ : std_logic;
signal \b2v_inst20.counter_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_5\ : std_logic;
signal \b2v_inst20.counter_1_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_6\ : std_logic;
signal \b2v_inst11.count_offZ0Z_3\ : std_logic;
signal \b2v_inst20.counterZ0Z_1\ : std_logic;
signal v33dsw_ok : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.count_offZ0Z_4\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\ : std_logic;
signal \b2v_inst11.count_off_0_4\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\ : std_logic;
signal \b2v_inst11.count_off_0_15\ : std_logic;
signal \b2v_inst11.count_off_0_5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\ : std_logic;
signal \b2v_inst11.count_offZ0Z_5\ : std_logic;
signal \b2v_inst11.count_off_0_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\ : std_logic;
signal \b2v_inst11.count_offZ0Z_6\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \b2v_inst20.un4_counter_1_and\ : std_logic;
signal \b2v_inst20.un4_counter_0\ : std_logic;
signal \b2v_inst20.un4_counter_2_and\ : std_logic;
signal \b2v_inst20.un4_counter_1\ : std_logic;
signal \b2v_inst20.un4_counter_2\ : std_logic;
signal \b2v_inst20.un4_counter_3\ : std_logic;
signal \b2v_inst20.un4_counter_5_and\ : std_logic;
signal \b2v_inst20.un4_counter_4\ : std_logic;
signal \b2v_inst20.un4_counter_5\ : std_logic;
signal \b2v_inst20.un4_counter_7_and\ : std_logic;
signal \b2v_inst20.un4_counter_6\ : std_logic;
signal b2v_inst20_un4_counter_7 : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_16\ : std_logic;
signal \b2v_inst20.counterZ0Z_17\ : std_logic;
signal \b2v_inst20.counterZ0Z_18\ : std_logic;
signal \b2v_inst20.counterZ0Z_19\ : std_logic;
signal \b2v_inst20.un4_counter_4_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_15\ : std_logic;
signal \b2v_inst20.counterZ0Z_13\ : std_logic;
signal \b2v_inst20.counterZ0Z_14\ : std_logic;
signal \b2v_inst20.counterZ0Z_12\ : std_logic;
signal \b2v_inst20.un4_counter_3_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_24\ : std_logic;
signal \b2v_inst20.counterZ0Z_26\ : std_logic;
signal \b2v_inst20.counterZ0Z_25\ : std_logic;
signal \b2v_inst20.counterZ0Z_27\ : std_logic;
signal \b2v_inst20.un4_counter_6_and\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_axb_6\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_s_7\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_i\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_axb_4_l_fx\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_axb_7_l_fx\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_axb_7\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i\ : std_logic;
signal pch_pwrok : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i_0_8\ : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i_0_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_4_c_RNIPKTZ0Z9\ : std_logic;
signal \b2v_inst5.count_1_5\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9\ : std_logic;
signal \b2v_inst5.count_1_6\ : std_logic;
signal \b2v_inst5.countZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst5.count_1_13\ : std_logic;
signal \b2v_inst5.countZ0Z_3\ : std_logic;
signal \b2v_inst5.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_1\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_0_c_RNILCPZ0Z9\ : std_logic;
signal \b2v_inst5.count_1_1\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2\ : std_logic;
signal \b2v_inst5.count_1_12\ : std_logic;
signal \b2v_inst5.count_1_14\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\ : std_logic;
signal \b2v_inst5.countZ0Z_14\ : std_logic;
signal \b2v_inst5.countZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_12\ : std_logic;
signal \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_0\ : std_logic;
signal \b2v_inst5.curr_state_0_1\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst5.count_1_0\ : std_logic;
signal \b2v_inst5.count_rst_14\ : std_logic;
signal \b2v_inst5.count_i_0\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst5.count_1_15\ : std_logic;
signal \b2v_inst5.count_rst\ : std_logic;
signal \b2v_inst5.countZ0Z_15\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.N_51\ : std_logic;
signal \b2v_inst5.m4_0\ : std_logic;
signal \curr_state_RNID8DP1_0_0_cascade_\ : std_logic;
signal \N_413\ : std_logic;
signal \b2v_inst5.curr_state_0_0\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst5.N_2856_i\ : std_logic;
signal \b2v_inst5.curr_state_RNIZ0Z_1\ : std_logic;
signal \b2v_inst5.N_2856_i_cascade_\ : std_logic;
signal \b2v_inst11.count_off_0_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\ : std_logic;
signal \b2v_inst11.count_offZ0Z_7\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_11\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_9\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_10\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_8\ : std_logic;
signal \b2v_inst11.count_off_RNI_1Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m0_0_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\ : std_logic;
signal \b2v_inst11.count_off_0_8\ : std_logic;
signal \b2v_inst11.count_offZ0Z_8\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\ : std_logic;
signal \b2v_inst11.count_off_0_9\ : std_logic;
signal \b2v_inst11.N_76_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNICMPB4Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_1_m2_1_cascade_\ : std_logic;
signal \b2v_inst11.func_state_cascade_\ : std_logic;
signal \b2v_inst11.N_339\ : std_logic;
signal \b2v_inst11.N_339_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI6IFF4Z0Z_1\ : std_logic;
signal \b2v_inst36.DSW_PWROK_0\ : std_logic;
signal \b2v_inst36.curr_state_RNI3E27Z0Z_0\ : std_logic;
signal dsw_pwrok : std_logic;
signal \b2v_inst11.func_state_1_m2_1\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_1\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_51_and_i_a3_0_1_cascade_\ : std_logic;
signal vpp_ok : std_logic;
signal \VCCST_EN_i_0_o3_0_cascade_\ : std_logic;
signal vddq_en : std_logic;
signal \b2v_inst11.count_clk_en_0_xZ0Z1_cascade_\ : std_logic;
signal \b2v_inst11.N_335\ : std_logic;
signal \v5s_enn_cascade_\ : std_logic;
signal \b2v_inst20.counterZ0Z_0\ : std_logic;
signal \b2v_inst20.un4_counter_0_and\ : std_logic;
signal \b2v_inst20.counter_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_2\ : std_logic;
signal \b2v_inst20.counter_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_3\ : std_logic;
signal \b2v_inst20.counter_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVKZ0_cascade_\ : std_logic;
signal \b2v_inst11.N_236\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\ : std_logic;
signal \b2v_inst11.N_295\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i\ : std_logic;
signal \b2v_inst11.N_3055_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_14Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m3_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_0\ : std_logic;
signal \b2v_inst11.N_19_i_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m0_ns_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m0\ : std_logic;
signal \b2v_inst11.g0_4_1_cascade_\ : std_logic;
signal \b2v_inst11.N_293_0\ : std_logic;
signal \b2v_inst11.g0_3_2_0\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_a2_1_4_cascade_\ : std_logic;
signal \b2v_inst11.N_363_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_s_3_sf\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_7\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_i_1\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_i_8\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_0_8\ : std_logic;
signal \b2v_inst6.count_rst_11_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_3_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_11\ : std_logic;
signal \b2v_inst6.count_0_3\ : std_logic;
signal \b2v_inst6.count_rst_10\ : std_logic;
signal \b2v_inst6.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst6.count_0_4\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_11\ : std_logic;
signal \b2v_inst5.count_1_7\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_6_c_RNIROVZ0Z9\ : std_logic;
signal \b2v_inst5.countZ0Z_7\ : std_logic;
signal \b2v_inst5.count_rst_3\ : std_logic;
signal \b2v_inst5.count_1_11\ : std_logic;
signal \b2v_inst5.countZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_1_c_RNIMEQZ0Z9\ : std_logic;
signal \b2v_inst5.count_1_2\ : std_logic;
signal \b2v_inst5.countZ0Z_2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\ : std_logic;
signal \b2v_inst5.count_1_3\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_10_cascade_\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_9\ : std_logic;
signal \b2v_inst5.countZ0Z_5\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_1\ : std_logic;
signal \b2v_inst5.countZ0Z_6\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_10\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst5.count_rst_4\ : std_logic;
signal \b2v_inst5.count_1_10\ : std_logic;
signal \b2v_inst5.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_4\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_11\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_5_cascade_\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_12\ : std_logic;
signal \b2v_inst5.N_1_i_cascade_\ : std_logic;
signal \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\ : std_logic;
signal \b2v_inst5.count_1_9\ : std_logic;
signal \b2v_inst5.countZ0Z_13\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12_THRU_CO\ : std_logic;
signal \b2v_inst5.count_rst_1\ : std_logic;
signal \b2v_inst5.N_1_i\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst5.countZ0Z_9\ : std_logic;
signal \b2v_inst5.count_0_sqmuxa\ : std_logic;
signal \b2v_inst5.count_rst_5\ : std_logic;
signal v33a_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal v1p8a_ok : std_logic;
signal v5a_ok : std_logic;
signal vr_ready_vccinaux : std_logic;
signal vr_ready_vccin : std_logic;
signal \b2v_inst6.N_192_cascade_\ : std_logic;
signal \b2v_inst6.N_241_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNIG8KAHZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1\ : std_logic;
signal \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.N_428_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNITV5AUZ0Z_7\ : std_logic;
signal \b2v_inst11.count_clk_RNILG61T1Z0Z_5\ : std_logic;
signal \b2v_inst11.un1_func_state25_4_i_a2_sxZ0_cascade_\ : std_logic;
signal \rsmrstn_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_0_2\ : std_logic;
signal \b2v_inst20_un4_counter_7_THRU_CO\ : std_logic;
signal \b2v_inst11.func_state_1_ss0_i_0_o3_0\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_331_N\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_a3_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_332_N\ : std_logic;
signal \b2v_inst11.func_state_RNI_2Z0Z_1\ : std_logic;
signal \b2v_inst11.N_337_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m2s2_i_1\ : std_logic;
signal \b2v_inst11.N_76\ : std_logic;
signal \b2v_inst11.func_state_RNI6IFF4_0Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_1_m2_0_cascade_\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m2_0\ : std_logic;
signal \VCCST_EN_i_0_o3_0\ : std_logic;
signal \b2v_inst11.func_stateZ1Z_0\ : std_logic;
signal \b2v_inst11.count_clk_en_0\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_3_1\ : std_logic;
signal \b2v_inst11.d_N_5\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_5_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.N_293\ : std_logic;
signal \b2v_inst11.N_365\ : std_logic;
signal \b2v_inst11.N_159_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_9Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m3_d_ns_1_0_cascade_\ : std_logic;
signal \b2v_inst11.g1_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNIDQ4A1Z0Z_5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m4_rn_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_11Z0Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m4_rn_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m4\ : std_logic;
signal \b2v_inst11.N_3057_0\ : std_logic;
signal \b2v_inst11.g1_0_0_0\ : std_logic;
signal \b2v_inst11.N_3055_0_0\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.g0_0_1\ : std_logic;
signal \b2v_inst11.g1_0_1_0\ : std_logic;
signal \b2v_inst11.g0_3_2\ : std_logic;
signal \b2v_inst11.g2_1_0_1_cascade_\ : std_logic;
signal \b2v_inst11.g2_1_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_10Z0Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNIPKS23Z0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08UZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNI5AV24Z0Z_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNIPKS23Z0Z_4\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.un1_i3_mux_cascade_\ : std_logic;
signal \b2v_inst11.d_i3_mux\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_0\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_0\ : std_logic;
signal \b2v_inst11.mult1_un138_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_2\ : std_logic;
signal \b2v_inst11.mult1_un131_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_2\ : std_logic;
signal \b2v_inst11.mult1_un124_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_2\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un110_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un103_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un96_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_7\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_9\ : std_logic;
signal \b2v_inst11.mult1_un68_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_11\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \b2v_inst11.CO2\ : std_logic;
signal \b2v_inst11.mult1_un61_sum\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_13\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_6\ : std_logic;
signal \b2v_inst11.mult1_un89_sum\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_8_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_9_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_6\ : std_logic;
signal \b2v_inst6.count_rst_5\ : std_logic;
signal \b2v_inst6.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst6.count_0_9\ : std_logic;
signal \b2v_inst6.count_0_8\ : std_logic;
signal \N_607_g\ : std_logic;
signal \b2v_inst6.N_394_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_1_1\ : std_logic;
signal \b2v_inst6.m6_i_a3_cascade_\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_1_0\ : std_logic;
signal \b2v_inst6.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst6.count_RNICV5H1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\ : std_logic;
signal \N_222\ : std_logic;
signal \b2v_inst6.N_2992_i_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_8\ : std_logic;
signal v5s_ok : std_logic;
signal v33s_ok : std_logic;
signal vccinaux_en : std_logic;
signal \b2v_inst6.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst6.curr_state_RNIKIRD1Z0Z_0\ : std_logic;
signal \b2v_inst6.N_276_0\ : std_logic;
signal \b2v_inst6.curr_state_RNIKIRD1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_ok_0\ : std_logic;
signal \b2v_inst6.N_2992_i\ : std_logic;
signal \b2v_inst6.N_3011_i\ : std_logic;
signal \b2v_inst6.N_192\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_1_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_0\ : std_logic;
signal \b2v_inst11.count_clk_0_1\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_1\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1\ : std_logic;
signal \b2v_inst11.N_379\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.N_190\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_3\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_3\ : std_logic;
signal \b2v_inst11.N_428\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\ : std_logic;
signal \b2v_inst11.func_state_1_m2_am_1_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNINCPR4Z0Z_0\ : std_logic;
signal \b2v_inst11.N_382\ : std_logic;
signal \b2v_inst11.N_315\ : std_logic;
signal vccst_en : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.count_clk_RNIG510TZ0Z_5\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_1\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_\ : std_logic;
signal \b2v_inst11.count_off_enZ0\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.N_382_N\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3_fast\ : std_logic;
signal \RSMRSTn_0\ : std_logic;
signal \b2v_inst11.g0_4_sx_cascade_\ : std_logic;
signal \curr_state_RNID8DP1_0_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0_0\ : std_logic;
signal \b2v_inst11.N_160_i\ : std_logic;
signal \b2v_inst11.N_160_i_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI5DLRZ0Z_0\ : std_logic;
signal \b2v_inst11.N_366\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_313_N\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2BZ0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_0\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_8Z0Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_2\ : std_logic;
signal \b2v_inst11.N_19_i\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \b2v_inst11.N_186_i_cascade_\ : std_logic;
signal \b2v_inst11.N_309\ : std_logic;
signal \b2v_inst11.un1_dutycycle_96_0_a3_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_25_and_i_0_1_0\ : std_logic;
signal \b2v_inst11.N_186_i\ : std_logic;
signal \b2v_inst11.N_117_f0_1\ : std_logic;
signal v5s_enn : std_logic;
signal \b2v_inst11.N_117_f0_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_2\ : std_logic;
signal \b2v_inst11.N_73\ : std_logic;
signal \b2v_inst11.dutycycle_eena_1\ : std_logic;
signal \b2v_inst11.N_159\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.N_363\ : std_logic;
signal \b2v_inst11.func_state_RNI_1Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_7_cascade_\ : std_logic;
signal \b2v_inst11.N_2943_i\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1Z0Z_1\ : std_logic;
signal \b2v_inst11.N_360_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\ : std_logic;
signal \b2v_inst11.N_234_N\ : std_logic;
signal \b2v_inst11.dutycycle_eena_9\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_12\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_eena_7\ : std_logic;
signal \b2v_inst11.N_6_0\ : std_logic;
signal \b2v_inst11.N_8_cascade_\ : std_logic;
signal \b2v_inst11.N_355\ : std_logic;
signal \b2v_inst11.g0_6_a5_0_0_cascade_\ : std_logic;
signal \b2v_inst11.g0_6_a5_2_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_7\ : std_logic;
signal \b2v_inst11.CO2_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_axb_6_i_l_fx\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_axb_5_i_l_ofx\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_2\ : std_logic;
signal \b2v_inst11.mult1_un47_sum1_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_15\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_6\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_15\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_10\ : std_logic;
signal \b2v_inst11.N_11_cascade_\ : std_logic;
signal \b2v_inst11.N_35_0\ : std_logic;
signal \b2v_inst11.N_13_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_11\ : std_logic;
signal \b2v_inst11.g0_6_a5_1_0\ : std_logic;
signal \b2v_inst6.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_7_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_3_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst6.count_0_11\ : std_logic;
signal \b2v_inst6.N_394\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_4\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_8\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_13\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_10\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_12\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_11\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o2_4_cascade_\ : std_logic;
signal \b2v_inst11.N_175\ : std_logic;
signal \b2v_inst11.count_clk_0_10\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_1\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_0\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_3\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_10\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_11\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_10_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_12\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_13\ : std_logic;
signal \b2v_inst11.func_state_RNIIGCET1_0_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14\ : std_logic;
signal \b2v_inst11.count_clk_1_11\ : std_logic;
signal \b2v_inst11.count_clk_0_11\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_7\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_8\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_8\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_9\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_9\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.N_369\ : std_logic;
signal \b2v_inst11.count_clk_en_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_14\ : std_logic;
signal \b2v_inst11.N_417\ : std_logic;
signal \b2v_inst11.func_state_RNID7Q51Z0Z_0\ : std_logic;
signal \b2v_inst11.count_off_RNI_1Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNI6M5R2Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_RNIJGA54Z0Z_1\ : std_logic;
signal \b2v_inst11.count_clk_1_14\ : std_logic;
signal \b2v_inst11.count_clk_0_14\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.N_2904_i_cascade_\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_s1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4_s1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_9Z0Z_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_s1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_s1\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_s1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10_s1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_s1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14_s1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_6\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EGZ0Z1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_11\ : std_logic;
signal \b2v_inst11.dutycycle_rst_6\ : std_logic;
signal \b2v_inst11.dutycycle\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_2\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_s0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3_s0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_10Z0Z_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_s0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_s0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_s0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_axb_15_s0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_15\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14_s0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_12_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_3_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_31_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_31\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_55_0_tz\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_14_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_14_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_9\ : std_logic;
signal \b2v_inst11.N_2904_i\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_12\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_9\ : std_logic;
signal \b2v_inst11.i2_mux_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_5\ : std_logic;
signal \b2v_inst11.un1_N_5_cascade_\ : std_logic;
signal \b2v_inst11.un1_i2_mux_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_11\ : std_logic;
signal \b2v_inst6.count_rst_7\ : std_logic;
signal \b2v_inst6.count_0_7\ : std_logic;
signal \b2v_inst6.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst6.count_RNICV5H1Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_1\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_1_cascade_\ : std_logic;
signal \b2v_inst6.count_RNICV5H1Z0Z_1\ : std_logic;
signal \b2v_inst6.countZ0Z_11\ : std_logic;
signal \b2v_inst6.count_0_1\ : std_logic;
signal \b2v_inst6.count_1_i_a3_4_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_6_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_3_0_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_5_0\ : std_logic;
signal \b2v_inst6.count_0_5\ : std_logic;
signal \b2v_inst6.count_rst_9\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_5\ : std_logic;
signal \b2v_inst6.count_0_14\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_13_c_RNIR6IOZ0Z5\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_14\ : std_logic;
signal \b2v_inst6.countZ0Z_14\ : std_logic;
signal \b2v_inst6.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_12_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_1_0_cascade_\ : std_logic;
signal \b2v_inst6.count_0_2\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_1_c_RNIN2PZ0Z3\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_2\ : std_logic;
signal \b2v_inst6.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_0_0_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_7_0\ : std_logic;
signal \b2v_inst6.count_0_6\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_6\ : std_logic;
signal \b2v_inst6.count_rst_2\ : std_logic;
signal \b2v_inst6.count_0_12\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_11_c_RNI8RABZ0\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_12\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_10\ : std_logic;
signal \b2v_inst6.count_0_10\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_9_c_RNIVIZ0Z14\ : std_logic;
signal \b2v_inst6.count_rst_4\ : std_logic;
signal \b2v_inst6.countZ0Z_15\ : std_logic;
signal \b2v_inst6.count_0_13\ : std_logic;
signal \b2v_inst6.countZ0Z_15_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_2_0\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0\ : std_logic;
signal \b2v_inst6.count_rst_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_12\ : std_logic;
signal \b2v_inst11.count_clk_1_12\ : std_logic;
signal \b2v_inst11.count_clk_0_12\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_13\ : std_logic;
signal \b2v_inst11.count_clk_1_13\ : std_logic;
signal \b2v_inst11.count_clk_0_13\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_5\ : std_logic;
signal \b2v_inst11.count_clk_0_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_5\ : std_logic;
signal \b2v_inst11.count_clk_0_7\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_7\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_axb_2\ : std_logic;
signal \b2v_inst11.count_clk_0_2\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_15\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\ : std_logic;
signal \b2v_inst11.count_clk_0_15\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_6\ : std_logic;
signal \b2v_inst11.count_clk_en\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_6\ : std_logic;
signal \b2v_inst6.N_241\ : std_logic;
signal \b2v_inst6.countZ0Z_0\ : std_logic;
signal \b2v_inst6.N_2994_i\ : std_logic;
signal \b2v_inst6.N_2994_i_cascade_\ : std_logic;
signal \b2v_inst6.N_389\ : std_logic;
signal \b2v_inst6.count_0_0\ : std_logic;
signal \b2v_inst6.count_rst\ : std_logic;
signal \b2v_inst6.count_0_15\ : std_logic;
signal \b2v_inst6.count_en\ : std_logic;
signal \b2v_inst6.curr_state_RNICV5H1Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNI_4Z0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_s0_sf\ : std_logic;
signal \b2v_inst11.count_clk_RNIG510TZ0Z_7\ : std_logic;
signal \b2v_inst11.N_305\ : std_logic;
signal \b2v_inst11.N_306\ : std_logic;
signal \b2v_inst11.N_231_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_13_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4\ : std_logic;
signal \b2v_inst11.dutycycle_0_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_13\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_6_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNILF063Z0Z_6\ : std_logic;
signal \b2v_inst11.N_172\ : std_logic;
signal \b2v_inst11.N_185\ : std_logic;
signal \b2v_inst11.dutycycle_set_1\ : std_logic;
signal \b2v_inst11.dutycycle_set_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_14_0\ : std_logic;
signal \b2v_inst11.dutycycle_0_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJZ0Z9\ : std_logic;
signal \b2v_inst11.dutycycle_RNIM98E2Z0Z_3\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNIM98E2Z0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_9\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3_rep1\ : std_logic;
signal \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_32_and_i_0_c_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_32_and_i_0_d\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_33_and_i_0_c_0_cascade_\ : std_logic;
signal \b2v_inst11.N_153_N\ : std_logic;
signal \b2v_inst11.N_155_N_cascade_\ : std_logic;
signal \b2v_inst11.g0_0_1_0_cascade_\ : std_logic;
signal \b2v_inst11.g0_1_1\ : std_logic;
signal \b2v_inst11.g3_0_0\ : std_logic;
signal rsmrstn : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.g1_0_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_36_and_i_0_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_0_7\ : std_logic;
signal \b2v_inst11.g0_0_1_0\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_0_7_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_13\ : std_logic;
signal \b2v_inst11.dutycycle_en_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_5\ : std_logic;
signal \b2v_inst11.N_302\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_6\ : std_logic;
signal \b2v_inst11.N_301\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0\ : std_logic;
signal \b2v_inst11.dutycycle_en_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_14\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_0_3_tz_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_eena_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_0_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3\ : std_logic;
signal \b2v_inst11.g1_i_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena_2\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_eena_2_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_30_and_i_0_0_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_10\ : std_logic;
signal \b2v_inst11.N_140_N\ : std_logic;
signal \b2v_inst11.N_425\ : std_logic;
signal \b2v_inst11.N_158_N_cascade_\ : std_logic;
signal \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\ : std_logic;
signal \b2v_inst11.dutycycle_en_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3AZ0Z64\ : std_logic;
signal \b2v_inst11.dutycycle_en_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_15\ : std_logic;
signal \b2v_inst11.N_326_N\ : std_logic;
signal fpga_osc : std_logic;
signal \b2v_inst11.N_224_iZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s1_8\ : std_logic;
signal \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_s0_8\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_eena_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1_cascade_\ : std_logic;
signal \G_149\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_6\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_i2_mux_0\ : std_logic;
signal \b2v_inst11.un1_N_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_12\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_8\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_s_9_sf_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_12\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_1\ : std_logic;
signal \b2v_inst11.N_371_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNIDUQ02Z0Z_1\ : std_logic;
signal \b2v_inst11.g2_0_0Z0Z_0\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \b2v_inst11.func_state\ : std_logic;
signal \b2v_inst11.g2_3Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.N_200_i\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_0\ : std_logic;
signal slp_s3n : std_logic;
signal slp_s4n : std_logic;
signal \b2v_inst11.N_161\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    \SUSWARN_N_wire\ <= SUSWARN_N;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    \VCCINAUX_VR_PE_wire\ <= VCCINAUX_VR_PE;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    \VCCIN_VR_PE_wire\ <= VCCIN_VR_PE;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39838\,
            DIN => \N__39837\,
            DOUT => \N__39836\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39838\,
            PADOUT => \N__39837\,
            PADIN => \N__39836\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccinaux,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39829\,
            DIN => \N__39828\,
            DOUT => \N__39827\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39829\,
            PADOUT => \N__39828\,
            PADIN => \N__39827\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39820\,
            DIN => \N__39819\,
            DOUT => \N__39818\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39820\,
            PADOUT => \N__39819\,
            PADIN => \N__39818\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39811\,
            DIN => \N__39810\,
            DOUT => \N__39809\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39811\,
            PADOUT => \N__39810\,
            PADIN => \N__39809\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24846\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39802\,
            DIN => \N__39801\,
            DOUT => \N__39800\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39802\,
            PADOUT => \N__39801\,
            PADIN => \N__39800\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39793\,
            DIN => \N__39792\,
            DOUT => \N__39791\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39793\,
            PADOUT => \N__39792\,
            PADIN => \N__39791\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39784\,
            DIN => \N__39783\,
            DOUT => \N__39782\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39784\,
            PADOUT => \N__39783\,
            PADIN => \N__39782\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39775\,
            DIN => \N__39774\,
            DOUT => \N__39773\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39775\,
            PADOUT => \N__39774\,
            PADIN => \N__39773\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39766\,
            DIN => \N__39765\,
            DOUT => \N__39764\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39766\,
            PADOUT => \N__39765\,
            PADIN => \N__39764\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29116\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39757\,
            DIN => \N__39756\,
            DOUT => \N__39755\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39757\,
            PADOUT => \N__39756\,
            PADIN => \N__39755\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39748\,
            DIN => \N__39747\,
            DOUT => \N__39746\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39748\,
            PADOUT => \N__39747\,
            PADIN => \N__39746\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39739\,
            DIN => \N__39738\,
            DOUT => \N__39737\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39739\,
            PADOUT => \N__39738\,
            PADIN => \N__39737\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19878\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39730\,
            DIN => \N__39729\,
            DOUT => \N__39728\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39730\,
            PADOUT => \N__39729\,
            PADIN => \N__39728\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39721\,
            DIN => \N__39720\,
            DOUT => \N__39719\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39721\,
            PADOUT => \N__39720\,
            PADIN => \N__39719\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39712\,
            DIN => \N__39711\,
            DOUT => \N__39710\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39712\,
            PADOUT => \N__39711\,
            PADIN => \N__39710\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39703\,
            DIN => \N__39702\,
            DOUT => \N__39701\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39703\,
            PADOUT => \N__39702\,
            PADIN => \N__39701\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39694\,
            DIN => \N__39693\,
            DOUT => \N__39692\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39694\,
            PADOUT => \N__39693\,
            PADIN => \N__39692\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27984\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39685\,
            DIN => \N__39684\,
            DOUT => \N__39683\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39685\,
            PADOUT => \N__39684\,
            PADIN => \N__39683\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39676\,
            DIN => \N__39675\,
            DOUT => \N__39674\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39676\,
            PADOUT => \N__39675\,
            PADIN => \N__39674\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39667\,
            DIN => \N__39666\,
            DOUT => \N__39665\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39667\,
            PADOUT => \N__39666\,
            PADIN => \N__39665\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39658\,
            DIN => \N__39657\,
            DOUT => \N__39656\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39658\,
            PADOUT => \N__39657\,
            PADIN => \N__39656\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39649\,
            DIN => \N__39648\,
            DOUT => \N__39647\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39649\,
            PADOUT => \N__39648\,
            PADIN => \N__39647\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39640\,
            DIN => \N__39639\,
            DOUT => \N__39638\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39640\,
            PADOUT => \N__39639\,
            PADIN => \N__39638\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39631\,
            DIN => \N__39630\,
            DOUT => \N__39629\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39631\,
            PADOUT => \N__39630\,
            PADIN => \N__39629\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39622\,
            DIN => \N__39621\,
            DOUT => \N__39620\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39622\,
            PADOUT => \N__39621\,
            PADIN => \N__39620\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34842\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39613\,
            DIN => \N__39612\,
            DOUT => \N__39611\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39613\,
            PADOUT => \N__39612\,
            PADIN => \N__39611\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39604\,
            DIN => \N__39603\,
            DOUT => \N__39602\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39604\,
            PADOUT => \N__39603\,
            PADIN => \N__39602\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23941\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39595\,
            DIN => \N__39594\,
            DOUT => \N__39593\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39595\,
            PADOUT => \N__39594\,
            PADIN => \N__39593\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23945\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39586\,
            DIN => \N__39585\,
            DOUT => \N__39584\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39586\,
            PADOUT => \N__39585\,
            PADIN => \N__39584\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39577\,
            DIN => \N__39576\,
            DOUT => \N__39575\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39577\,
            PADOUT => \N__39576\,
            PADIN => \N__39575\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39568\,
            DIN => \N__39567\,
            DOUT => \N__39566\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39568\,
            PADOUT => \N__39567\,
            PADIN => \N__39566\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39559\,
            DIN => \N__39558\,
            DOUT => \N__39557\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39559\,
            PADOUT => \N__39558\,
            PADIN => \N__39557\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39550\,
            DIN => \N__39549\,
            DOUT => \N__39548\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39550\,
            PADOUT => \N__39549\,
            PADIN => \N__39548\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39541\,
            DIN => \N__39540\,
            DOUT => \N__39539\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39541\,
            PADOUT => \N__39540\,
            PADIN => \N__39539\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21369\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39532\,
            DIN => \N__39531\,
            DOUT => \N__39530\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39532\,
            PADOUT => \N__39531\,
            PADIN => \N__39530\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39523\,
            DIN => \N__39522\,
            DOUT => \N__39521\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39523\,
            PADOUT => \N__39522\,
            PADIN => \N__39521\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19848\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39514\,
            DIN => \N__39513\,
            DOUT => \N__39512\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39514\,
            PADOUT => \N__39513\,
            PADIN => \N__39512\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39505\,
            DIN => \N__39504\,
            DOUT => \N__39503\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39505\,
            PADOUT => \N__39504\,
            PADIN => \N__39503\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39496\,
            DIN => \N__39495\,
            DOUT => \N__39494\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39496\,
            PADOUT => \N__39495\,
            PADIN => \N__39494\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39487\,
            DIN => \N__39486\,
            DOUT => \N__39485\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39487\,
            PADOUT => \N__39486\,
            PADIN => \N__39485\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39478\,
            DIN => \N__39477\,
            DOUT => \N__39476\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39478\,
            PADOUT => \N__39477\,
            PADIN => \N__39476\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27668\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39469\,
            DIN => \N__39468\,
            DOUT => \N__39467\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39469\,
            PADOUT => \N__39468\,
            PADIN => \N__39467\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39460\,
            DIN => \N__39459\,
            DOUT => \N__39458\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39460\,
            PADOUT => \N__39459\,
            PADIN => \N__39458\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29117\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39451\,
            DIN => \N__39450\,
            DOUT => \N__39449\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39451\,
            PADOUT => \N__39450\,
            PADIN => \N__39449\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39442\,
            DIN => \N__39441\,
            DOUT => \N__39440\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39442\,
            PADOUT => \N__39441\,
            PADIN => \N__39440\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24735\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39433\,
            DIN => \N__39432\,
            DOUT => \N__39431\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39433\,
            PADOUT => \N__39432\,
            PADIN => \N__39431\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30945\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39424\,
            DIN => \N__39423\,
            DOUT => \N__39422\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39424\,
            PADOUT => \N__39423\,
            PADIN => \N__39422\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39415\,
            DIN => \N__39414\,
            DOUT => \N__39413\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39415\,
            PADOUT => \N__39414\,
            PADIN => \N__39413\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39406\,
            DIN => \N__39405\,
            DOUT => \N__39404\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39406\,
            PADOUT => \N__39405\,
            PADIN => \N__39404\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39397\,
            DIN => \N__39396\,
            DOUT => \N__39395\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39397\,
            PADOUT => \N__39396\,
            PADIN => \N__39395\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39388\,
            DIN => \N__39387\,
            DOUT => \N__39386\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39388\,
            PADOUT => \N__39387\,
            PADIN => \N__39386\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27675\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39379\,
            DIN => \N__39378\,
            DOUT => \N__39377\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39379\,
            PADOUT => \N__39378\,
            PADIN => \N__39377\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39370\,
            DIN => \N__39369\,
            DOUT => \N__39368\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39370\,
            PADOUT => \N__39369\,
            PADIN => \N__39368\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39361\,
            DIN => \N__39360\,
            DOUT => \N__39359\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39361\,
            PADOUT => \N__39360\,
            PADIN => \N__39359\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39352\,
            DIN => \N__39351\,
            DOUT => \N__39350\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39352\,
            PADOUT => \N__39351\,
            PADIN => \N__39350\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39343\,
            DIN => \N__39342\,
            DOUT => \N__39341\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39343\,
            PADOUT => \N__39342\,
            PADIN => \N__39341\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39334\,
            DIN => \N__39333\,
            DOUT => \N__39332\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39334\,
            PADOUT => \N__39333\,
            PADIN => \N__39332\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39325\,
            DIN => \N__39324\,
            DOUT => \N__39323\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39325\,
            PADOUT => \N__39324\,
            PADIN => \N__39323\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23952\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39316\,
            DIN => \N__39315\,
            DOUT => \N__39314\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39316\,
            PADOUT => \N__39315\,
            PADIN => \N__39314\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__9172\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39289\
        );

    \I__9171\ : InMux
    port map (
            O => \N__39296\,
            I => \N__39289\
        );

    \I__9170\ : InMux
    port map (
            O => \N__39295\,
            I => \N__39277\
        );

    \I__9169\ : InMux
    port map (
            O => \N__39294\,
            I => \N__39274\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__39289\,
            I => \N__39269\
        );

    \I__9167\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39266\
        );

    \I__9166\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39263\
        );

    \I__9165\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39256\
        );

    \I__9164\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39256\
        );

    \I__9163\ : InMux
    port map (
            O => \N__39284\,
            I => \N__39256\
        );

    \I__9162\ : InMux
    port map (
            O => \N__39283\,
            I => \N__39249\
        );

    \I__9161\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39249\
        );

    \I__9160\ : InMux
    port map (
            O => \N__39281\,
            I => \N__39249\
        );

    \I__9159\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39246\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__39277\,
            I => \N__39243\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__39274\,
            I => \N__39240\
        );

    \I__9156\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39237\
        );

    \I__9155\ : InMux
    port map (
            O => \N__39272\,
            I => \N__39234\
        );

    \I__9154\ : Sp12to4
    port map (
            O => \N__39269\,
            I => \N__39231\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__39266\,
            I => \N__39224\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__39263\,
            I => \N__39224\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__39256\,
            I => \N__39224\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__39249\,
            I => \N__39219\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__39246\,
            I => \N__39219\
        );

    \I__9148\ : Span4Mux_v
    port map (
            O => \N__39243\,
            I => \N__39214\
        );

    \I__9147\ : Span4Mux_h
    port map (
            O => \N__39240\,
            I => \N__39214\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__39237\,
            I => \N__39209\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__39234\,
            I => \N__39209\
        );

    \I__9144\ : Span12Mux_v
    port map (
            O => \N__39231\,
            I => \N__39206\
        );

    \I__9143\ : Span4Mux_v
    port map (
            O => \N__39224\,
            I => \N__39203\
        );

    \I__9142\ : Span12Mux_v
    port map (
            O => \N__39219\,
            I => \N__39200\
        );

    \I__9141\ : Span4Mux_v
    port map (
            O => \N__39214\,
            I => \N__39195\
        );

    \I__9140\ : Span4Mux_v
    port map (
            O => \N__39209\,
            I => \N__39195\
        );

    \I__9139\ : Odrv12
    port map (
            O => \N__39206\,
            I => gpio_fpga_soc_4
        );

    \I__9138\ : Odrv4
    port map (
            O => \N__39203\,
            I => gpio_fpga_soc_4
        );

    \I__9137\ : Odrv12
    port map (
            O => \N__39200\,
            I => gpio_fpga_soc_4
        );

    \I__9136\ : Odrv4
    port map (
            O => \N__39195\,
            I => gpio_fpga_soc_4
        );

    \I__9135\ : InMux
    port map (
            O => \N__39186\,
            I => \N__39172\
        );

    \I__9134\ : CascadeMux
    port map (
            O => \N__39185\,
            I => \N__39162\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__39184\,
            I => \N__39155\
        );

    \I__9132\ : InMux
    port map (
            O => \N__39183\,
            I => \N__39147\
        );

    \I__9131\ : InMux
    port map (
            O => \N__39182\,
            I => \N__39147\
        );

    \I__9130\ : InMux
    port map (
            O => \N__39181\,
            I => \N__39147\
        );

    \I__9129\ : CascadeMux
    port map (
            O => \N__39180\,
            I => \N__39143\
        );

    \I__9128\ : CascadeMux
    port map (
            O => \N__39179\,
            I => \N__39140\
        );

    \I__9127\ : CascadeMux
    port map (
            O => \N__39178\,
            I => \N__39136\
        );

    \I__9126\ : CascadeMux
    port map (
            O => \N__39177\,
            I => \N__39133\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__39176\,
            I => \N__39129\
        );

    \I__9124\ : InMux
    port map (
            O => \N__39175\,
            I => \N__39124\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__39172\,
            I => \N__39121\
        );

    \I__9122\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39118\
        );

    \I__9121\ : InMux
    port map (
            O => \N__39170\,
            I => \N__39102\
        );

    \I__9120\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39102\
        );

    \I__9119\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39102\
        );

    \I__9118\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39102\
        );

    \I__9117\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39102\
        );

    \I__9116\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39102\
        );

    \I__9115\ : InMux
    port map (
            O => \N__39162\,
            I => \N__39102\
        );

    \I__9114\ : CascadeMux
    port map (
            O => \N__39161\,
            I => \N__39099\
        );

    \I__9113\ : CascadeMux
    port map (
            O => \N__39160\,
            I => \N__39096\
        );

    \I__9112\ : CascadeMux
    port map (
            O => \N__39159\,
            I => \N__39088\
        );

    \I__9111\ : InMux
    port map (
            O => \N__39158\,
            I => \N__39077\
        );

    \I__9110\ : InMux
    port map (
            O => \N__39155\,
            I => \N__39077\
        );

    \I__9109\ : InMux
    port map (
            O => \N__39154\,
            I => \N__39077\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__39147\,
            I => \N__39074\
        );

    \I__9107\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39061\
        );

    \I__9106\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39061\
        );

    \I__9105\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39061\
        );

    \I__9104\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39061\
        );

    \I__9103\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39061\
        );

    \I__9102\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39061\
        );

    \I__9101\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39048\
        );

    \I__9100\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39048\
        );

    \I__9099\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39045\
        );

    \I__9098\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39042\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39035\
        );

    \I__9096\ : Span4Mux_s2_h
    port map (
            O => \N__39121\,
            I => \N__39035\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__39118\,
            I => \N__39035\
        );

    \I__9094\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39032\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__39102\,
            I => \N__39029\
        );

    \I__9092\ : InMux
    port map (
            O => \N__39099\,
            I => \N__39022\
        );

    \I__9091\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39022\
        );

    \I__9090\ : InMux
    port map (
            O => \N__39095\,
            I => \N__39022\
        );

    \I__9089\ : InMux
    port map (
            O => \N__39094\,
            I => \N__39019\
        );

    \I__9088\ : CascadeMux
    port map (
            O => \N__39093\,
            I => \N__39016\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__39092\,
            I => \N__39013\
        );

    \I__9086\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39007\
        );

    \I__9085\ : InMux
    port map (
            O => \N__39088\,
            I => \N__39007\
        );

    \I__9084\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39002\
        );

    \I__9083\ : InMux
    port map (
            O => \N__39086\,
            I => \N__39002\
        );

    \I__9082\ : CascadeMux
    port map (
            O => \N__39085\,
            I => \N__38998\
        );

    \I__9081\ : InMux
    port map (
            O => \N__39084\,
            I => \N__38995\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__39077\,
            I => \N__38992\
        );

    \I__9079\ : Span4Mux_s2_v
    port map (
            O => \N__39074\,
            I => \N__38987\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__38987\
        );

    \I__9077\ : CascadeMux
    port map (
            O => \N__39060\,
            I => \N__38984\
        );

    \I__9076\ : InMux
    port map (
            O => \N__39059\,
            I => \N__38971\
        );

    \I__9075\ : InMux
    port map (
            O => \N__39058\,
            I => \N__38971\
        );

    \I__9074\ : InMux
    port map (
            O => \N__39057\,
            I => \N__38971\
        );

    \I__9073\ : InMux
    port map (
            O => \N__39056\,
            I => \N__38971\
        );

    \I__9072\ : InMux
    port map (
            O => \N__39055\,
            I => \N__38968\
        );

    \I__9071\ : InMux
    port map (
            O => \N__39054\,
            I => \N__38964\
        );

    \I__9070\ : InMux
    port map (
            O => \N__39053\,
            I => \N__38961\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__39048\,
            I => \N__38958\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__39045\,
            I => \N__38945\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__39042\,
            I => \N__38945\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__39035\,
            I => \N__38945\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__39032\,
            I => \N__38945\
        );

    \I__9064\ : Span4Mux_s2_h
    port map (
            O => \N__39029\,
            I => \N__38945\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__39022\,
            I => \N__38945\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__39019\,
            I => \N__38942\
        );

    \I__9061\ : InMux
    port map (
            O => \N__39016\,
            I => \N__38935\
        );

    \I__9060\ : InMux
    port map (
            O => \N__39013\,
            I => \N__38935\
        );

    \I__9059\ : InMux
    port map (
            O => \N__39012\,
            I => \N__38935\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__39007\,
            I => \N__38930\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__39002\,
            I => \N__38930\
        );

    \I__9056\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38925\
        );

    \I__9055\ : InMux
    port map (
            O => \N__38998\,
            I => \N__38925\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__38995\,
            I => \N__38918\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__38992\,
            I => \N__38918\
        );

    \I__9052\ : Span4Mux_v
    port map (
            O => \N__38987\,
            I => \N__38918\
        );

    \I__9051\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38913\
        );

    \I__9050\ : InMux
    port map (
            O => \N__38983\,
            I => \N__38913\
        );

    \I__9049\ : InMux
    port map (
            O => \N__38982\,
            I => \N__38910\
        );

    \I__9048\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38905\
        );

    \I__9047\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38905\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__38971\,
            I => \N__38900\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__38968\,
            I => \N__38900\
        );

    \I__9044\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38897\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__38964\,
            I => \N__38888\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__38961\,
            I => \N__38888\
        );

    \I__9041\ : Span4Mux_s2_h
    port map (
            O => \N__38958\,
            I => \N__38888\
        );

    \I__9040\ : Span4Mux_v
    port map (
            O => \N__38945\,
            I => \N__38888\
        );

    \I__9039\ : Span4Mux_v
    port map (
            O => \N__38942\,
            I => \N__38877\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__38935\,
            I => \N__38877\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__38930\,
            I => \N__38877\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__38925\,
            I => \N__38877\
        );

    \I__9035\ : Span4Mux_h
    port map (
            O => \N__38918\,
            I => \N__38877\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__38913\,
            I => \b2v_inst11.func_state\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__38910\,
            I => \b2v_inst11.func_state\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__38905\,
            I => \b2v_inst11.func_state\
        );

    \I__9031\ : Odrv12
    port map (
            O => \N__38900\,
            I => \b2v_inst11.func_state\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__38897\,
            I => \b2v_inst11.func_state\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__38888\,
            I => \b2v_inst11.func_state\
        );

    \I__9028\ : Odrv4
    port map (
            O => \N__38877\,
            I => \b2v_inst11.func_state\
        );

    \I__9027\ : CascadeMux
    port map (
            O => \N__38862\,
            I => \b2v_inst11.g2_3Z0Z_0_cascade_\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__38859\,
            I => \N__38855\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__38858\,
            I => \N__38852\
        );

    \I__9024\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38839\
        );

    \I__9023\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38839\
        );

    \I__9022\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38839\
        );

    \I__9021\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38836\
        );

    \I__9020\ : CascadeMux
    port map (
            O => \N__38849\,
            I => \N__38833\
        );

    \I__9019\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38828\
        );

    \I__9018\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38825\
        );

    \I__9017\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38822\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__38839\,
            I => \N__38819\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__38836\,
            I => \N__38816\
        );

    \I__9014\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38809\
        );

    \I__9013\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38804\
        );

    \I__9012\ : InMux
    port map (
            O => \N__38831\,
            I => \N__38804\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__38828\,
            I => \N__38798\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__38825\,
            I => \N__38791\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__38822\,
            I => \N__38791\
        );

    \I__9008\ : Span4Mux_v
    port map (
            O => \N__38819\,
            I => \N__38791\
        );

    \I__9007\ : Span4Mux_h
    port map (
            O => \N__38816\,
            I => \N__38788\
        );

    \I__9006\ : InMux
    port map (
            O => \N__38815\,
            I => \N__38781\
        );

    \I__9005\ : InMux
    port map (
            O => \N__38814\,
            I => \N__38781\
        );

    \I__9004\ : InMux
    port map (
            O => \N__38813\,
            I => \N__38781\
        );

    \I__9003\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38778\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38773\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__38804\,
            I => \N__38773\
        );

    \I__9000\ : InMux
    port map (
            O => \N__38803\,
            I => \N__38766\
        );

    \I__8999\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38766\
        );

    \I__8998\ : InMux
    port map (
            O => \N__38801\,
            I => \N__38766\
        );

    \I__8997\ : Span4Mux_h
    port map (
            O => \N__38798\,
            I => \N__38761\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__38791\,
            I => \N__38761\
        );

    \I__8995\ : Span4Mux_v
    port map (
            O => \N__38788\,
            I => \N__38758\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__38781\,
            I => \N__38749\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__38778\,
            I => \N__38749\
        );

    \I__8992\ : Span12Mux_s2_v
    port map (
            O => \N__38773\,
            I => \N__38749\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__38766\,
            I => \N__38749\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__38761\,
            I => \b2v_inst11.N_200_i\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__38758\,
            I => \b2v_inst11.N_200_i\
        );

    \I__8988\ : Odrv12
    port map (
            O => \N__38749\,
            I => \b2v_inst11.N_200_i\
        );

    \I__8987\ : CascadeMux
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__8986\ : InMux
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__8984\ : Odrv12
    port map (
            O => \N__38733\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_0\
        );

    \I__8983\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38726\
        );

    \I__8982\ : CascadeMux
    port map (
            O => \N__38729\,
            I => \N__38719\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__38726\,
            I => \N__38714\
        );

    \I__8980\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38711\
        );

    \I__8979\ : InMux
    port map (
            O => \N__38724\,
            I => \N__38708\
        );

    \I__8978\ : CascadeMux
    port map (
            O => \N__38723\,
            I => \N__38705\
        );

    \I__8977\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38697\
        );

    \I__8976\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38697\
        );

    \I__8975\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38697\
        );

    \I__8974\ : CascadeMux
    port map (
            O => \N__38717\,
            I => \N__38694\
        );

    \I__8973\ : Span4Mux_v
    port map (
            O => \N__38714\,
            I => \N__38688\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__38711\,
            I => \N__38688\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__38708\,
            I => \N__38685\
        );

    \I__8970\ : InMux
    port map (
            O => \N__38705\,
            I => \N__38680\
        );

    \I__8969\ : InMux
    port map (
            O => \N__38704\,
            I => \N__38680\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38671\
        );

    \I__8967\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38666\
        );

    \I__8966\ : InMux
    port map (
            O => \N__38693\,
            I => \N__38666\
        );

    \I__8965\ : Span4Mux_h
    port map (
            O => \N__38688\,
            I => \N__38659\
        );

    \I__8964\ : Span4Mux_h
    port map (
            O => \N__38685\,
            I => \N__38659\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__38680\,
            I => \N__38659\
        );

    \I__8962\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38652\
        );

    \I__8961\ : InMux
    port map (
            O => \N__38678\,
            I => \N__38652\
        );

    \I__8960\ : InMux
    port map (
            O => \N__38677\,
            I => \N__38652\
        );

    \I__8959\ : CascadeMux
    port map (
            O => \N__38676\,
            I => \N__38649\
        );

    \I__8958\ : CascadeMux
    port map (
            O => \N__38675\,
            I => \N__38646\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__38674\,
            I => \N__38642\
        );

    \I__8956\ : Span4Mux_v
    port map (
            O => \N__38671\,
            I => \N__38632\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__38666\,
            I => \N__38632\
        );

    \I__8954\ : Span4Mux_s3_h
    port map (
            O => \N__38659\,
            I => \N__38632\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__38652\,
            I => \N__38632\
        );

    \I__8952\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38627\
        );

    \I__8951\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38627\
        );

    \I__8950\ : InMux
    port map (
            O => \N__38645\,
            I => \N__38622\
        );

    \I__8949\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38622\
        );

    \I__8948\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38619\
        );

    \I__8947\ : Span4Mux_v
    port map (
            O => \N__38632\,
            I => \N__38616\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38608\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__38622\,
            I => \N__38608\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__38619\,
            I => \N__38608\
        );

    \I__8943\ : IoSpan4Mux
    port map (
            O => \N__38616\,
            I => \N__38605\
        );

    \I__8942\ : InMux
    port map (
            O => \N__38615\,
            I => \N__38602\
        );

    \I__8941\ : Span4Mux_v
    port map (
            O => \N__38608\,
            I => \N__38595\
        );

    \I__8940\ : Span4Mux_s1_h
    port map (
            O => \N__38605\,
            I => \N__38595\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__38602\,
            I => \N__38595\
        );

    \I__8938\ : Span4Mux_h
    port map (
            O => \N__38595\,
            I => \N__38592\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__38592\,
            I => \N__38584\
        );

    \I__8936\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38579\
        );

    \I__8935\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38579\
        );

    \I__8934\ : InMux
    port map (
            O => \N__38589\,
            I => \N__38572\
        );

    \I__8933\ : InMux
    port map (
            O => \N__38588\,
            I => \N__38572\
        );

    \I__8932\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38572\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__38584\,
            I => slp_s3n
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__38579\,
            I => slp_s3n
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__38572\,
            I => slp_s3n
        );

    \I__8928\ : CascadeMux
    port map (
            O => \N__38565\,
            I => \N__38557\
        );

    \I__8927\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38547\
        );

    \I__8926\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38547\
        );

    \I__8925\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38544\
        );

    \I__8924\ : InMux
    port map (
            O => \N__38561\,
            I => \N__38539\
        );

    \I__8923\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38539\
        );

    \I__8922\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38530\
        );

    \I__8921\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38530\
        );

    \I__8920\ : InMux
    port map (
            O => \N__38555\,
            I => \N__38530\
        );

    \I__8919\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38530\
        );

    \I__8918\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38518\
        );

    \I__8917\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38518\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38510\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__38544\,
            I => \N__38510\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__38539\,
            I => \N__38505\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__38530\,
            I => \N__38505\
        );

    \I__8912\ : InMux
    port map (
            O => \N__38529\,
            I => \N__38502\
        );

    \I__8911\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38499\
        );

    \I__8910\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38488\
        );

    \I__8909\ : InMux
    port map (
            O => \N__38526\,
            I => \N__38488\
        );

    \I__8908\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38488\
        );

    \I__8907\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38488\
        );

    \I__8906\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38488\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__38518\,
            I => \N__38485\
        );

    \I__8904\ : InMux
    port map (
            O => \N__38517\,
            I => \N__38477\
        );

    \I__8903\ : InMux
    port map (
            O => \N__38516\,
            I => \N__38477\
        );

    \I__8902\ : InMux
    port map (
            O => \N__38515\,
            I => \N__38477\
        );

    \I__8901\ : Span4Mux_v
    port map (
            O => \N__38510\,
            I => \N__38472\
        );

    \I__8900\ : Span4Mux_v
    port map (
            O => \N__38505\,
            I => \N__38472\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__38502\,
            I => \N__38469\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__38499\,
            I => \N__38466\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__38488\,
            I => \N__38463\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__38485\,
            I => \N__38460\
        );

    \I__8895\ : InMux
    port map (
            O => \N__38484\,
            I => \N__38457\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__38477\,
            I => \N__38454\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__38472\,
            I => \N__38447\
        );

    \I__8892\ : Span4Mux_s3_h
    port map (
            O => \N__38469\,
            I => \N__38447\
        );

    \I__8891\ : Span4Mux_h
    port map (
            O => \N__38466\,
            I => \N__38447\
        );

    \I__8890\ : IoSpan4Mux
    port map (
            O => \N__38463\,
            I => \N__38444\
        );

    \I__8889\ : Sp12to4
    port map (
            O => \N__38460\,
            I => \N__38439\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__38457\,
            I => \N__38439\
        );

    \I__8887\ : Span12Mux_s8_h
    port map (
            O => \N__38454\,
            I => \N__38436\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__38447\,
            I => \N__38433\
        );

    \I__8885\ : IoSpan4Mux
    port map (
            O => \N__38444\,
            I => \N__38430\
        );

    \I__8884\ : Span12Mux_s8_h
    port map (
            O => \N__38439\,
            I => \N__38427\
        );

    \I__8883\ : Odrv12
    port map (
            O => \N__38436\,
            I => slp_s4n
        );

    \I__8882\ : Odrv4
    port map (
            O => \N__38433\,
            I => slp_s4n
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__38430\,
            I => slp_s4n
        );

    \I__8880\ : Odrv12
    port map (
            O => \N__38427\,
            I => slp_s4n
        );

    \I__8879\ : CascadeMux
    port map (
            O => \N__38418\,
            I => \N__38413\
        );

    \I__8878\ : CascadeMux
    port map (
            O => \N__38417\,
            I => \N__38410\
        );

    \I__8877\ : CascadeMux
    port map (
            O => \N__38416\,
            I => \N__38405\
        );

    \I__8876\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38399\
        );

    \I__8875\ : InMux
    port map (
            O => \N__38410\,
            I => \N__38399\
        );

    \I__8874\ : InMux
    port map (
            O => \N__38409\,
            I => \N__38392\
        );

    \I__8873\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38392\
        );

    \I__8872\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38392\
        );

    \I__8871\ : InMux
    port map (
            O => \N__38404\,
            I => \N__38388\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__38399\,
            I => \N__38383\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38383\
        );

    \I__8868\ : CascadeMux
    port map (
            O => \N__38391\,
            I => \N__38380\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__38388\,
            I => \N__38377\
        );

    \I__8866\ : Span4Mux_h
    port map (
            O => \N__38383\,
            I => \N__38374\
        );

    \I__8865\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38371\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__38377\,
            I => \N__38368\
        );

    \I__8863\ : Sp12to4
    port map (
            O => \N__38374\,
            I => \N__38363\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38363\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__38368\,
            I => \N__38360\
        );

    \I__8860\ : Span12Mux_s10_v
    port map (
            O => \N__38363\,
            I => \N__38357\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__38360\,
            I => \b2v_inst11.N_161\
        );

    \I__8858\ : Odrv12
    port map (
            O => \N__38357\,
            I => \b2v_inst11.N_161\
        );

    \I__8857\ : CascadeMux
    port map (
            O => \N__38352\,
            I => \N__38348\
        );

    \I__8856\ : CascadeMux
    port map (
            O => \N__38351\,
            I => \N__38333\
        );

    \I__8855\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38321\
        );

    \I__8854\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38321\
        );

    \I__8853\ : InMux
    port map (
            O => \N__38346\,
            I => \N__38321\
        );

    \I__8852\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38316\
        );

    \I__8851\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38316\
        );

    \I__8850\ : CascadeMux
    port map (
            O => \N__38343\,
            I => \N__38313\
        );

    \I__8849\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38306\
        );

    \I__8848\ : CascadeMux
    port map (
            O => \N__38341\,
            I => \N__38303\
        );

    \I__8847\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38296\
        );

    \I__8846\ : InMux
    port map (
            O => \N__38339\,
            I => \N__38296\
        );

    \I__8845\ : InMux
    port map (
            O => \N__38338\,
            I => \N__38296\
        );

    \I__8844\ : InMux
    port map (
            O => \N__38337\,
            I => \N__38292\
        );

    \I__8843\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38287\
        );

    \I__8842\ : InMux
    port map (
            O => \N__38333\,
            I => \N__38287\
        );

    \I__8841\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38280\
        );

    \I__8840\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38280\
        );

    \I__8839\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38280\
        );

    \I__8838\ : InMux
    port map (
            O => \N__38329\,
            I => \N__38275\
        );

    \I__8837\ : InMux
    port map (
            O => \N__38328\,
            I => \N__38275\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__38321\,
            I => \N__38271\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38268\
        );

    \I__8834\ : InMux
    port map (
            O => \N__38313\,
            I => \N__38259\
        );

    \I__8833\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38259\
        );

    \I__8832\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38259\
        );

    \I__8831\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38259\
        );

    \I__8830\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38254\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__38306\,
            I => \N__38251\
        );

    \I__8828\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38248\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__38296\,
            I => \N__38245\
        );

    \I__8826\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38242\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38237\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__38287\,
            I => \N__38237\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__38280\,
            I => \N__38232\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__38275\,
            I => \N__38232\
        );

    \I__8821\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38229\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__38271\,
            I => \N__38220\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__38268\,
            I => \N__38220\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__38259\,
            I => \N__38220\
        );

    \I__8817\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38215\
        );

    \I__8816\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38215\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__38254\,
            I => \N__38204\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__38251\,
            I => \N__38204\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38204\
        );

    \I__8812\ : Span4Mux_s1_v
    port map (
            O => \N__38245\,
            I => \N__38204\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38204\
        );

    \I__8810\ : Span4Mux_v
    port map (
            O => \N__38237\,
            I => \N__38197\
        );

    \I__8809\ : Span4Mux_v
    port map (
            O => \N__38232\,
            I => \N__38197\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__38229\,
            I => \N__38197\
        );

    \I__8807\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38194\
        );

    \I__8806\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38191\
        );

    \I__8805\ : Span4Mux_v
    port map (
            O => \N__38220\,
            I => \N__38188\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__38215\,
            I => \N__38183\
        );

    \I__8803\ : Span4Mux_v
    port map (
            O => \N__38204\,
            I => \N__38183\
        );

    \I__8802\ : Span4Mux_v
    port map (
            O => \N__38197\,
            I => \N__38180\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__38194\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__38191\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__38188\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__38183\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__38180\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__38169\,
            I => \N__38163\
        );

    \I__8795\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38155\
        );

    \I__8794\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38145\
        );

    \I__8793\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38145\
        );

    \I__8792\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38145\
        );

    \I__8791\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38145\
        );

    \I__8790\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38140\
        );

    \I__8789\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38140\
        );

    \I__8788\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38137\
        );

    \I__8787\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38132\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__38155\,
            I => \N__38127\
        );

    \I__8785\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38124\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__38145\,
            I => \N__38118\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38115\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__38137\,
            I => \N__38112\
        );

    \I__8781\ : InMux
    port map (
            O => \N__38136\,
            I => \N__38109\
        );

    \I__8780\ : CascadeMux
    port map (
            O => \N__38135\,
            I => \N__38103\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__38132\,
            I => \N__38100\
        );

    \I__8778\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38095\
        );

    \I__8777\ : InMux
    port map (
            O => \N__38130\,
            I => \N__38095\
        );

    \I__8776\ : Span4Mux_h
    port map (
            O => \N__38127\,
            I => \N__38092\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__38124\,
            I => \N__38089\
        );

    \I__8774\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38086\
        );

    \I__8773\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38081\
        );

    \I__8772\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38081\
        );

    \I__8771\ : Span4Mux_s2_v
    port map (
            O => \N__38118\,
            I => \N__38076\
        );

    \I__8770\ : Span4Mux_v
    port map (
            O => \N__38115\,
            I => \N__38076\
        );

    \I__8769\ : Span12Mux_v
    port map (
            O => \N__38112\,
            I => \N__38071\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38071\
        );

    \I__8767\ : InMux
    port map (
            O => \N__38108\,
            I => \N__38064\
        );

    \I__8766\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38064\
        );

    \I__8765\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38064\
        );

    \I__8764\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38061\
        );

    \I__8763\ : Span4Mux_v
    port map (
            O => \N__38100\,
            I => \N__38054\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__38095\,
            I => \N__38054\
        );

    \I__8761\ : Span4Mux_h
    port map (
            O => \N__38092\,
            I => \N__38054\
        );

    \I__8760\ : Odrv4
    port map (
            O => \N__38089\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__38086\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__38081\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8757\ : Odrv4
    port map (
            O => \N__38076\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8756\ : Odrv12
    port map (
            O => \N__38071\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__38064\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__38061\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__38054\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__38037\,
            I => \N__38024\
        );

    \I__8751\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38019\
        );

    \I__8750\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38014\
        );

    \I__8749\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38014\
        );

    \I__8748\ : CascadeMux
    port map (
            O => \N__38033\,
            I => \N__38011\
        );

    \I__8747\ : InMux
    port map (
            O => \N__38032\,
            I => \N__38008\
        );

    \I__8746\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38003\
        );

    \I__8745\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38003\
        );

    \I__8744\ : InMux
    port map (
            O => \N__38029\,
            I => \N__37994\
        );

    \I__8743\ : InMux
    port map (
            O => \N__38028\,
            I => \N__37994\
        );

    \I__8742\ : InMux
    port map (
            O => \N__38027\,
            I => \N__37994\
        );

    \I__8741\ : InMux
    port map (
            O => \N__38024\,
            I => \N__37994\
        );

    \I__8740\ : InMux
    port map (
            O => \N__38023\,
            I => \N__37991\
        );

    \I__8739\ : CascadeMux
    port map (
            O => \N__38022\,
            I => \N__37988\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__38019\,
            I => \N__37985\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__38014\,
            I => \N__37982\
        );

    \I__8736\ : InMux
    port map (
            O => \N__38011\,
            I => \N__37977\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__38008\,
            I => \N__37974\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__38003\,
            I => \N__37969\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__37994\,
            I => \N__37969\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__37991\,
            I => \N__37966\
        );

    \I__8731\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37963\
        );

    \I__8730\ : Span12Mux_s10_v
    port map (
            O => \N__37985\,
            I => \N__37958\
        );

    \I__8729\ : Span12Mux_s5_v
    port map (
            O => \N__37982\,
            I => \N__37958\
        );

    \I__8728\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37953\
        );

    \I__8727\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37953\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__37977\,
            I => \N__37942\
        );

    \I__8725\ : Span4Mux_h
    port map (
            O => \N__37974\,
            I => \N__37942\
        );

    \I__8724\ : Span4Mux_s3_v
    port map (
            O => \N__37969\,
            I => \N__37942\
        );

    \I__8723\ : Span4Mux_h
    port map (
            O => \N__37966\,
            I => \N__37942\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37942\
        );

    \I__8721\ : Odrv12
    port map (
            O => \N__37958\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__37953\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__37942\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__8718\ : CascadeMux
    port map (
            O => \N__37935\,
            I => \N__37931\
        );

    \I__8717\ : CascadeMux
    port map (
            O => \N__37934\,
            I => \N__37924\
        );

    \I__8716\ : InMux
    port map (
            O => \N__37931\,
            I => \N__37920\
        );

    \I__8715\ : InMux
    port map (
            O => \N__37930\,
            I => \N__37917\
        );

    \I__8714\ : CascadeMux
    port map (
            O => \N__37929\,
            I => \N__37912\
        );

    \I__8713\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37907\
        );

    \I__8712\ : InMux
    port map (
            O => \N__37927\,
            I => \N__37904\
        );

    \I__8711\ : InMux
    port map (
            O => \N__37924\,
            I => \N__37899\
        );

    \I__8710\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37899\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__37920\,
            I => \N__37896\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__37917\,
            I => \N__37893\
        );

    \I__8707\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37888\
        );

    \I__8706\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37888\
        );

    \I__8705\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37885\
        );

    \I__8704\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37882\
        );

    \I__8703\ : CascadeMux
    port map (
            O => \N__37910\,
            I => \N__37878\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__37907\,
            I => \N__37865\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__37904\,
            I => \N__37865\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__37899\,
            I => \N__37862\
        );

    \I__8699\ : Span4Mux_v
    port map (
            O => \N__37896\,
            I => \N__37855\
        );

    \I__8698\ : Span4Mux_v
    port map (
            O => \N__37893\,
            I => \N__37855\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__37888\,
            I => \N__37855\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37850\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__37882\,
            I => \N__37850\
        );

    \I__8694\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37843\
        );

    \I__8693\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37843\
        );

    \I__8692\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37843\
        );

    \I__8691\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37840\
        );

    \I__8690\ : CascadeMux
    port map (
            O => \N__37875\,
            I => \N__37837\
        );

    \I__8689\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37832\
        );

    \I__8688\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37832\
        );

    \I__8687\ : InMux
    port map (
            O => \N__37872\,
            I => \N__37825\
        );

    \I__8686\ : InMux
    port map (
            O => \N__37871\,
            I => \N__37825\
        );

    \I__8685\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37825\
        );

    \I__8684\ : Span4Mux_s1_v
    port map (
            O => \N__37865\,
            I => \N__37820\
        );

    \I__8683\ : Span4Mux_v
    port map (
            O => \N__37862\,
            I => \N__37820\
        );

    \I__8682\ : Span4Mux_h
    port map (
            O => \N__37855\,
            I => \N__37817\
        );

    \I__8681\ : Span4Mux_v
    port map (
            O => \N__37850\,
            I => \N__37812\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__37843\,
            I => \N__37812\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__37840\,
            I => \N__37809\
        );

    \I__8678\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37806\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__37832\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__37825\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8675\ : Odrv4
    port map (
            O => \N__37820\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__37817\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8673\ : Odrv4
    port map (
            O => \N__37812\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8672\ : Odrv12
    port map (
            O => \N__37809\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__37806\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__8670\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37788\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__37788\,
            I => \b2v_inst11.un1_i2_mux_0\
        );

    \I__8668\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37782\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__37782\,
            I => \b2v_inst11.un1_N_5\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__37779\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_\
        );

    \I__8665\ : InMux
    port map (
            O => \N__37776\,
            I => \N__37773\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__37773\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_12\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__37770\,
            I => \N__37758\
        );

    \I__8662\ : CascadeMux
    port map (
            O => \N__37769\,
            I => \N__37753\
        );

    \I__8661\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37750\
        );

    \I__8660\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37743\
        );

    \I__8659\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37740\
        );

    \I__8658\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37731\
        );

    \I__8657\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37731\
        );

    \I__8656\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37731\
        );

    \I__8655\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37731\
        );

    \I__8654\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37724\
        );

    \I__8653\ : InMux
    port map (
            O => \N__37758\,
            I => \N__37724\
        );

    \I__8652\ : InMux
    port map (
            O => \N__37757\,
            I => \N__37724\
        );

    \I__8651\ : InMux
    port map (
            O => \N__37756\,
            I => \N__37721\
        );

    \I__8650\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37718\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37715\
        );

    \I__8648\ : InMux
    port map (
            O => \N__37749\,
            I => \N__37706\
        );

    \I__8647\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37706\
        );

    \I__8646\ : InMux
    port map (
            O => \N__37747\,
            I => \N__37706\
        );

    \I__8645\ : InMux
    port map (
            O => \N__37746\,
            I => \N__37706\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__37743\,
            I => \N__37701\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__37740\,
            I => \N__37698\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__37731\,
            I => \N__37693\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__37724\,
            I => \N__37693\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37690\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__37718\,
            I => \N__37687\
        );

    \I__8638\ : Span4Mux_v
    port map (
            O => \N__37715\,
            I => \N__37682\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__37706\,
            I => \N__37682\
        );

    \I__8636\ : InMux
    port map (
            O => \N__37705\,
            I => \N__37677\
        );

    \I__8635\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37677\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__37701\,
            I => \N__37670\
        );

    \I__8633\ : Span4Mux_v
    port map (
            O => \N__37698\,
            I => \N__37670\
        );

    \I__8632\ : Span4Mux_v
    port map (
            O => \N__37693\,
            I => \N__37670\
        );

    \I__8631\ : Span4Mux_s2_v
    port map (
            O => \N__37690\,
            I => \N__37665\
        );

    \I__8630\ : Span4Mux_s2_h
    port map (
            O => \N__37687\,
            I => \N__37665\
        );

    \I__8629\ : Odrv4
    port map (
            O => \N__37682\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__37677\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__8627\ : Odrv4
    port map (
            O => \N__37670\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__8626\ : Odrv4
    port map (
            O => \N__37665\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__8625\ : CascadeMux
    port map (
            O => \N__37656\,
            I => \b2v_inst11.un1_dutycycle_53_s_9_sf_cascade_\
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__8623\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37647\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__37647\,
            I => \N__37644\
        );

    \I__8621\ : Odrv12
    port map (
            O => \N__37644\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_12\
        );

    \I__8620\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37638\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__37638\,
            I => \N__37635\
        );

    \I__8618\ : Span4Mux_h
    port map (
            O => \N__37635\,
            I => \N__37632\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__37632\,
            I => \N__37629\
        );

    \I__8616\ : Span4Mux_v
    port map (
            O => \N__37629\,
            I => \N__37626\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__37626\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_1\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__37623\,
            I => \b2v_inst11.N_371_cascade_\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__37620\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_cascade_\
        );

    \I__8612\ : InMux
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__37614\,
            I => \N__37611\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__37611\,
            I => \N__37608\
        );

    \I__8609\ : Span4Mux_v
    port map (
            O => \N__37608\,
            I => \N__37605\
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__37605\,
            I => \b2v_inst11.func_state_RNIDUQ02Z0Z_1\
        );

    \I__8607\ : InMux
    port map (
            O => \N__37602\,
            I => \N__37599\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__37599\,
            I => \b2v_inst11.g2_0_0Z0Z_0\
        );

    \I__8605\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37590\
        );

    \I__8604\ : CascadeMux
    port map (
            O => \N__37595\,
            I => \N__37585\
        );

    \I__8603\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37579\
        );

    \I__8602\ : InMux
    port map (
            O => \N__37593\,
            I => \N__37576\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__37590\,
            I => \N__37573\
        );

    \I__8600\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37570\
        );

    \I__8599\ : InMux
    port map (
            O => \N__37588\,
            I => \N__37565\
        );

    \I__8598\ : InMux
    port map (
            O => \N__37585\,
            I => \N__37565\
        );

    \I__8597\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37560\
        );

    \I__8596\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37560\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__37582\,
            I => \N__37557\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__37579\,
            I => \N__37554\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__37576\,
            I => \N__37549\
        );

    \I__8592\ : Span4Mux_s3_h
    port map (
            O => \N__37573\,
            I => \N__37549\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__37570\,
            I => \N__37544\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37544\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__37560\,
            I => \N__37541\
        );

    \I__8588\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37537\
        );

    \I__8587\ : Span4Mux_v
    port map (
            O => \N__37554\,
            I => \N__37534\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__37549\,
            I => \N__37527\
        );

    \I__8585\ : Span4Mux_s2_v
    port map (
            O => \N__37544\,
            I => \N__37527\
        );

    \I__8584\ : Span4Mux_s2_v
    port map (
            O => \N__37541\,
            I => \N__37527\
        );

    \I__8583\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37524\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__37537\,
            I => \N__37519\
        );

    \I__8581\ : Span4Mux_h
    port map (
            O => \N__37534\,
            I => \N__37519\
        );

    \I__8580\ : Odrv4
    port map (
            O => \N__37527\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__37524\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__8578\ : Odrv4
    port map (
            O => \N__37519\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__8577\ : CascadeMux
    port map (
            O => \N__37512\,
            I => \N__37503\
        );

    \I__8576\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37495\
        );

    \I__8575\ : InMux
    port map (
            O => \N__37510\,
            I => \N__37495\
        );

    \I__8574\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37492\
        );

    \I__8573\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37489\
        );

    \I__8572\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37486\
        );

    \I__8571\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37477\
        );

    \I__8570\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37477\
        );

    \I__8569\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37477\
        );

    \I__8568\ : InMux
    port map (
            O => \N__37501\,
            I => \N__37477\
        );

    \I__8567\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37474\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__37495\,
            I => \N__37471\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__37492\,
            I => \N__37468\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__37489\,
            I => \N__37465\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__37486\,
            I => \N__37462\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__37477\,
            I => \N__37459\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__37474\,
            I => \N__37454\
        );

    \I__8560\ : Span4Mux_s2_h
    port map (
            O => \N__37471\,
            I => \N__37454\
        );

    \I__8559\ : Span4Mux_v
    port map (
            O => \N__37468\,
            I => \N__37449\
        );

    \I__8558\ : Span4Mux_v
    port map (
            O => \N__37465\,
            I => \N__37449\
        );

    \I__8557\ : Span4Mux_s2_h
    port map (
            O => \N__37462\,
            I => \N__37446\
        );

    \I__8556\ : Span4Mux_s2_h
    port map (
            O => \N__37459\,
            I => \N__37441\
        );

    \I__8555\ : Span4Mux_v
    port map (
            O => \N__37454\,
            I => \N__37441\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__37449\,
            I => \b2v_inst11.N_140_N\
        );

    \I__8553\ : Odrv4
    port map (
            O => \N__37446\,
            I => \b2v_inst11.N_140_N\
        );

    \I__8552\ : Odrv4
    port map (
            O => \N__37441\,
            I => \b2v_inst11.N_140_N\
        );

    \I__8551\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37417\
        );

    \I__8550\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37417\
        );

    \I__8549\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37417\
        );

    \I__8548\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37417\
        );

    \I__8547\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37412\
        );

    \I__8546\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37412\
        );

    \I__8545\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37409\
        );

    \I__8544\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37403\
        );

    \I__8543\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37403\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__37417\,
            I => \N__37399\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__37412\,
            I => \N__37394\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__37409\,
            I => \N__37394\
        );

    \I__8539\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37391\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__37403\,
            I => \N__37388\
        );

    \I__8537\ : InMux
    port map (
            O => \N__37402\,
            I => \N__37385\
        );

    \I__8536\ : Span4Mux_s0_h
    port map (
            O => \N__37399\,
            I => \N__37380\
        );

    \I__8535\ : Span4Mux_v
    port map (
            O => \N__37394\,
            I => \N__37380\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__37391\,
            I => \N__37375\
        );

    \I__8533\ : Span4Mux_s3_h
    port map (
            O => \N__37388\,
            I => \N__37375\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__37385\,
            I => \N__37372\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__37380\,
            I => \b2v_inst11.N_425\
        );

    \I__8530\ : Odrv4
    port map (
            O => \N__37375\,
            I => \b2v_inst11.N_425\
        );

    \I__8529\ : Odrv4
    port map (
            O => \N__37372\,
            I => \b2v_inst11.N_425\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__37365\,
            I => \b2v_inst11.N_158_N_cascade_\
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__37362\,
            I => \N__37358\
        );

    \I__8526\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37351\
        );

    \I__8525\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37351\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__37357\,
            I => \N__37347\
        );

    \I__8523\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37337\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__37351\,
            I => \N__37334\
        );

    \I__8521\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37327\
        );

    \I__8520\ : InMux
    port map (
            O => \N__37347\,
            I => \N__37327\
        );

    \I__8519\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37327\
        );

    \I__8518\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37324\
        );

    \I__8517\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37320\
        );

    \I__8516\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37317\
        );

    \I__8515\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37311\
        );

    \I__8514\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37311\
        );

    \I__8513\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37308\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37305\
        );

    \I__8511\ : Span4Mux_v
    port map (
            O => \N__37334\,
            I => \N__37300\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__37327\,
            I => \N__37300\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37297\
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__37323\,
            I => \N__37294\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__37320\,
            I => \N__37284\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37284\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__37316\,
            I => \N__37279\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__37311\,
            I => \N__37272\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__37308\,
            I => \N__37272\
        );

    \I__8502\ : Span4Mux_v
    port map (
            O => \N__37305\,
            I => \N__37265\
        );

    \I__8501\ : Span4Mux_v
    port map (
            O => \N__37300\,
            I => \N__37265\
        );

    \I__8500\ : Span4Mux_h
    port map (
            O => \N__37297\,
            I => \N__37265\
        );

    \I__8499\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37262\
        );

    \I__8498\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37257\
        );

    \I__8497\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37257\
        );

    \I__8496\ : InMux
    port map (
            O => \N__37291\,
            I => \N__37254\
        );

    \I__8495\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37249\
        );

    \I__8494\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37249\
        );

    \I__8493\ : Span4Mux_h
    port map (
            O => \N__37284\,
            I => \N__37246\
        );

    \I__8492\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37241\
        );

    \I__8491\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37241\
        );

    \I__8490\ : InMux
    port map (
            O => \N__37279\,
            I => \N__37234\
        );

    \I__8489\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37234\
        );

    \I__8488\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37234\
        );

    \I__8487\ : Span4Mux_h
    port map (
            O => \N__37272\,
            I => \N__37229\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__37265\,
            I => \N__37229\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__37262\,
            I => \N__37224\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__37257\,
            I => \N__37224\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__37254\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__37249\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8481\ : Odrv4
    port map (
            O => \N__37246\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__37241\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__37234\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__37229\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8477\ : Odrv12
    port map (
            O => \N__37224\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__8476\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37206\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__37206\,
            I => \b2v_inst11.dutycycle_en_12\
        );

    \I__8474\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37197\
        );

    \I__8473\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37197\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__37197\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3AZ0Z64\
        );

    \I__8471\ : CascadeMux
    port map (
            O => \N__37194\,
            I => \b2v_inst11.dutycycle_en_12_cascade_\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__37191\,
            I => \N__37187\
        );

    \I__8469\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37182\
        );

    \I__8468\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37182\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__37182\,
            I => \b2v_inst11.dutycycleZ0Z_15\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__37179\,
            I => \N__37175\
        );

    \I__8465\ : InMux
    port map (
            O => \N__37178\,
            I => \N__37172\
        );

    \I__8464\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37169\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37165\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__37169\,
            I => \N__37162\
        );

    \I__8461\ : InMux
    port map (
            O => \N__37168\,
            I => \N__37159\
        );

    \I__8460\ : Span12Mux_s8_v
    port map (
            O => \N__37165\,
            I => \N__37154\
        );

    \I__8459\ : Span12Mux_s0_h
    port map (
            O => \N__37162\,
            I => \N__37154\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__37159\,
            I => \b2v_inst11.N_326_N\
        );

    \I__8457\ : Odrv12
    port map (
            O => \N__37154\,
            I => \b2v_inst11.N_326_N\
        );

    \I__8456\ : ClkMux
    port map (
            O => \N__37149\,
            I => \N__37145\
        );

    \I__8455\ : ClkMux
    port map (
            O => \N__37148\,
            I => \N__37136\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37131\
        );

    \I__8453\ : ClkMux
    port map (
            O => \N__37144\,
            I => \N__37128\
        );

    \I__8452\ : ClkMux
    port map (
            O => \N__37143\,
            I => \N__37122\
        );

    \I__8451\ : ClkMux
    port map (
            O => \N__37142\,
            I => \N__37119\
        );

    \I__8450\ : ClkMux
    port map (
            O => \N__37141\,
            I => \N__37116\
        );

    \I__8449\ : ClkMux
    port map (
            O => \N__37140\,
            I => \N__37113\
        );

    \I__8448\ : ClkMux
    port map (
            O => \N__37139\,
            I => \N__37110\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__37136\,
            I => \N__37105\
        );

    \I__8446\ : ClkMux
    port map (
            O => \N__37135\,
            I => \N__37102\
        );

    \I__8445\ : ClkMux
    port map (
            O => \N__37134\,
            I => \N__37096\
        );

    \I__8444\ : Span4Mux_s1_h
    port map (
            O => \N__37131\,
            I => \N__37092\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__37128\,
            I => \N__37089\
        );

    \I__8442\ : ClkMux
    port map (
            O => \N__37127\,
            I => \N__37082\
        );

    \I__8441\ : ClkMux
    port map (
            O => \N__37126\,
            I => \N__37079\
        );

    \I__8440\ : ClkMux
    port map (
            O => \N__37125\,
            I => \N__37076\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37073\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__37119\,
            I => \N__37064\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37055\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__37113\,
            I => \N__37055\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__37110\,
            I => \N__37055\
        );

    \I__8434\ : ClkMux
    port map (
            O => \N__37109\,
            I => \N__37052\
        );

    \I__8433\ : ClkMux
    port map (
            O => \N__37108\,
            I => \N__37049\
        );

    \I__8432\ : Span4Mux_v
    port map (
            O => \N__37105\,
            I => \N__37044\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__37102\,
            I => \N__37044\
        );

    \I__8430\ : ClkMux
    port map (
            O => \N__37101\,
            I => \N__37041\
        );

    \I__8429\ : ClkMux
    port map (
            O => \N__37100\,
            I => \N__37038\
        );

    \I__8428\ : ClkMux
    port map (
            O => \N__37099\,
            I => \N__37035\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__37096\,
            I => \N__37031\
        );

    \I__8426\ : ClkMux
    port map (
            O => \N__37095\,
            I => \N__37028\
        );

    \I__8425\ : Span4Mux_v
    port map (
            O => \N__37092\,
            I => \N__37022\
        );

    \I__8424\ : Span4Mux_s1_h
    port map (
            O => \N__37089\,
            I => \N__37022\
        );

    \I__8423\ : ClkMux
    port map (
            O => \N__37088\,
            I => \N__37019\
        );

    \I__8422\ : ClkMux
    port map (
            O => \N__37087\,
            I => \N__37015\
        );

    \I__8421\ : ClkMux
    port map (
            O => \N__37086\,
            I => \N__37011\
        );

    \I__8420\ : ClkMux
    port map (
            O => \N__37085\,
            I => \N__37008\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__37082\,
            I => \N__37003\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__37079\,
            I => \N__36998\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__37076\,
            I => \N__36993\
        );

    \I__8416\ : Span4Mux_v
    port map (
            O => \N__37073\,
            I => \N__36990\
        );

    \I__8415\ : ClkMux
    port map (
            O => \N__37072\,
            I => \N__36987\
        );

    \I__8414\ : ClkMux
    port map (
            O => \N__37071\,
            I => \N__36984\
        );

    \I__8413\ : ClkMux
    port map (
            O => \N__37070\,
            I => \N__36981\
        );

    \I__8412\ : ClkMux
    port map (
            O => \N__37069\,
            I => \N__36977\
        );

    \I__8411\ : ClkMux
    port map (
            O => \N__37068\,
            I => \N__36974\
        );

    \I__8410\ : ClkMux
    port map (
            O => \N__37067\,
            I => \N__36970\
        );

    \I__8409\ : Span4Mux_s2_h
    port map (
            O => \N__37064\,
            I => \N__36962\
        );

    \I__8408\ : ClkMux
    port map (
            O => \N__37063\,
            I => \N__36959\
        );

    \I__8407\ : ClkMux
    port map (
            O => \N__37062\,
            I => \N__36956\
        );

    \I__8406\ : Span4Mux_v
    port map (
            O => \N__37055\,
            I => \N__36948\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__37052\,
            I => \N__36948\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__36948\
        );

    \I__8403\ : Span4Mux_v
    port map (
            O => \N__37044\,
            I => \N__36943\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__37041\,
            I => \N__36943\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__37038\,
            I => \N__36939\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__37035\,
            I => \N__36936\
        );

    \I__8399\ : ClkMux
    port map (
            O => \N__37034\,
            I => \N__36933\
        );

    \I__8398\ : Span4Mux_v
    port map (
            O => \N__37031\,
            I => \N__36928\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__37028\,
            I => \N__36928\
        );

    \I__8396\ : ClkMux
    port map (
            O => \N__37027\,
            I => \N__36925\
        );

    \I__8395\ : Span4Mux_h
    port map (
            O => \N__37022\,
            I => \N__36922\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__37019\,
            I => \N__36919\
        );

    \I__8393\ : ClkMux
    port map (
            O => \N__37018\,
            I => \N__36916\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__37015\,
            I => \N__36913\
        );

    \I__8391\ : ClkMux
    port map (
            O => \N__37014\,
            I => \N__36910\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__37011\,
            I => \N__36906\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__37008\,
            I => \N__36903\
        );

    \I__8388\ : ClkMux
    port map (
            O => \N__37007\,
            I => \N__36900\
        );

    \I__8387\ : ClkMux
    port map (
            O => \N__37006\,
            I => \N__36895\
        );

    \I__8386\ : Span4Mux_s1_h
    port map (
            O => \N__37003\,
            I => \N__36892\
        );

    \I__8385\ : ClkMux
    port map (
            O => \N__37002\,
            I => \N__36886\
        );

    \I__8384\ : ClkMux
    port map (
            O => \N__37001\,
            I => \N__36883\
        );

    \I__8383\ : Span4Mux_v
    port map (
            O => \N__36998\,
            I => \N__36880\
        );

    \I__8382\ : ClkMux
    port map (
            O => \N__36997\,
            I => \N__36877\
        );

    \I__8381\ : ClkMux
    port map (
            O => \N__36996\,
            I => \N__36874\
        );

    \I__8380\ : Span4Mux_h
    port map (
            O => \N__36993\,
            I => \N__36863\
        );

    \I__8379\ : Span4Mux_h
    port map (
            O => \N__36990\,
            I => \N__36863\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__36987\,
            I => \N__36863\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__36984\,
            I => \N__36863\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__36981\,
            I => \N__36858\
        );

    \I__8375\ : ClkMux
    port map (
            O => \N__36980\,
            I => \N__36855\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36850\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36850\
        );

    \I__8372\ : ClkMux
    port map (
            O => \N__36973\,
            I => \N__36847\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__36970\,
            I => \N__36844\
        );

    \I__8370\ : ClkMux
    port map (
            O => \N__36969\,
            I => \N__36841\
        );

    \I__8369\ : ClkMux
    port map (
            O => \N__36968\,
            I => \N__36837\
        );

    \I__8368\ : ClkMux
    port map (
            O => \N__36967\,
            I => \N__36831\
        );

    \I__8367\ : ClkMux
    port map (
            O => \N__36966\,
            I => \N__36827\
        );

    \I__8366\ : ClkMux
    port map (
            O => \N__36965\,
            I => \N__36824\
        );

    \I__8365\ : Span4Mux_h
    port map (
            O => \N__36962\,
            I => \N__36817\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__36959\,
            I => \N__36817\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__36956\,
            I => \N__36814\
        );

    \I__8362\ : ClkMux
    port map (
            O => \N__36955\,
            I => \N__36811\
        );

    \I__8361\ : Span4Mux_v
    port map (
            O => \N__36948\,
            I => \N__36805\
        );

    \I__8360\ : Span4Mux_v
    port map (
            O => \N__36943\,
            I => \N__36805\
        );

    \I__8359\ : ClkMux
    port map (
            O => \N__36942\,
            I => \N__36802\
        );

    \I__8358\ : Span4Mux_s1_h
    port map (
            O => \N__36939\,
            I => \N__36793\
        );

    \I__8357\ : Span4Mux_v
    port map (
            O => \N__36936\,
            I => \N__36793\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__36933\,
            I => \N__36793\
        );

    \I__8355\ : Span4Mux_v
    port map (
            O => \N__36928\,
            I => \N__36788\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__36925\,
            I => \N__36788\
        );

    \I__8353\ : Span4Mux_v
    port map (
            O => \N__36922\,
            I => \N__36781\
        );

    \I__8352\ : Span4Mux_v
    port map (
            O => \N__36919\,
            I => \N__36781\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__36916\,
            I => \N__36781\
        );

    \I__8350\ : Span4Mux_v
    port map (
            O => \N__36913\,
            I => \N__36776\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__36910\,
            I => \N__36776\
        );

    \I__8348\ : ClkMux
    port map (
            O => \N__36909\,
            I => \N__36771\
        );

    \I__8347\ : Span4Mux_s1_h
    port map (
            O => \N__36906\,
            I => \N__36768\
        );

    \I__8346\ : Span4Mux_s1_h
    port map (
            O => \N__36903\,
            I => \N__36765\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__36900\,
            I => \N__36762\
        );

    \I__8344\ : ClkMux
    port map (
            O => \N__36899\,
            I => \N__36759\
        );

    \I__8343\ : ClkMux
    port map (
            O => \N__36898\,
            I => \N__36756\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__36895\,
            I => \N__36752\
        );

    \I__8341\ : Span4Mux_h
    port map (
            O => \N__36892\,
            I => \N__36749\
        );

    \I__8340\ : ClkMux
    port map (
            O => \N__36891\,
            I => \N__36746\
        );

    \I__8339\ : ClkMux
    port map (
            O => \N__36890\,
            I => \N__36741\
        );

    \I__8338\ : ClkMux
    port map (
            O => \N__36889\,
            I => \N__36738\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__36886\,
            I => \N__36733\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__36883\,
            I => \N__36733\
        );

    \I__8335\ : Span4Mux_h
    port map (
            O => \N__36880\,
            I => \N__36726\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__36877\,
            I => \N__36726\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__36874\,
            I => \N__36726\
        );

    \I__8332\ : ClkMux
    port map (
            O => \N__36873\,
            I => \N__36723\
        );

    \I__8331\ : ClkMux
    port map (
            O => \N__36872\,
            I => \N__36720\
        );

    \I__8330\ : Span4Mux_v
    port map (
            O => \N__36863\,
            I => \N__36716\
        );

    \I__8329\ : ClkMux
    port map (
            O => \N__36862\,
            I => \N__36713\
        );

    \I__8328\ : ClkMux
    port map (
            O => \N__36861\,
            I => \N__36710\
        );

    \I__8327\ : Span4Mux_s3_h
    port map (
            O => \N__36858\,
            I => \N__36704\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__36855\,
            I => \N__36704\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__36850\,
            I => \N__36695\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__36847\,
            I => \N__36695\
        );

    \I__8323\ : Span4Mux_s3_h
    port map (
            O => \N__36844\,
            I => \N__36695\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__36841\,
            I => \N__36695\
        );

    \I__8321\ : ClkMux
    port map (
            O => \N__36840\,
            I => \N__36692\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__36837\,
            I => \N__36689\
        );

    \I__8319\ : ClkMux
    port map (
            O => \N__36836\,
            I => \N__36686\
        );

    \I__8318\ : ClkMux
    port map (
            O => \N__36835\,
            I => \N__36683\
        );

    \I__8317\ : ClkMux
    port map (
            O => \N__36834\,
            I => \N__36680\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__36831\,
            I => \N__36677\
        );

    \I__8315\ : ClkMux
    port map (
            O => \N__36830\,
            I => \N__36674\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__36827\,
            I => \N__36668\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__36824\,
            I => \N__36668\
        );

    \I__8312\ : ClkMux
    port map (
            O => \N__36823\,
            I => \N__36665\
        );

    \I__8311\ : ClkMux
    port map (
            O => \N__36822\,
            I => \N__36662\
        );

    \I__8310\ : Span4Mux_v
    port map (
            O => \N__36817\,
            I => \N__36655\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__36814\,
            I => \N__36655\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__36811\,
            I => \N__36655\
        );

    \I__8307\ : ClkMux
    port map (
            O => \N__36810\,
            I => \N__36652\
        );

    \I__8306\ : IoSpan4Mux
    port map (
            O => \N__36805\,
            I => \N__36647\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__36802\,
            I => \N__36647\
        );

    \I__8304\ : ClkMux
    port map (
            O => \N__36801\,
            I => \N__36644\
        );

    \I__8303\ : ClkMux
    port map (
            O => \N__36800\,
            I => \N__36641\
        );

    \I__8302\ : Span4Mux_v
    port map (
            O => \N__36793\,
            I => \N__36636\
        );

    \I__8301\ : Span4Mux_v
    port map (
            O => \N__36788\,
            I => \N__36633\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__36781\,
            I => \N__36628\
        );

    \I__8299\ : Span4Mux_h
    port map (
            O => \N__36776\,
            I => \N__36628\
        );

    \I__8298\ : ClkMux
    port map (
            O => \N__36775\,
            I => \N__36625\
        );

    \I__8297\ : ClkMux
    port map (
            O => \N__36774\,
            I => \N__36622\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__36771\,
            I => \N__36619\
        );

    \I__8295\ : Span4Mux_h
    port map (
            O => \N__36768\,
            I => \N__36612\
        );

    \I__8294\ : Span4Mux_h
    port map (
            O => \N__36765\,
            I => \N__36612\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__36762\,
            I => \N__36612\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__36759\,
            I => \N__36608\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__36756\,
            I => \N__36605\
        );

    \I__8290\ : ClkMux
    port map (
            O => \N__36755\,
            I => \N__36602\
        );

    \I__8289\ : Span4Mux_s1_h
    port map (
            O => \N__36752\,
            I => \N__36599\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__36749\,
            I => \N__36594\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36594\
        );

    \I__8286\ : ClkMux
    port map (
            O => \N__36745\,
            I => \N__36591\
        );

    \I__8285\ : ClkMux
    port map (
            O => \N__36744\,
            I => \N__36588\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__36741\,
            I => \N__36585\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__36738\,
            I => \N__36582\
        );

    \I__8282\ : Span4Mux_v
    port map (
            O => \N__36733\,
            I => \N__36573\
        );

    \I__8281\ : Span4Mux_v
    port map (
            O => \N__36726\,
            I => \N__36573\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__36723\,
            I => \N__36573\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__36720\,
            I => \N__36573\
        );

    \I__8278\ : ClkMux
    port map (
            O => \N__36719\,
            I => \N__36570\
        );

    \I__8277\ : Span4Mux_h
    port map (
            O => \N__36716\,
            I => \N__36565\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__36713\,
            I => \N__36565\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__36710\,
            I => \N__36562\
        );

    \I__8274\ : ClkMux
    port map (
            O => \N__36709\,
            I => \N__36559\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__36704\,
            I => \N__36544\
        );

    \I__8272\ : Span4Mux_v
    port map (
            O => \N__36695\,
            I => \N__36544\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__36692\,
            I => \N__36544\
        );

    \I__8270\ : Span4Mux_s3_h
    port map (
            O => \N__36689\,
            I => \N__36544\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__36686\,
            I => \N__36544\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__36683\,
            I => \N__36544\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__36680\,
            I => \N__36544\
        );

    \I__8266\ : Span4Mux_s2_h
    port map (
            O => \N__36677\,
            I => \N__36541\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36538\
        );

    \I__8264\ : ClkMux
    port map (
            O => \N__36673\,
            I => \N__36535\
        );

    \I__8263\ : Span4Mux_h
    port map (
            O => \N__36668\,
            I => \N__36528\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__36665\,
            I => \N__36528\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__36662\,
            I => \N__36528\
        );

    \I__8260\ : Span4Mux_v
    port map (
            O => \N__36655\,
            I => \N__36523\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__36652\,
            I => \N__36523\
        );

    \I__8258\ : Span4Mux_s0_v
    port map (
            O => \N__36647\,
            I => \N__36516\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__36644\,
            I => \N__36516\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__36641\,
            I => \N__36516\
        );

    \I__8255\ : ClkMux
    port map (
            O => \N__36640\,
            I => \N__36513\
        );

    \I__8254\ : ClkMux
    port map (
            O => \N__36639\,
            I => \N__36509\
        );

    \I__8253\ : Span4Mux_h
    port map (
            O => \N__36636\,
            I => \N__36498\
        );

    \I__8252\ : Span4Mux_h
    port map (
            O => \N__36633\,
            I => \N__36498\
        );

    \I__8251\ : Span4Mux_h
    port map (
            O => \N__36628\,
            I => \N__36498\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__36625\,
            I => \N__36498\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__36622\,
            I => \N__36498\
        );

    \I__8248\ : Span4Mux_v
    port map (
            O => \N__36619\,
            I => \N__36493\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__36612\,
            I => \N__36493\
        );

    \I__8246\ : ClkMux
    port map (
            O => \N__36611\,
            I => \N__36490\
        );

    \I__8245\ : Span4Mux_s1_h
    port map (
            O => \N__36608\,
            I => \N__36487\
        );

    \I__8244\ : Span4Mux_s2_h
    port map (
            O => \N__36605\,
            I => \N__36482\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__36602\,
            I => \N__36482\
        );

    \I__8242\ : Span4Mux_h
    port map (
            O => \N__36599\,
            I => \N__36473\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__36594\,
            I => \N__36473\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__36591\,
            I => \N__36473\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__36588\,
            I => \N__36473\
        );

    \I__8238\ : IoSpan4Mux
    port map (
            O => \N__36585\,
            I => \N__36470\
        );

    \I__8237\ : Span4Mux_h
    port map (
            O => \N__36582\,
            I => \N__36463\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__36573\,
            I => \N__36463\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__36570\,
            I => \N__36463\
        );

    \I__8234\ : Span4Mux_v
    port map (
            O => \N__36565\,
            I => \N__36454\
        );

    \I__8233\ : Span4Mux_s3_h
    port map (
            O => \N__36562\,
            I => \N__36454\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__36559\,
            I => \N__36454\
        );

    \I__8231\ : Span4Mux_v
    port map (
            O => \N__36544\,
            I => \N__36454\
        );

    \I__8230\ : Span4Mux_v
    port map (
            O => \N__36541\,
            I => \N__36447\
        );

    \I__8229\ : Span4Mux_s2_h
    port map (
            O => \N__36538\,
            I => \N__36447\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__36535\,
            I => \N__36447\
        );

    \I__8227\ : Span4Mux_v
    port map (
            O => \N__36528\,
            I => \N__36438\
        );

    \I__8226\ : Span4Mux_v
    port map (
            O => \N__36523\,
            I => \N__36438\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__36516\,
            I => \N__36438\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__36513\,
            I => \N__36438\
        );

    \I__8223\ : ClkMux
    port map (
            O => \N__36512\,
            I => \N__36433\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36428\
        );

    \I__8221\ : Span4Mux_s2_v
    port map (
            O => \N__36498\,
            I => \N__36428\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__36493\,
            I => \N__36424\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__36490\,
            I => \N__36421\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__36487\,
            I => \N__36414\
        );

    \I__8217\ : Span4Mux_h
    port map (
            O => \N__36482\,
            I => \N__36414\
        );

    \I__8216\ : Span4Mux_v
    port map (
            O => \N__36473\,
            I => \N__36414\
        );

    \I__8215\ : IoSpan4Mux
    port map (
            O => \N__36470\,
            I => \N__36407\
        );

    \I__8214\ : IoSpan4Mux
    port map (
            O => \N__36463\,
            I => \N__36407\
        );

    \I__8213\ : IoSpan4Mux
    port map (
            O => \N__36454\,
            I => \N__36407\
        );

    \I__8212\ : IoSpan4Mux
    port map (
            O => \N__36447\,
            I => \N__36402\
        );

    \I__8211\ : IoSpan4Mux
    port map (
            O => \N__36438\,
            I => \N__36402\
        );

    \I__8210\ : ClkMux
    port map (
            O => \N__36437\,
            I => \N__36399\
        );

    \I__8209\ : ClkMux
    port map (
            O => \N__36436\,
            I => \N__36396\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__36433\,
            I => \N__36391\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__36428\,
            I => \N__36391\
        );

    \I__8206\ : ClkMux
    port map (
            O => \N__36427\,
            I => \N__36388\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__36424\,
            I => fpga_osc
        );

    \I__8204\ : Odrv12
    port map (
            O => \N__36421\,
            I => fpga_osc
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__36414\,
            I => fpga_osc
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__36407\,
            I => fpga_osc
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__36402\,
            I => fpga_osc
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__36399\,
            I => fpga_osc
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__36396\,
            I => fpga_osc
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__36391\,
            I => fpga_osc
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__36388\,
            I => fpga_osc
        );

    \I__8196\ : SRMux
    port map (
            O => \N__36369\,
            I => \N__36363\
        );

    \I__8195\ : SRMux
    port map (
            O => \N__36368\,
            I => \N__36358\
        );

    \I__8194\ : SRMux
    port map (
            O => \N__36367\,
            I => \N__36355\
        );

    \I__8193\ : SRMux
    port map (
            O => \N__36366\,
            I => \N__36352\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__36363\,
            I => \N__36349\
        );

    \I__8191\ : SRMux
    port map (
            O => \N__36362\,
            I => \N__36345\
        );

    \I__8190\ : SRMux
    port map (
            O => \N__36361\,
            I => \N__36342\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__36358\,
            I => \N__36338\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__36355\,
            I => \N__36333\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__36352\,
            I => \N__36333\
        );

    \I__8186\ : Span4Mux_s0_h
    port map (
            O => \N__36349\,
            I => \N__36330\
        );

    \I__8185\ : SRMux
    port map (
            O => \N__36348\,
            I => \N__36327\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__36345\,
            I => \N__36321\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__36342\,
            I => \N__36318\
        );

    \I__8182\ : SRMux
    port map (
            O => \N__36341\,
            I => \N__36315\
        );

    \I__8181\ : Span4Mux_v
    port map (
            O => \N__36338\,
            I => \N__36310\
        );

    \I__8180\ : Span4Mux_v
    port map (
            O => \N__36333\,
            I => \N__36310\
        );

    \I__8179\ : Span4Mux_s2_v
    port map (
            O => \N__36330\,
            I => \N__36305\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__36327\,
            I => \N__36305\
        );

    \I__8177\ : SRMux
    port map (
            O => \N__36326\,
            I => \N__36302\
        );

    \I__8176\ : SRMux
    port map (
            O => \N__36325\,
            I => \N__36299\
        );

    \I__8175\ : SRMux
    port map (
            O => \N__36324\,
            I => \N__36296\
        );

    \I__8174\ : Span4Mux_s3_h
    port map (
            O => \N__36321\,
            I => \N__36291\
        );

    \I__8173\ : Span4Mux_s3_h
    port map (
            O => \N__36318\,
            I => \N__36291\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36288\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__36310\,
            I => \N__36285\
        );

    \I__8170\ : Span4Mux_v
    port map (
            O => \N__36305\,
            I => \N__36282\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__36302\,
            I => \N__36279\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__36299\,
            I => \N__36274\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__36296\,
            I => \N__36274\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__36291\,
            I => \N__36271\
        );

    \I__8165\ : Span4Mux_v
    port map (
            O => \N__36288\,
            I => \N__36266\
        );

    \I__8164\ : Span4Mux_h
    port map (
            O => \N__36285\,
            I => \N__36266\
        );

    \I__8163\ : Span4Mux_v
    port map (
            O => \N__36282\,
            I => \N__36263\
        );

    \I__8162\ : Span4Mux_v
    port map (
            O => \N__36279\,
            I => \N__36256\
        );

    \I__8161\ : Span4Mux_v
    port map (
            O => \N__36274\,
            I => \N__36256\
        );

    \I__8160\ : Span4Mux_s3_h
    port map (
            O => \N__36271\,
            I => \N__36256\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__36266\,
            I => \N__36253\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__36263\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__36256\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__36253\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__8155\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36243\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__36243\,
            I => \N__36240\
        );

    \I__8153\ : Span4Mux_s1_h
    port map (
            O => \N__36240\,
            I => \N__36237\
        );

    \I__8152\ : Span4Mux_v
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__36234\,
            I => \b2v_inst11.un1_dutycycle_94_s1_8\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__36231\,
            I => \N__36217\
        );

    \I__8149\ : CascadeMux
    port map (
            O => \N__36230\,
            I => \N__36212\
        );

    \I__8148\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36200\
        );

    \I__8147\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36191\
        );

    \I__8146\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36191\
        );

    \I__8145\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36191\
        );

    \I__8144\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36191\
        );

    \I__8143\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36188\
        );

    \I__8142\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36185\
        );

    \I__8141\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36182\
        );

    \I__8140\ : CascadeMux
    port map (
            O => \N__36221\,
            I => \N__36179\
        );

    \I__8139\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36170\
        );

    \I__8138\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36163\
        );

    \I__8137\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36163\
        );

    \I__8136\ : InMux
    port map (
            O => \N__36215\,
            I => \N__36163\
        );

    \I__8135\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36158\
        );

    \I__8134\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36158\
        );

    \I__8133\ : InMux
    port map (
            O => \N__36210\,
            I => \N__36151\
        );

    \I__8132\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36151\
        );

    \I__8131\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36151\
        );

    \I__8130\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36140\
        );

    \I__8129\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36140\
        );

    \I__8128\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36140\
        );

    \I__8127\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36140\
        );

    \I__8126\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36140\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__36200\,
            I => \N__36129\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__36191\,
            I => \N__36129\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36129\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__36185\,
            I => \N__36129\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__36182\,
            I => \N__36129\
        );

    \I__8120\ : InMux
    port map (
            O => \N__36179\,
            I => \N__36126\
        );

    \I__8119\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36117\
        );

    \I__8118\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36117\
        );

    \I__8117\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36117\
        );

    \I__8116\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36117\
        );

    \I__8115\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36114\
        );

    \I__8114\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36111\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__36170\,
            I => \N__36096\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36096\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__36158\,
            I => \N__36096\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__36151\,
            I => \N__36096\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__36140\,
            I => \N__36096\
        );

    \I__8108\ : Span4Mux_v
    port map (
            O => \N__36129\,
            I => \N__36096\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__36126\,
            I => \N__36096\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__36117\,
            I => \N__36091\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__36114\,
            I => \N__36091\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__36111\,
            I => \N__36088\
        );

    \I__8103\ : Span4Mux_v
    port map (
            O => \N__36096\,
            I => \N__36085\
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__36091\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__8101\ : Odrv12
    port map (
            O => \N__36088\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__8100\ : Odrv4
    port map (
            O => \N__36085\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__36078\,
            I => \N__36075\
        );

    \I__8098\ : InMux
    port map (
            O => \N__36075\,
            I => \N__36072\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__36072\,
            I => \b2v_inst11.un1_dutycycle_94_s0_8\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__36069\,
            I => \N__36065\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__36068\,
            I => \N__36062\
        );

    \I__8094\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36054\
        );

    \I__8093\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36051\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__36061\,
            I => \N__36046\
        );

    \I__8091\ : CascadeMux
    port map (
            O => \N__36060\,
            I => \N__36043\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__36059\,
            I => \N__36038\
        );

    \I__8089\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36032\
        );

    \I__8088\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36032\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__36054\,
            I => \N__36027\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__36051\,
            I => \N__36027\
        );

    \I__8085\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36024\
        );

    \I__8084\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36021\
        );

    \I__8083\ : InMux
    port map (
            O => \N__36046\,
            I => \N__36016\
        );

    \I__8082\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36013\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__36042\,
            I => \N__36006\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__36041\,
            I => \N__36001\
        );

    \I__8079\ : InMux
    port map (
            O => \N__36038\,
            I => \N__35998\
        );

    \I__8078\ : InMux
    port map (
            O => \N__36037\,
            I => \N__35995\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__36032\,
            I => \N__35992\
        );

    \I__8076\ : Span4Mux_s3_v
    port map (
            O => \N__36027\,
            I => \N__35985\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__36024\,
            I => \N__35985\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__35985\
        );

    \I__8073\ : InMux
    port map (
            O => \N__36020\,
            I => \N__35980\
        );

    \I__8072\ : InMux
    port map (
            O => \N__36019\,
            I => \N__35980\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__36016\,
            I => \N__35975\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__36013\,
            I => \N__35975\
        );

    \I__8069\ : InMux
    port map (
            O => \N__36012\,
            I => \N__35970\
        );

    \I__8068\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35970\
        );

    \I__8067\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35967\
        );

    \I__8066\ : InMux
    port map (
            O => \N__36009\,
            I => \N__35964\
        );

    \I__8065\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35959\
        );

    \I__8064\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35959\
        );

    \I__8063\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35956\
        );

    \I__8062\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35953\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__35998\,
            I => \N__35948\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__35995\,
            I => \N__35948\
        );

    \I__8059\ : Span4Mux_v
    port map (
            O => \N__35992\,
            I => \N__35941\
        );

    \I__8058\ : Span4Mux_v
    port map (
            O => \N__35985\,
            I => \N__35941\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__35980\,
            I => \N__35932\
        );

    \I__8056\ : Span4Mux_s3_v
    port map (
            O => \N__35975\,
            I => \N__35932\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__35970\,
            I => \N__35932\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__35967\,
            I => \N__35932\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__35964\,
            I => \N__35921\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__35959\,
            I => \N__35921\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__35956\,
            I => \N__35921\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__35953\,
            I => \N__35921\
        );

    \I__8049\ : Span4Mux_s3_v
    port map (
            O => \N__35948\,
            I => \N__35921\
        );

    \I__8048\ : InMux
    port map (
            O => \N__35947\,
            I => \N__35914\
        );

    \I__8047\ : InMux
    port map (
            O => \N__35946\,
            I => \N__35914\
        );

    \I__8046\ : Span4Mux_s0_h
    port map (
            O => \N__35941\,
            I => \N__35907\
        );

    \I__8045\ : Span4Mux_v
    port map (
            O => \N__35932\,
            I => \N__35907\
        );

    \I__8044\ : Span4Mux_v
    port map (
            O => \N__35921\,
            I => \N__35907\
        );

    \I__8043\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35902\
        );

    \I__8042\ : InMux
    port map (
            O => \N__35919\,
            I => \N__35902\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__35914\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__8040\ : Odrv4
    port map (
            O => \N__35907\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__35902\,
            I => \b2v_inst11.dutycycleZ1Z_5\
        );

    \I__8038\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35892\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__35892\,
            I => \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1\
        );

    \I__8036\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35883\
        );

    \I__8035\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35883\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__35883\,
            I => \b2v_inst11.dutycycleZ1Z_8\
        );

    \I__8033\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35874\
        );

    \I__8032\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35874\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__35874\,
            I => \N__35871\
        );

    \I__8030\ : Odrv12
    port map (
            O => \N__35871\,
            I => \b2v_inst11.dutycycle_eena_3\
        );

    \I__8029\ : CascadeMux
    port map (
            O => \N__35868\,
            I => \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1_cascade_\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__35865\,
            I => \N__35861\
        );

    \I__8027\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35853\
        );

    \I__8026\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35849\
        );

    \I__8025\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35846\
        );

    \I__8024\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35838\
        );

    \I__8023\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35838\
        );

    \I__8022\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35838\
        );

    \I__8021\ : CascadeMux
    port map (
            O => \N__35856\,
            I => \N__35824\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__35853\,
            I => \N__35821\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__35852\,
            I => \N__35818\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__35849\,
            I => \N__35812\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__35846\,
            I => \N__35812\
        );

    \I__8016\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35809\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__35838\,
            I => \N__35805\
        );

    \I__8014\ : InMux
    port map (
            O => \N__35837\,
            I => \N__35800\
        );

    \I__8013\ : InMux
    port map (
            O => \N__35836\,
            I => \N__35800\
        );

    \I__8012\ : InMux
    port map (
            O => \N__35835\,
            I => \N__35793\
        );

    \I__8011\ : InMux
    port map (
            O => \N__35834\,
            I => \N__35793\
        );

    \I__8010\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35783\
        );

    \I__8009\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35783\
        );

    \I__8008\ : CascadeMux
    port map (
            O => \N__35831\,
            I => \N__35776\
        );

    \I__8007\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35771\
        );

    \I__8006\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35771\
        );

    \I__8005\ : IoInMux
    port map (
            O => \N__35828\,
            I => \N__35768\
        );

    \I__8004\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35765\
        );

    \I__8003\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35762\
        );

    \I__8002\ : Span4Mux_s1_h
    port map (
            O => \N__35821\,
            I => \N__35759\
        );

    \I__8001\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35754\
        );

    \I__8000\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35754\
        );

    \I__7999\ : Span4Mux_s1_h
    port map (
            O => \N__35812\,
            I => \N__35751\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35748\
        );

    \I__7997\ : InMux
    port map (
            O => \N__35808\,
            I => \N__35745\
        );

    \I__7996\ : Span4Mux_s2_h
    port map (
            O => \N__35805\,
            I => \N__35742\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35739\
        );

    \I__7994\ : InMux
    port map (
            O => \N__35799\,
            I => \N__35736\
        );

    \I__7993\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35733\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__35793\,
            I => \N__35730\
        );

    \I__7991\ : InMux
    port map (
            O => \N__35792\,
            I => \N__35723\
        );

    \I__7990\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35723\
        );

    \I__7989\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35723\
        );

    \I__7988\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35720\
        );

    \I__7987\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35717\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__35783\,
            I => \N__35714\
        );

    \I__7985\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35711\
        );

    \I__7984\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35708\
        );

    \I__7983\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35701\
        );

    \I__7982\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35701\
        );

    \I__7981\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35701\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35698\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__35768\,
            I => \N__35695\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35692\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__35762\,
            I => \N__35681\
        );

    \I__7976\ : Span4Mux_v
    port map (
            O => \N__35759\,
            I => \N__35681\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__35754\,
            I => \N__35681\
        );

    \I__7974\ : Span4Mux_v
    port map (
            O => \N__35751\,
            I => \N__35681\
        );

    \I__7973\ : Span4Mux_s1_h
    port map (
            O => \N__35748\,
            I => \N__35681\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__35745\,
            I => \N__35678\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__35742\,
            I => \N__35675\
        );

    \I__7970\ : Span4Mux_s2_h
    port map (
            O => \N__35739\,
            I => \N__35670\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__35736\,
            I => \N__35670\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__35733\,
            I => \N__35661\
        );

    \I__7967\ : Span4Mux_s2_h
    port map (
            O => \N__35730\,
            I => \N__35661\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__35723\,
            I => \N__35661\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35661\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35658\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__35714\,
            I => \N__35653\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__35711\,
            I => \N__35653\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__35708\,
            I => \N__35646\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35646\
        );

    \I__7959\ : Span4Mux_s2_h
    port map (
            O => \N__35698\,
            I => \N__35646\
        );

    \I__7958\ : Span4Mux_s3_v
    port map (
            O => \N__35695\,
            I => \N__35643\
        );

    \I__7957\ : Span4Mux_v
    port map (
            O => \N__35692\,
            I => \N__35638\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__35681\,
            I => \N__35638\
        );

    \I__7955\ : Span12Mux_s5_h
    port map (
            O => \N__35678\,
            I => \N__35633\
        );

    \I__7954\ : Sp12to4
    port map (
            O => \N__35675\,
            I => \N__35633\
        );

    \I__7953\ : Span4Mux_h
    port map (
            O => \N__35670\,
            I => \N__35628\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__35661\,
            I => \N__35628\
        );

    \I__7951\ : Span4Mux_s2_h
    port map (
            O => \N__35658\,
            I => \N__35621\
        );

    \I__7950\ : Span4Mux_v
    port map (
            O => \N__35653\,
            I => \N__35621\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__35646\,
            I => \N__35621\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__35643\,
            I => \G_149\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__35638\,
            I => \G_149\
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__35633\,
            I => \G_149\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__35628\,
            I => \G_149\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__35621\,
            I => \G_149\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__35610\,
            I => \b2v_inst11.dutycycleZ0Z_4_cascade_\
        );

    \I__7942\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35604\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35601\
        );

    \I__7940\ : Span4Mux_s1_h
    port map (
            O => \N__35601\,
            I => \N__35598\
        );

    \I__7939\ : Odrv4
    port map (
            O => \N__35598\,
            I => \b2v_inst11.un1_dutycycle_94_s1_10\
        );

    \I__7938\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35592\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__35592\,
            I => \b2v_inst11.un1_dutycycle_94_s0_10\
        );

    \I__7936\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35586\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__35586\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__35583\,
            I => \N__35580\
        );

    \I__7933\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35574\
        );

    \I__7932\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35574\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__35574\,
            I => \b2v_inst11.dutycycleZ1Z_10\
        );

    \I__7930\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35565\
        );

    \I__7929\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35565\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__35565\,
            I => \N__35562\
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__35562\,
            I => \b2v_inst11.dutycycle_eena_4\
        );

    \I__7926\ : CascadeMux
    port map (
            O => \N__35559\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642_cascade_\
        );

    \I__7925\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35549\
        );

    \I__7924\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35549\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__35554\,
            I => \N__35546\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__35549\,
            I => \N__35541\
        );

    \I__7921\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35538\
        );

    \I__7920\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35531\
        );

    \I__7919\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35531\
        );

    \I__7918\ : Span4Mux_s1_v
    port map (
            O => \N__35541\,
            I => \N__35527\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__35538\,
            I => \N__35524\
        );

    \I__7916\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35519\
        );

    \I__7915\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35519\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35516\
        );

    \I__7913\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35513\
        );

    \I__7912\ : Span4Mux_v
    port map (
            O => \N__35527\,
            I => \N__35510\
        );

    \I__7911\ : Span4Mux_h
    port map (
            O => \N__35524\,
            I => \N__35507\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__35519\,
            I => \N__35502\
        );

    \I__7909\ : Span4Mux_h
    port map (
            O => \N__35516\,
            I => \N__35502\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__35513\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__7907\ : Odrv4
    port map (
            O => \N__35510\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__7906\ : Odrv4
    port map (
            O => \N__35507\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__35502\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__35493\,
            I => \b2v_inst11.dutycycleZ0Z_3_cascade_\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__35490\,
            I => \N__35487\
        );

    \I__7902\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35481\
        );

    \I__7901\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35481\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__35481\,
            I => \N__35478\
        );

    \I__7899\ : Span4Mux_s3_v
    port map (
            O => \N__35478\,
            I => \N__35475\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__35475\,
            I => \b2v_inst11.un1_dutycycle_53_44_0_1\
        );

    \I__7897\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35469\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35458\
        );

    \I__7895\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35455\
        );

    \I__7894\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35450\
        );

    \I__7893\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35450\
        );

    \I__7892\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35445\
        );

    \I__7891\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35445\
        );

    \I__7890\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35442\
        );

    \I__7889\ : CascadeMux
    port map (
            O => \N__35462\,
            I => \N__35439\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__35461\,
            I => \N__35436\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__35458\,
            I => \N__35429\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__35455\,
            I => \N__35429\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__35450\,
            I => \N__35424\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__35445\,
            I => \N__35424\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__35442\,
            I => \N__35419\
        );

    \I__7882\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35416\
        );

    \I__7881\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35413\
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__35435\,
            I => \N__35410\
        );

    \I__7879\ : InMux
    port map (
            O => \N__35434\,
            I => \N__35407\
        );

    \I__7878\ : Span4Mux_s3_v
    port map (
            O => \N__35429\,
            I => \N__35404\
        );

    \I__7877\ : Span4Mux_s3_v
    port map (
            O => \N__35424\,
            I => \N__35401\
        );

    \I__7876\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35398\
        );

    \I__7875\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35395\
        );

    \I__7874\ : Span4Mux_s3_v
    port map (
            O => \N__35419\,
            I => \N__35388\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35388\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__35413\,
            I => \N__35388\
        );

    \I__7871\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35385\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__35407\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__35404\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__35401\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__35398\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__35395\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__35388\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__35385\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__7863\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35367\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__35367\,
            I => \N__35364\
        );

    \I__7861\ : Odrv4
    port map (
            O => \N__35364\,
            I => \b2v_inst11.g1_i_0\
        );

    \I__7860\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35358\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35355\
        );

    \I__7858\ : Span4Mux_v
    port map (
            O => \N__35355\,
            I => \N__35352\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__35352\,
            I => \b2v_inst11.dutycycle_eena_2\
        );

    \I__7856\ : InMux
    port map (
            O => \N__35349\,
            I => \N__35346\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__35346\,
            I => \N__35342\
        );

    \I__7854\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35339\
        );

    \I__7853\ : Span4Mux_v
    port map (
            O => \N__35342\,
            I => \N__35336\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__35339\,
            I => \N__35331\
        );

    \I__7851\ : Span4Mux_s0_h
    port map (
            O => \N__35336\,
            I => \N__35331\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__35331\,
            I => \b2v_inst11.dutycycleZ1Z_9\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__35328\,
            I => \b2v_inst11.dutycycle_eena_2_cascade_\
        );

    \I__7848\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35322\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__35322\,
            I => \N__35319\
        );

    \I__7846\ : Span4Mux_h
    port map (
            O => \N__35319\,
            I => \N__35315\
        );

    \I__7845\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35312\
        );

    \I__7844\ : Span4Mux_v
    port map (
            O => \N__35315\,
            I => \N__35309\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__35312\,
            I => \N__35306\
        );

    \I__7842\ : Odrv4
    port map (
            O => \N__35309\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1\
        );

    \I__7841\ : Odrv4
    port map (
            O => \N__35306\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__35301\,
            I => \b2v_inst11.dutycycleZ0Z_0_cascade_\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__35298\,
            I => \N__35295\
        );

    \I__7838\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35292\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__35292\,
            I => \b2v_inst11.un1_clk_100khz_30_and_i_0_0_1\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__35289\,
            I => \N__35286\
        );

    \I__7835\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35283\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__35283\,
            I => \b2v_inst11.un1_dutycycle_94_s0_5\
        );

    \I__7833\ : InMux
    port map (
            O => \N__35280\,
            I => \N__35277\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__35277\,
            I => \N__35274\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__35274\,
            I => \b2v_inst11.un1_dutycycle_94_s1_5\
        );

    \I__7830\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35268\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__35268\,
            I => \N__35265\
        );

    \I__7828\ : Odrv12
    port map (
            O => \N__35265\,
            I => \b2v_inst11.N_302\
        );

    \I__7827\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35259\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__35259\,
            I => \N__35256\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__35256\,
            I => \N__35253\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__35253\,
            I => \b2v_inst11.un1_dutycycle_94_s1_6\
        );

    \I__7823\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__35247\,
            I => \b2v_inst11.un1_dutycycle_94_s0_6\
        );

    \I__7821\ : InMux
    port map (
            O => \N__35244\,
            I => \N__35241\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__35241\,
            I => \N__35238\
        );

    \I__7819\ : Span4Mux_s0_h
    port map (
            O => \N__35238\,
            I => \N__35235\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__35235\,
            I => \b2v_inst11.N_301\
        );

    \I__7817\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35229\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__35229\,
            I => \N__35226\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__35226\,
            I => \b2v_inst11.un1_dutycycle_94_s1_14\
        );

    \I__7814\ : InMux
    port map (
            O => \N__35223\,
            I => \N__35220\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__35220\,
            I => \N__35217\
        );

    \I__7812\ : Odrv4
    port map (
            O => \N__35217\,
            I => \b2v_inst11.un1_dutycycle_94_s0_14\
        );

    \I__7811\ : CascadeMux
    port map (
            O => \N__35214\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0_cascade_\
        );

    \I__7810\ : InMux
    port map (
            O => \N__35211\,
            I => \N__35206\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__35210\,
            I => \N__35200\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__35209\,
            I => \N__35196\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__35206\,
            I => \N__35190\
        );

    \I__7806\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35185\
        );

    \I__7805\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35182\
        );

    \I__7804\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35177\
        );

    \I__7803\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35177\
        );

    \I__7802\ : InMux
    port map (
            O => \N__35199\,
            I => \N__35170\
        );

    \I__7801\ : InMux
    port map (
            O => \N__35196\,
            I => \N__35170\
        );

    \I__7800\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35170\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__35194\,
            I => \N__35166\
        );

    \I__7798\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35163\
        );

    \I__7797\ : Span4Mux_v
    port map (
            O => \N__35190\,
            I => \N__35160\
        );

    \I__7796\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35157\
        );

    \I__7795\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35154\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__35185\,
            I => \N__35149\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__35182\,
            I => \N__35149\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35146\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__35143\
        );

    \I__7790\ : InMux
    port map (
            O => \N__35169\,
            I => \N__35138\
        );

    \I__7789\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35138\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__35163\,
            I => \N__35135\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__35160\,
            I => \N__35120\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__35157\,
            I => \N__35120\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__35154\,
            I => \N__35120\
        );

    \I__7784\ : Span4Mux_v
    port map (
            O => \N__35149\,
            I => \N__35120\
        );

    \I__7783\ : Span4Mux_h
    port map (
            O => \N__35146\,
            I => \N__35120\
        );

    \I__7782\ : Span4Mux_h
    port map (
            O => \N__35143\,
            I => \N__35120\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__35138\,
            I => \N__35120\
        );

    \I__7780\ : Odrv12
    port map (
            O => \N__35135\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__7779\ : Odrv4
    port map (
            O => \N__35120\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__7778\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__35112\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0\
        );

    \I__7776\ : InMux
    port map (
            O => \N__35109\,
            I => \N__35103\
        );

    \I__7775\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35103\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__7773\ : Odrv12
    port map (
            O => \N__35100\,
            I => \b2v_inst11.dutycycle_en_11\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__35097\,
            I => \N__35094\
        );

    \I__7771\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35088\
        );

    \I__7770\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35088\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__35088\,
            I => \b2v_inst11.dutycycleZ0Z_14\
        );

    \I__7768\ : CascadeMux
    port map (
            O => \N__35085\,
            I => \N__35080\
        );

    \I__7767\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35077\
        );

    \I__7766\ : CascadeMux
    port map (
            O => \N__35083\,
            I => \N__35074\
        );

    \I__7765\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35071\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__35077\,
            I => \N__35066\
        );

    \I__7763\ : InMux
    port map (
            O => \N__35074\,
            I => \N__35063\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__35071\,
            I => \N__35060\
        );

    \I__7761\ : InMux
    port map (
            O => \N__35070\,
            I => \N__35057\
        );

    \I__7760\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35054\
        );

    \I__7759\ : Span4Mux_v
    port map (
            O => \N__35066\,
            I => \N__35049\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__35063\,
            I => \N__35049\
        );

    \I__7757\ : Span4Mux_s3_v
    port map (
            O => \N__35060\,
            I => \N__35046\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__35057\,
            I => \N__35043\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__35054\,
            I => \N__35038\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__35049\,
            I => \N__35038\
        );

    \I__7753\ : Odrv4
    port map (
            O => \N__35046\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_10\
        );

    \I__7752\ : Odrv12
    port map (
            O => \N__35043\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_10\
        );

    \I__7751\ : Odrv4
    port map (
            O => \N__35038\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_10\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__35031\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_\
        );

    \I__7749\ : InMux
    port map (
            O => \N__35028\,
            I => \N__35020\
        );

    \I__7748\ : InMux
    port map (
            O => \N__35027\,
            I => \N__35020\
        );

    \I__7747\ : CascadeMux
    port map (
            O => \N__35026\,
            I => \N__35017\
        );

    \I__7746\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35012\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__35020\,
            I => \N__35003\
        );

    \I__7744\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34997\
        );

    \I__7743\ : InMux
    port map (
            O => \N__35016\,
            I => \N__34997\
        );

    \I__7742\ : InMux
    port map (
            O => \N__35015\,
            I => \N__34994\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__35012\,
            I => \N__34990\
        );

    \I__7740\ : InMux
    port map (
            O => \N__35011\,
            I => \N__34987\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__35010\,
            I => \N__34983\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__35009\,
            I => \N__34979\
        );

    \I__7737\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34969\
        );

    \I__7736\ : InMux
    port map (
            O => \N__35007\,
            I => \N__34969\
        );

    \I__7735\ : InMux
    port map (
            O => \N__35006\,
            I => \N__34969\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__35003\,
            I => \N__34966\
        );

    \I__7733\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34963\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__34997\,
            I => \N__34959\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__34994\,
            I => \N__34956\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__34993\,
            I => \N__34950\
        );

    \I__7729\ : Span4Mux_s3_h
    port map (
            O => \N__34990\,
            I => \N__34947\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34944\
        );

    \I__7727\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34941\
        );

    \I__7726\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34936\
        );

    \I__7725\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34936\
        );

    \I__7724\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34933\
        );

    \I__7723\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34926\
        );

    \I__7722\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34926\
        );

    \I__7721\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34926\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34923\
        );

    \I__7719\ : Sp12to4
    port map (
            O => \N__34966\,
            I => \N__34918\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34918\
        );

    \I__7717\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34915\
        );

    \I__7716\ : Span4Mux_s3_v
    port map (
            O => \N__34959\,
            I => \N__34910\
        );

    \I__7715\ : Span4Mux_s0_h
    port map (
            O => \N__34956\,
            I => \N__34910\
        );

    \I__7714\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34901\
        );

    \I__7713\ : InMux
    port map (
            O => \N__34954\,
            I => \N__34901\
        );

    \I__7712\ : InMux
    port map (
            O => \N__34953\,
            I => \N__34901\
        );

    \I__7711\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34901\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__34947\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7709\ : Odrv12
    port map (
            O => \N__34944\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__34941\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__34936\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__34933\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__34926\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7704\ : Odrv4
    port map (
            O => \N__34923\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7703\ : Odrv12
    port map (
            O => \N__34918\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__34915\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__34910\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__34901\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__7699\ : CascadeMux
    port map (
            O => \N__34878\,
            I => \b2v_inst11.un1_dutycycle_53_44_0_3_tz_1_cascade_\
        );

    \I__7698\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34871\
        );

    \I__7697\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34868\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34865\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__34868\,
            I => \N__34862\
        );

    \I__7694\ : Span4Mux_s3_v
    port map (
            O => \N__34865\,
            I => \N__34859\
        );

    \I__7693\ : Odrv4
    port map (
            O => \N__34862\,
            I => \b2v_inst11.un1_dutycycle_53_44_1\
        );

    \I__7692\ : Odrv4
    port map (
            O => \N__34859\,
            I => \b2v_inst11.un1_dutycycle_53_44_1\
        );

    \I__7691\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34851\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__34851\,
            I => \N__34848\
        );

    \I__7689\ : Span4Mux_s3_h
    port map (
            O => \N__34848\,
            I => \N__34845\
        );

    \I__7688\ : Odrv4
    port map (
            O => \N__34845\,
            I => \b2v_inst11.g3_0_0\
        );

    \I__7687\ : IoInMux
    port map (
            O => \N__34842\,
            I => \N__34839\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34834\
        );

    \I__7685\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34830\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__34837\,
            I => \N__34827\
        );

    \I__7683\ : IoSpan4Mux
    port map (
            O => \N__34834\,
            I => \N__34824\
        );

    \I__7682\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34820\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__34830\,
            I => \N__34814\
        );

    \I__7680\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34811\
        );

    \I__7679\ : IoSpan4Mux
    port map (
            O => \N__34824\,
            I => \N__34808\
        );

    \I__7678\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34805\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34802\
        );

    \I__7676\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34797\
        );

    \I__7675\ : CascadeMux
    port map (
            O => \N__34818\,
            I => \N__34794\
        );

    \I__7674\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34791\
        );

    \I__7673\ : Span4Mux_v
    port map (
            O => \N__34814\,
            I => \N__34786\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__34811\,
            I => \N__34786\
        );

    \I__7671\ : Span4Mux_s3_v
    port map (
            O => \N__34808\,
            I => \N__34781\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__34805\,
            I => \N__34781\
        );

    \I__7669\ : Span4Mux_s3_h
    port map (
            O => \N__34802\,
            I => \N__34778\
        );

    \I__7668\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34775\
        );

    \I__7667\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34772\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__34797\,
            I => \N__34766\
        );

    \I__7665\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34763\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__34791\,
            I => \N__34760\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__34786\,
            I => \N__34757\
        );

    \I__7662\ : Span4Mux_v
    port map (
            O => \N__34781\,
            I => \N__34748\
        );

    \I__7661\ : Span4Mux_h
    port map (
            O => \N__34778\,
            I => \N__34748\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__34775\,
            I => \N__34748\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__34772\,
            I => \N__34748\
        );

    \I__7658\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34741\
        );

    \I__7657\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34741\
        );

    \I__7656\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34741\
        );

    \I__7655\ : Span4Mux_s3_h
    port map (
            O => \N__34766\,
            I => \N__34738\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__34763\,
            I => rsmrstn
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__34760\,
            I => rsmrstn
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__34757\,
            I => rsmrstn
        );

    \I__7651\ : Odrv4
    port map (
            O => \N__34748\,
            I => rsmrstn
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__34741\,
            I => rsmrstn
        );

    \I__7649\ : Odrv4
    port map (
            O => \N__34738\,
            I => rsmrstn
        );

    \I__7648\ : CascadeMux
    port map (
            O => \N__34725\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_7_cascade_\
        );

    \I__7647\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34719\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__34719\,
            I => \b2v_inst11.g1_0_0\
        );

    \I__7645\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34713\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__34713\,
            I => \b2v_inst11.un1_clk_100khz_36_and_i_0_0\
        );

    \I__7643\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34707\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__34707\,
            I => \N__34704\
        );

    \I__7641\ : Span4Mux_s1_h
    port map (
            O => \N__34704\,
            I => \N__34701\
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__34701\,
            I => \b2v_inst11.un1_dutycycle_94_s1_7\
        );

    \I__7639\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34695\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34692\
        );

    \I__7637\ : Span4Mux_s0_h
    port map (
            O => \N__34692\,
            I => \N__34689\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__34689\,
            I => \b2v_inst11.un1_dutycycle_94_s0_7\
        );

    \I__7635\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34683\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__34683\,
            I => \b2v_inst11.un1_dutycycle_94_0_7\
        );

    \I__7633\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__34677\,
            I => \b2v_inst11.g0_0_1_0\
        );

    \I__7631\ : InMux
    port map (
            O => \N__34674\,
            I => \N__34668\
        );

    \I__7630\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34668\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__34668\,
            I => \b2v_inst11.dutycycleZ1Z_7\
        );

    \I__7628\ : CascadeMux
    port map (
            O => \N__34665\,
            I => \b2v_inst11.un1_dutycycle_94_0_7_cascade_\
        );

    \I__7627\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34659\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__34659\,
            I => \N__34656\
        );

    \I__7625\ : Span4Mux_s1_h
    port map (
            O => \N__34656\,
            I => \N__34653\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__34653\,
            I => \b2v_inst11.un1_dutycycle_94_s1_13\
        );

    \I__7623\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34647\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__34647\,
            I => \N__34644\
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__34644\,
            I => \b2v_inst11.un1_dutycycle_94_s0_13\
        );

    \I__7620\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34638\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__34638\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0\
        );

    \I__7618\ : CascadeMux
    port map (
            O => \N__34635\,
            I => \N__34632\
        );

    \I__7617\ : InMux
    port map (
            O => \N__34632\,
            I => \N__34626\
        );

    \I__7616\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34626\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__34626\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__7614\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34617\
        );

    \I__7613\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34617\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__34617\,
            I => \N__34614\
        );

    \I__7611\ : Odrv12
    port map (
            O => \N__34614\,
            I => \b2v_inst11.dutycycle_en_10\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__34611\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0_cascade_\
        );

    \I__7609\ : CascadeMux
    port map (
            O => \N__34608\,
            I => \N__34601\
        );

    \I__7608\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34595\
        );

    \I__7607\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34592\
        );

    \I__7606\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34588\
        );

    \I__7605\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34585\
        );

    \I__7604\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34580\
        );

    \I__7603\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34580\
        );

    \I__7602\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34575\
        );

    \I__7601\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34575\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__34595\,
            I => \N__34570\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__34592\,
            I => \N__34570\
        );

    \I__7598\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34564\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__34588\,
            I => \N__34560\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34557\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__34580\,
            I => \N__34552\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34552\
        );

    \I__7593\ : Span4Mux_v
    port map (
            O => \N__34570\,
            I => \N__34549\
        );

    \I__7592\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34544\
        );

    \I__7591\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34544\
        );

    \I__7590\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34541\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34538\
        );

    \I__7588\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34535\
        );

    \I__7587\ : Span4Mux_v
    port map (
            O => \N__34560\,
            I => \N__34528\
        );

    \I__7586\ : Span4Mux_v
    port map (
            O => \N__34557\,
            I => \N__34528\
        );

    \I__7585\ : Span4Mux_v
    port map (
            O => \N__34552\,
            I => \N__34528\
        );

    \I__7584\ : Span4Mux_s0_h
    port map (
            O => \N__34549\,
            I => \N__34521\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34521\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34521\
        );

    \I__7581\ : Odrv12
    port map (
            O => \N__34538\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__34535\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__34528\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__34521\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__34512\,
            I => \b2v_inst11.un1_clk_100khz_32_and_i_0_c_0_cascade_\
        );

    \I__7576\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34503\
        );

    \I__7575\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34503\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__34503\,
            I => \b2v_inst11.un1_clk_100khz_32_and_i_0_d\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__34500\,
            I => \b2v_inst11.un1_clk_100khz_33_and_i_0_c_0_cascade_\
        );

    \I__7572\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34494\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__34494\,
            I => \b2v_inst11.N_153_N\
        );

    \I__7570\ : CascadeMux
    port map (
            O => \N__34491\,
            I => \b2v_inst11.N_155_N_cascade_\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__34488\,
            I => \b2v_inst11.g0_0_1_0_cascade_\
        );

    \I__7568\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34482\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__34482\,
            I => \b2v_inst11.g0_1_1\
        );

    \I__7566\ : CascadeMux
    port map (
            O => \N__34479\,
            I => \b2v_inst11.dutycycle_set_1_cascade_\
        );

    \I__7565\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34473\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34470\
        );

    \I__7563\ : Span4Mux_s0_h
    port map (
            O => \N__34470\,
            I => \N__34467\
        );

    \I__7562\ : Span4Mux_h
    port map (
            O => \N__34467\,
            I => \N__34463\
        );

    \I__7561\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34460\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__34463\,
            I => \b2v_inst11.dutycycle_eena_14_0\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__34460\,
            I => \b2v_inst11.dutycycle_eena_14_0\
        );

    \I__7558\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34452\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__34452\,
            I => \N__34448\
        );

    \I__7556\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34445\
        );

    \I__7555\ : Span4Mux_h
    port map (
            O => \N__34448\,
            I => \N__34442\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__34445\,
            I => \b2v_inst11.dutycycle_0_5\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__34442\,
            I => \b2v_inst11.dutycycle_0_5\
        );

    \I__7552\ : CascadeMux
    port map (
            O => \N__34437\,
            I => \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3_cascade_\
        );

    \I__7551\ : InMux
    port map (
            O => \N__34434\,
            I => \N__34431\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__34431\,
            I => \N__34428\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__34428\,
            I => \N__34425\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__34425\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJZ0Z9\
        );

    \I__7547\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34419\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__34419\,
            I => \b2v_inst11.dutycycle_RNIM98E2Z0Z_3\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__34416\,
            I => \N__34413\
        );

    \I__7544\ : InMux
    port map (
            O => \N__34413\,
            I => \N__34408\
        );

    \I__7543\ : InMux
    port map (
            O => \N__34412\,
            I => \N__34403\
        );

    \I__7542\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34403\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__34408\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__34403\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__34398\,
            I => \b2v_inst11.dutycycle_RNIM98E2Z0Z_3_cascade_\
        );

    \I__7538\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34392\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__34392\,
            I => \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3\
        );

    \I__7536\ : InMux
    port map (
            O => \N__34389\,
            I => \N__34384\
        );

    \I__7535\ : InMux
    port map (
            O => \N__34388\,
            I => \N__34373\
        );

    \I__7534\ : InMux
    port map (
            O => \N__34387\,
            I => \N__34373\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__34384\,
            I => \N__34370\
        );

    \I__7532\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34363\
        );

    \I__7531\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34363\
        );

    \I__7530\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34357\
        );

    \I__7529\ : InMux
    port map (
            O => \N__34380\,
            I => \N__34357\
        );

    \I__7528\ : CascadeMux
    port map (
            O => \N__34379\,
            I => \N__34351\
        );

    \I__7527\ : InMux
    port map (
            O => \N__34378\,
            I => \N__34348\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34343\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__34370\,
            I => \N__34343\
        );

    \I__7524\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34338\
        );

    \I__7523\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34338\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__34363\,
            I => \N__34335\
        );

    \I__7521\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34332\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__34357\,
            I => \N__34329\
        );

    \I__7519\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34324\
        );

    \I__7518\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34324\
        );

    \I__7517\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34319\
        );

    \I__7516\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34316\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34309\
        );

    \I__7514\ : Span4Mux_h
    port map (
            O => \N__34343\,
            I => \N__34309\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__34338\,
            I => \N__34309\
        );

    \I__7512\ : Span4Mux_s3_v
    port map (
            O => \N__34335\,
            I => \N__34306\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__34332\,
            I => \N__34303\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__34329\,
            I => \N__34298\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__34324\,
            I => \N__34298\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__34323\,
            I => \N__34295\
        );

    \I__7507\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34292\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__34319\,
            I => \N__34285\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34285\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__34309\,
            I => \N__34285\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__34306\,
            I => \N__34278\
        );

    \I__7502\ : Span4Mux_h
    port map (
            O => \N__34303\,
            I => \N__34278\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__34298\,
            I => \N__34278\
        );

    \I__7500\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34275\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__34292\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__7498\ : Odrv4
    port map (
            O => \N__34285\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__34278\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__34275\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__7495\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34262\
        );

    \I__7494\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34255\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__34262\,
            I => \N__34252\
        );

    \I__7492\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34242\
        );

    \I__7491\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34242\
        );

    \I__7490\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34242\
        );

    \I__7489\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34242\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34235\
        );

    \I__7487\ : Span4Mux_s1_h
    port map (
            O => \N__34252\,
            I => \N__34235\
        );

    \I__7486\ : InMux
    port map (
            O => \N__34251\,
            I => \N__34232\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__34242\,
            I => \N__34229\
        );

    \I__7484\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34224\
        );

    \I__7483\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34224\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__34235\,
            I => \N__34221\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__34232\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__34229\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__34224\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__34221\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__34212\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3_cascade_\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__34209\,
            I => \N__34206\
        );

    \I__7475\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34203\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34200\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__34200\,
            I => \N__34197\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__34197\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_s0_sf\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__34194\,
            I => \N__34190\
        );

    \I__7470\ : CascadeMux
    port map (
            O => \N__34193\,
            I => \N__34184\
        );

    \I__7469\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34178\
        );

    \I__7468\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34178\
        );

    \I__7467\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34175\
        );

    \I__7466\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34170\
        );

    \I__7465\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34170\
        );

    \I__7464\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34167\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__34178\,
            I => \N__34156\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__34175\,
            I => \N__34156\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__34170\,
            I => \N__34156\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34156\
        );

    \I__7459\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34153\
        );

    \I__7458\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34150\
        );

    \I__7457\ : Span4Mux_v
    port map (
            O => \N__34156\,
            I => \N__34147\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__34153\,
            I => \N__34144\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__34150\,
            I => \N__34141\
        );

    \I__7454\ : Span4Mux_v
    port map (
            O => \N__34147\,
            I => \N__34136\
        );

    \I__7453\ : Span4Mux_v
    port map (
            O => \N__34144\,
            I => \N__34136\
        );

    \I__7452\ : Odrv12
    port map (
            O => \N__34141\,
            I => \b2v_inst11.count_clk_RNIG510TZ0Z_7\
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__34136\,
            I => \b2v_inst11.count_clk_RNIG510TZ0Z_7\
        );

    \I__7450\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__34128\,
            I => \N__34125\
        );

    \I__7448\ : Span4Mux_s0_h
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__34122\,
            I => \b2v_inst11.N_305\
        );

    \I__7446\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34116\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__34116\,
            I => \N__34113\
        );

    \I__7444\ : Odrv12
    port map (
            O => \N__34113\,
            I => \b2v_inst11.N_306\
        );

    \I__7443\ : CascadeMux
    port map (
            O => \N__34110\,
            I => \b2v_inst11.N_231_N_cascade_\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__34107\,
            I => \b2v_inst11.dutycycle_eena_13_cascade_\
        );

    \I__7441\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34101\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__34101\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4\
        );

    \I__7439\ : InMux
    port map (
            O => \N__34098\,
            I => \N__34092\
        );

    \I__7438\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34092\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__34092\,
            I => \b2v_inst11.dutycycle_0_6\
        );

    \I__7436\ : CascadeMux
    port map (
            O => \N__34089\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4_cascade_\
        );

    \I__7435\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34083\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__34083\,
            I => \b2v_inst11.dutycycle_eena_13\
        );

    \I__7433\ : InMux
    port map (
            O => \N__34080\,
            I => \N__34077\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__34077\,
            I => \N__34074\
        );

    \I__7431\ : Span4Mux_s2_h
    port map (
            O => \N__34074\,
            I => \N__34071\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__34071\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__34068\,
            I => \b2v_inst11.dutycycleZ1Z_6_cascade_\
        );

    \I__7428\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34062\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__34062\,
            I => \b2v_inst11.dutycycle_RNILF063Z0Z_6\
        );

    \I__7426\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34055\
        );

    \I__7425\ : InMux
    port map (
            O => \N__34058\,
            I => \N__34052\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__34055\,
            I => \N__34042\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__34052\,
            I => \N__34042\
        );

    \I__7422\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34037\
        );

    \I__7421\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34037\
        );

    \I__7420\ : CascadeMux
    port map (
            O => \N__34049\,
            I => \N__34033\
        );

    \I__7419\ : CascadeMux
    port map (
            O => \N__34048\,
            I => \N__34027\
        );

    \I__7418\ : CascadeMux
    port map (
            O => \N__34047\,
            I => \N__34021\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__34042\,
            I => \N__34018\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__34037\,
            I => \N__34015\
        );

    \I__7415\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34008\
        );

    \I__7414\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34008\
        );

    \I__7413\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34008\
        );

    \I__7412\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34005\
        );

    \I__7411\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34000\
        );

    \I__7410\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34000\
        );

    \I__7409\ : InMux
    port map (
            O => \N__34026\,
            I => \N__33995\
        );

    \I__7408\ : InMux
    port map (
            O => \N__34025\,
            I => \N__33995\
        );

    \I__7407\ : InMux
    port map (
            O => \N__34024\,
            I => \N__33992\
        );

    \I__7406\ : InMux
    port map (
            O => \N__34021\,
            I => \N__33989\
        );

    \I__7405\ : IoSpan4Mux
    port map (
            O => \N__34018\,
            I => \N__33984\
        );

    \I__7404\ : Span4Mux_h
    port map (
            O => \N__34015\,
            I => \N__33984\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__33981\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__33976\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__34000\,
            I => \N__33976\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__33995\,
            I => \N__33973\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__33992\,
            I => \N__33970\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__33989\,
            I => \N__33967\
        );

    \I__7397\ : Span4Mux_s1_h
    port map (
            O => \N__33984\,
            I => \N__33964\
        );

    \I__7396\ : Span4Mux_h
    port map (
            O => \N__33981\,
            I => \N__33961\
        );

    \I__7395\ : Span4Mux_v
    port map (
            O => \N__33976\,
            I => \N__33958\
        );

    \I__7394\ : Span12Mux_s1_h
    port map (
            O => \N__33973\,
            I => \N__33955\
        );

    \I__7393\ : Odrv12
    port map (
            O => \N__33970\,
            I => \b2v_inst11.N_172\
        );

    \I__7392\ : Odrv12
    port map (
            O => \N__33967\,
            I => \b2v_inst11.N_172\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__33964\,
            I => \b2v_inst11.N_172\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__33961\,
            I => \b2v_inst11.N_172\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__33958\,
            I => \b2v_inst11.N_172\
        );

    \I__7388\ : Odrv12
    port map (
            O => \N__33955\,
            I => \b2v_inst11.N_172\
        );

    \I__7387\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33935\
        );

    \I__7386\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33935\
        );

    \I__7385\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33932\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__33935\,
            I => \N__33929\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__33932\,
            I => \b2v_inst11.N_185\
        );

    \I__7382\ : Odrv12
    port map (
            O => \N__33929\,
            I => \b2v_inst11.N_185\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__33924\,
            I => \N__33921\
        );

    \I__7380\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33918\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__33918\,
            I => \N__33915\
        );

    \I__7378\ : Span4Mux_h
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__33912\,
            I => \b2v_inst11.dutycycle_set_1\
        );

    \I__7376\ : InMux
    port map (
            O => \N__33909\,
            I => \N__33906\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__33906\,
            I => \N__33902\
        );

    \I__7374\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33899\
        );

    \I__7373\ : Odrv4
    port map (
            O => \N__33902\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__33899\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__7371\ : InMux
    port map (
            O => \N__33894\,
            I => \N__33888\
        );

    \I__7370\ : InMux
    port map (
            O => \N__33893\,
            I => \N__33888\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__33888\,
            I => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\
        );

    \I__7368\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33882\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__33882\,
            I => \b2v_inst11.count_clk_0_15\
        );

    \I__7366\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33876\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__33876\,
            I => \N__33873\
        );

    \I__7364\ : Span4Mux_h
    port map (
            O => \N__33873\,
            I => \N__33870\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__33870\,
            I => \N__33866\
        );

    \I__7362\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33863\
        );

    \I__7361\ : Span4Mux_v
    port map (
            O => \N__33866\,
            I => \N__33860\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__33863\,
            I => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__33860\,
            I => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\
        );

    \I__7358\ : InMux
    port map (
            O => \N__33855\,
            I => \N__33852\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__33852\,
            I => \N__33849\
        );

    \I__7356\ : Span4Mux_s1_h
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__33846\,
            I => \N__33843\
        );

    \I__7354\ : Span4Mux_h
    port map (
            O => \N__33843\,
            I => \N__33840\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__33840\,
            I => \b2v_inst11.count_clk_0_6\
        );

    \I__7352\ : CEMux
    port map (
            O => \N__33837\,
            I => \N__33832\
        );

    \I__7351\ : CEMux
    port map (
            O => \N__33836\,
            I => \N__33827\
        );

    \I__7350\ : CEMux
    port map (
            O => \N__33835\,
            I => \N__33819\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__33832\,
            I => \N__33816\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__33831\,
            I => \N__33813\
        );

    \I__7347\ : CascadeMux
    port map (
            O => \N__33830\,
            I => \N__33804\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33798\
        );

    \I__7345\ : CascadeMux
    port map (
            O => \N__33826\,
            I => \N__33793\
        );

    \I__7344\ : CascadeMux
    port map (
            O => \N__33825\,
            I => \N__33790\
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__33824\,
            I => \N__33787\
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__33823\,
            I => \N__33783\
        );

    \I__7341\ : CEMux
    port map (
            O => \N__33822\,
            I => \N__33780\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33777\
        );

    \I__7339\ : Span4Mux_h
    port map (
            O => \N__33816\,
            I => \N__33774\
        );

    \I__7338\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33769\
        );

    \I__7337\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33769\
        );

    \I__7336\ : CascadeMux
    port map (
            O => \N__33811\,
            I => \N__33764\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__33810\,
            I => \N__33760\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__33809\,
            I => \N__33757\
        );

    \I__7333\ : CEMux
    port map (
            O => \N__33808\,
            I => \N__33753\
        );

    \I__7332\ : InMux
    port map (
            O => \N__33807\,
            I => \N__33744\
        );

    \I__7331\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33744\
        );

    \I__7330\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33744\
        );

    \I__7329\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33744\
        );

    \I__7328\ : CEMux
    port map (
            O => \N__33801\,
            I => \N__33741\
        );

    \I__7327\ : Span4Mux_v
    port map (
            O => \N__33798\,
            I => \N__33738\
        );

    \I__7326\ : CEMux
    port map (
            O => \N__33797\,
            I => \N__33733\
        );

    \I__7325\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33733\
        );

    \I__7324\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33719\
        );

    \I__7323\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33719\
        );

    \I__7322\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33719\
        );

    \I__7321\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33719\
        );

    \I__7320\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33719\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33716\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__33777\,
            I => \N__33711\
        );

    \I__7317\ : Span4Mux_h
    port map (
            O => \N__33774\,
            I => \N__33711\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__33769\,
            I => \N__33708\
        );

    \I__7315\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33695\
        );

    \I__7314\ : CEMux
    port map (
            O => \N__33767\,
            I => \N__33695\
        );

    \I__7313\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33695\
        );

    \I__7312\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33695\
        );

    \I__7311\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33695\
        );

    \I__7310\ : InMux
    port map (
            O => \N__33757\,
            I => \N__33695\
        );

    \I__7309\ : CEMux
    port map (
            O => \N__33756\,
            I => \N__33692\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__33753\,
            I => \N__33689\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33686\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33681\
        );

    \I__7305\ : Span4Mux_h
    port map (
            O => \N__33738\,
            I => \N__33681\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__33733\,
            I => \N__33678\
        );

    \I__7303\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33671\
        );

    \I__7302\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33671\
        );

    \I__7301\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33671\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33668\
        );

    \I__7299\ : Span4Mux_s0_h
    port map (
            O => \N__33716\,
            I => \N__33659\
        );

    \I__7298\ : Span4Mux_v
    port map (
            O => \N__33711\,
            I => \N__33659\
        );

    \I__7297\ : Span4Mux_h
    port map (
            O => \N__33708\,
            I => \N__33659\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33659\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__33692\,
            I => \N__33652\
        );

    \I__7294\ : Span4Mux_h
    port map (
            O => \N__33689\,
            I => \N__33652\
        );

    \I__7293\ : Span4Mux_h
    port map (
            O => \N__33686\,
            I => \N__33652\
        );

    \I__7292\ : Odrv4
    port map (
            O => \N__33681\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__7291\ : Odrv12
    port map (
            O => \N__33678\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__33671\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__33668\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__33659\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__7287\ : Odrv4
    port map (
            O => \N__33652\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__7286\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33635\
        );

    \I__7285\ : InMux
    port map (
            O => \N__33638\,
            I => \N__33632\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__33635\,
            I => \N__33626\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__33632\,
            I => \N__33626\
        );

    \I__7282\ : CascadeMux
    port map (
            O => \N__33631\,
            I => \N__33623\
        );

    \I__7281\ : Span4Mux_h
    port map (
            O => \N__33626\,
            I => \N__33620\
        );

    \I__7280\ : InMux
    port map (
            O => \N__33623\,
            I => \N__33617\
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__33620\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__33617\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__7277\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33608\
        );

    \I__7276\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33605\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__33608\,
            I => \N__33602\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__33605\,
            I => \N__33599\
        );

    \I__7273\ : Span4Mux_s3_h
    port map (
            O => \N__33602\,
            I => \N__33596\
        );

    \I__7272\ : Odrv4
    port map (
            O => \N__33599\,
            I => \b2v_inst6.N_241\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__33596\,
            I => \b2v_inst6.N_241\
        );

    \I__7270\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33585\
        );

    \I__7269\ : CascadeMux
    port map (
            O => \N__33590\,
            I => \N__33582\
        );

    \I__7268\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33577\
        );

    \I__7267\ : InMux
    port map (
            O => \N__33588\,
            I => \N__33577\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__33585\,
            I => \N__33574\
        );

    \I__7265\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33571\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__33577\,
            I => \N__33568\
        );

    \I__7263\ : Span4Mux_s2_h
    port map (
            O => \N__33574\,
            I => \N__33565\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__33571\,
            I => \N__33560\
        );

    \I__7261\ : Span4Mux_s1_v
    port map (
            O => \N__33568\,
            I => \N__33560\
        );

    \I__7260\ : Span4Mux_v
    port map (
            O => \N__33565\,
            I => \N__33557\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__33560\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__33557\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7257\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33546\
        );

    \I__7256\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33546\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__33546\,
            I => \N__33543\
        );

    \I__7254\ : Span4Mux_s2_v
    port map (
            O => \N__33543\,
            I => \N__33540\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__33540\,
            I => \N__33537\
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__33537\,
            I => \b2v_inst6.N_2994_i\
        );

    \I__7251\ : CascadeMux
    port map (
            O => \N__33534\,
            I => \b2v_inst6.N_2994_i_cascade_\
        );

    \I__7250\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33526\
        );

    \I__7249\ : InMux
    port map (
            O => \N__33530\,
            I => \N__33521\
        );

    \I__7248\ : InMux
    port map (
            O => \N__33529\,
            I => \N__33521\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__33526\,
            I => \N__33518\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__33521\,
            I => \N__33515\
        );

    \I__7245\ : Odrv12
    port map (
            O => \N__33518\,
            I => \b2v_inst6.N_389\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__33515\,
            I => \b2v_inst6.N_389\
        );

    \I__7243\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__33507\,
            I => \N__33504\
        );

    \I__7241\ : Span4Mux_s2_v
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__7240\ : Span4Mux_v
    port map (
            O => \N__33501\,
            I => \N__33498\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__33495\,
            I => \b2v_inst6.count_0_0\
        );

    \I__7237\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__33489\,
            I => \N__33485\
        );

    \I__7235\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33482\
        );

    \I__7234\ : Span4Mux_v
    port map (
            O => \N__33485\,
            I => \N__33479\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__33482\,
            I => \b2v_inst6.count_rst\
        );

    \I__7232\ : Odrv4
    port map (
            O => \N__33479\,
            I => \b2v_inst6.count_rst\
        );

    \I__7231\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33471\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__33471\,
            I => \N__33468\
        );

    \I__7229\ : Odrv12
    port map (
            O => \N__33468\,
            I => \b2v_inst6.count_0_15\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__33465\,
            I => \N__33447\
        );

    \I__7227\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33438\
        );

    \I__7226\ : CEMux
    port map (
            O => \N__33463\,
            I => \N__33438\
        );

    \I__7225\ : InMux
    port map (
            O => \N__33462\,
            I => \N__33435\
        );

    \I__7224\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33430\
        );

    \I__7223\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33430\
        );

    \I__7222\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33427\
        );

    \I__7221\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33422\
        );

    \I__7220\ : CEMux
    port map (
            O => \N__33457\,
            I => \N__33422\
        );

    \I__7219\ : CEMux
    port map (
            O => \N__33456\,
            I => \N__33419\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__33455\,
            I => \N__33414\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__33454\,
            I => \N__33411\
        );

    \I__7216\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33398\
        );

    \I__7215\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33398\
        );

    \I__7214\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33398\
        );

    \I__7213\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33398\
        );

    \I__7212\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33389\
        );

    \I__7211\ : InMux
    port map (
            O => \N__33446\,
            I => \N__33389\
        );

    \I__7210\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33389\
        );

    \I__7209\ : CEMux
    port map (
            O => \N__33444\,
            I => \N__33389\
        );

    \I__7208\ : CascadeMux
    port map (
            O => \N__33443\,
            I => \N__33380\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__33438\,
            I => \N__33374\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__33435\,
            I => \N__33367\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__33430\,
            I => \N__33367\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__33427\,
            I => \N__33367\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33364\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__33419\,
            I => \N__33361\
        );

    \I__7201\ : CEMux
    port map (
            O => \N__33418\,
            I => \N__33358\
        );

    \I__7200\ : CEMux
    port map (
            O => \N__33417\,
            I => \N__33355\
        );

    \I__7199\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33350\
        );

    \I__7198\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33350\
        );

    \I__7197\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33347\
        );

    \I__7196\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33342\
        );

    \I__7195\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33342\
        );

    \I__7194\ : CEMux
    port map (
            O => \N__33407\,
            I => \N__33337\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__33398\,
            I => \N__33334\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__33389\,
            I => \N__33331\
        );

    \I__7191\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33326\
        );

    \I__7190\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33326\
        );

    \I__7189\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33319\
        );

    \I__7188\ : CEMux
    port map (
            O => \N__33385\,
            I => \N__33319\
        );

    \I__7187\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33319\
        );

    \I__7186\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33308\
        );

    \I__7185\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33308\
        );

    \I__7184\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33308\
        );

    \I__7183\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33308\
        );

    \I__7182\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33308\
        );

    \I__7181\ : Span4Mux_s2_v
    port map (
            O => \N__33374\,
            I => \N__33305\
        );

    \I__7180\ : Span4Mux_s2_v
    port map (
            O => \N__33367\,
            I => \N__33302\
        );

    \I__7179\ : Span4Mux_v
    port map (
            O => \N__33364\,
            I => \N__33297\
        );

    \I__7178\ : Span4Mux_s2_v
    port map (
            O => \N__33361\,
            I => \N__33297\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__33358\,
            I => \N__33288\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__33355\,
            I => \N__33288\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33288\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__33347\,
            I => \N__33288\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__33342\,
            I => \N__33285\
        );

    \I__7172\ : InMux
    port map (
            O => \N__33341\,
            I => \N__33280\
        );

    \I__7171\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33280\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__33337\,
            I => \N__33277\
        );

    \I__7169\ : Span12Mux_s6_v
    port map (
            O => \N__33334\,
            I => \N__33274\
        );

    \I__7168\ : Sp12to4
    port map (
            O => \N__33331\,
            I => \N__33265\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__33326\,
            I => \N__33265\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33265\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__33308\,
            I => \N__33265\
        );

    \I__7164\ : Span4Mux_v
    port map (
            O => \N__33305\,
            I => \N__33260\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__33302\,
            I => \N__33260\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__33297\,
            I => \N__33251\
        );

    \I__7161\ : Span4Mux_s2_v
    port map (
            O => \N__33288\,
            I => \N__33251\
        );

    \I__7160\ : Span4Mux_s2_v
    port map (
            O => \N__33285\,
            I => \N__33251\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__33280\,
            I => \N__33251\
        );

    \I__7158\ : Odrv4
    port map (
            O => \N__33277\,
            I => \b2v_inst6.count_en\
        );

    \I__7157\ : Odrv12
    port map (
            O => \N__33274\,
            I => \b2v_inst6.count_en\
        );

    \I__7156\ : Odrv12
    port map (
            O => \N__33265\,
            I => \b2v_inst6.count_en\
        );

    \I__7155\ : Odrv4
    port map (
            O => \N__33260\,
            I => \b2v_inst6.count_en\
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__33251\,
            I => \b2v_inst6.count_en\
        );

    \I__7153\ : SRMux
    port map (
            O => \N__33240\,
            I => \N__33232\
        );

    \I__7152\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33224\
        );

    \I__7151\ : SRMux
    port map (
            O => \N__33238\,
            I => \N__33224\
        );

    \I__7150\ : SRMux
    port map (
            O => \N__33237\,
            I => \N__33213\
        );

    \I__7149\ : SRMux
    port map (
            O => \N__33236\,
            I => \N__33210\
        );

    \I__7148\ : CascadeMux
    port map (
            O => \N__33235\,
            I => \N__33205\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__33232\,
            I => \N__33199\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__33231\,
            I => \N__33192\
        );

    \I__7145\ : CascadeMux
    port map (
            O => \N__33230\,
            I => \N__33189\
        );

    \I__7144\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33183\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33180\
        );

    \I__7142\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33175\
        );

    \I__7141\ : SRMux
    port map (
            O => \N__33222\,
            I => \N__33175\
        );

    \I__7140\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33164\
        );

    \I__7139\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33164\
        );

    \I__7138\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33164\
        );

    \I__7137\ : InMux
    port map (
            O => \N__33218\,
            I => \N__33164\
        );

    \I__7136\ : InMux
    port map (
            O => \N__33217\,
            I => \N__33164\
        );

    \I__7135\ : SRMux
    port map (
            O => \N__33216\,
            I => \N__33152\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__33213\,
            I => \N__33147\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__33210\,
            I => \N__33147\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__33209\,
            I => \N__33144\
        );

    \I__7131\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33126\
        );

    \I__7130\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33126\
        );

    \I__7129\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33126\
        );

    \I__7128\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33126\
        );

    \I__7127\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33126\
        );

    \I__7126\ : Span4Mux_s2_h
    port map (
            O => \N__33199\,
            I => \N__33123\
        );

    \I__7125\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33118\
        );

    \I__7124\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33118\
        );

    \I__7123\ : SRMux
    port map (
            O => \N__33196\,
            I => \N__33107\
        );

    \I__7122\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33107\
        );

    \I__7121\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33107\
        );

    \I__7120\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33107\
        );

    \I__7119\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33107\
        );

    \I__7118\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33102\
        );

    \I__7117\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33102\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33098\
        );

    \I__7115\ : Span4Mux_v
    port map (
            O => \N__33180\,
            I => \N__33093\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__33175\,
            I => \N__33093\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__33164\,
            I => \N__33090\
        );

    \I__7112\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33085\
        );

    \I__7111\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33085\
        );

    \I__7110\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33076\
        );

    \I__7109\ : SRMux
    port map (
            O => \N__33160\,
            I => \N__33076\
        );

    \I__7108\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33076\
        );

    \I__7107\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33076\
        );

    \I__7106\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33069\
        );

    \I__7105\ : InMux
    port map (
            O => \N__33156\,
            I => \N__33069\
        );

    \I__7104\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33069\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__33152\,
            I => \N__33066\
        );

    \I__7102\ : Span4Mux_s3_v
    port map (
            O => \N__33147\,
            I => \N__33063\
        );

    \I__7101\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33054\
        );

    \I__7100\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33054\
        );

    \I__7099\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33054\
        );

    \I__7098\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33054\
        );

    \I__7097\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33045\
        );

    \I__7096\ : InMux
    port map (
            O => \N__33139\,
            I => \N__33045\
        );

    \I__7095\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33045\
        );

    \I__7094\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33045\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__33126\,
            I => \N__33042\
        );

    \I__7092\ : Span4Mux_s0_v
    port map (
            O => \N__33123\,
            I => \N__33033\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33033\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__33107\,
            I => \N__33033\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__33102\,
            I => \N__33033\
        );

    \I__7088\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33030\
        );

    \I__7087\ : Span4Mux_v
    port map (
            O => \N__33098\,
            I => \N__33025\
        );

    \I__7086\ : Span4Mux_s2_v
    port map (
            O => \N__33093\,
            I => \N__33025\
        );

    \I__7085\ : Span4Mux_s2_h
    port map (
            O => \N__33090\,
            I => \N__33022\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__33085\,
            I => \N__33015\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33015\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33015\
        );

    \I__7081\ : Span4Mux_s3_h
    port map (
            O => \N__33066\,
            I => \N__33006\
        );

    \I__7080\ : Span4Mux_s3_h
    port map (
            O => \N__33063\,
            I => \N__33006\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33006\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__33006\
        );

    \I__7077\ : Span4Mux_s2_h
    port map (
            O => \N__33042\,
            I => \N__33003\
        );

    \I__7076\ : Span4Mux_s2_h
    port map (
            O => \N__33033\,
            I => \N__33000\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__33030\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__33025\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7073\ : Odrv4
    port map (
            O => \N__33022\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7072\ : Odrv12
    port map (
            O => \N__33015\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7071\ : Odrv4
    port map (
            O => \N__33006\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__33003\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7069\ : Odrv4
    port map (
            O => \N__33000\,
            I => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__7067\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32979\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32976\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__32976\,
            I => \b2v_inst11.func_state_RNI_4Z0Z_1\
        );

    \I__7064\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32970\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__32970\,
            I => \b2v_inst11.un1_count_clk_2_axb_5\
        );

    \I__7062\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32961\
        );

    \I__7061\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32961\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__32961\,
            I => \b2v_inst11.count_clk_0_5\
        );

    \I__7059\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32949\
        );

    \I__7058\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32949\
        );

    \I__7057\ : InMux
    port map (
            O => \N__32956\,
            I => \N__32949\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__32949\,
            I => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__32946\,
            I => \N__32941\
        );

    \I__7054\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32934\
        );

    \I__7053\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32934\
        );

    \I__7052\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32934\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__7050\ : Odrv12
    port map (
            O => \N__32931\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__7049\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32921\
        );

    \I__7047\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32918\
        );

    \I__7046\ : Span4Mux_s1_h
    port map (
            O => \N__32921\,
            I => \N__32915\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__32918\,
            I => \b2v_inst11.count_clk_0_7\
        );

    \I__7044\ : Odrv4
    port map (
            O => \N__32915\,
            I => \b2v_inst11.count_clk_0_7\
        );

    \I__7043\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32904\
        );

    \I__7042\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32904\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32900\
        );

    \I__7040\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32897\
        );

    \I__7039\ : Odrv4
    port map (
            O => \N__32900\,
            I => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__32897\,
            I => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\
        );

    \I__7037\ : CascadeMux
    port map (
            O => \N__32892\,
            I => \N__32889\
        );

    \I__7036\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32886\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__32886\,
            I => \b2v_inst11.un1_count_clk_2_axb_7\
        );

    \I__7034\ : CascadeMux
    port map (
            O => \N__32883\,
            I => \N__32880\
        );

    \I__7033\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32874\
        );

    \I__7032\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32874\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__32874\,
            I => \N__32870\
        );

    \I__7030\ : CascadeMux
    port map (
            O => \N__32873\,
            I => \N__32867\
        );

    \I__7029\ : Span4Mux_v
    port map (
            O => \N__32870\,
            I => \N__32864\
        );

    \I__7028\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32861\
        );

    \I__7027\ : Odrv4
    port map (
            O => \N__32864\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__32861\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__7025\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32850\
        );

    \I__7024\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32850\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__32850\,
            I => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\
        );

    \I__7022\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32844\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__32844\,
            I => \b2v_inst11.count_clk_0_4\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__32841\,
            I => \N__32838\
        );

    \I__7019\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32835\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__32835\,
            I => \b2v_inst11.un1_count_clk_2_axb_2\
        );

    \I__7017\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32826\
        );

    \I__7016\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32826\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__32826\,
            I => \b2v_inst11.count_clk_0_2\
        );

    \I__7014\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32814\
        );

    \I__7013\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32814\
        );

    \I__7012\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32814\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__32814\,
            I => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\
        );

    \I__7010\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32805\
        );

    \I__7009\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32805\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32802\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__32799\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__7005\ : CascadeMux
    port map (
            O => \N__32796\,
            I => \N__32792\
        );

    \I__7004\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32784\
        );

    \I__7003\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32784\
        );

    \I__7002\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32784\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__32784\,
            I => \b2v_inst6.un2_count_1_cry_9_c_RNIVIZ0Z14\
        );

    \I__7000\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32778\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__32778\,
            I => \b2v_inst6.count_rst_4\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__32775\,
            I => \N__32772\
        );

    \I__6997\ : InMux
    port map (
            O => \N__32772\,
            I => \N__32769\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__32769\,
            I => \b2v_inst6.countZ0Z_15\
        );

    \I__6995\ : CascadeMux
    port map (
            O => \N__32766\,
            I => \N__32763\
        );

    \I__6994\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32759\
        );

    \I__6993\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32756\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__32759\,
            I => \b2v_inst6.count_0_13\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__32756\,
            I => \b2v_inst6.count_0_13\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__32751\,
            I => \b2v_inst6.countZ0Z_15_cascade_\
        );

    \I__6989\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32745\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__32745\,
            I => \N__32742\
        );

    \I__6987\ : Odrv4
    port map (
            O => \N__32742\,
            I => \b2v_inst6.count_1_i_a3_2_0\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__32739\,
            I => \N__32735\
        );

    \I__6985\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32729\
        );

    \I__6984\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32729\
        );

    \I__6983\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32726\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__32729\,
            I => \b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__32726\,
            I => \b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0\
        );

    \I__6980\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32718\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__32718\,
            I => \b2v_inst6.count_rst_1\
        );

    \I__6978\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__32712\,
            I => \b2v_inst11.un1_count_clk_2_axb_12\
        );

    \I__6976\ : CascadeMux
    port map (
            O => \N__32709\,
            I => \N__32706\
        );

    \I__6975\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32703\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32698\
        );

    \I__6973\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32693\
        );

    \I__6972\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32693\
        );

    \I__6971\ : Odrv4
    port map (
            O => \N__32698\,
            I => \b2v_inst11.count_clk_1_12\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__32693\,
            I => \b2v_inst11.count_clk_1_12\
        );

    \I__6969\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32684\
        );

    \I__6968\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32681\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__32684\,
            I => \b2v_inst11.count_clk_0_12\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__32681\,
            I => \b2v_inst11.count_clk_0_12\
        );

    \I__6965\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32673\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__32673\,
            I => \b2v_inst11.un1_count_clk_2_axb_13\
        );

    \I__6963\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32667\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32662\
        );

    \I__6961\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32657\
        );

    \I__6960\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32657\
        );

    \I__6959\ : Odrv4
    port map (
            O => \N__32662\,
            I => \b2v_inst11.count_clk_1_13\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__32657\,
            I => \b2v_inst11.count_clk_1_13\
        );

    \I__6957\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32648\
        );

    \I__6956\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32645\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__32648\,
            I => \b2v_inst11.count_clk_0_13\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__32645\,
            I => \b2v_inst11.count_clk_0_13\
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__32640\,
            I => \b2v_inst6.countZ0Z_6_cascade_\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__32637\,
            I => \b2v_inst6.count_1_i_a3_0_0_cascade_\
        );

    \I__6951\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32631\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__32631\,
            I => \b2v_inst6.count_1_i_a3_7_0\
        );

    \I__6949\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32622\
        );

    \I__6948\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32622\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__32622\,
            I => \b2v_inst6.count_0_6\
        );

    \I__6946\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32615\
        );

    \I__6945\ : CascadeMux
    port map (
            O => \N__32618\,
            I => \N__32612\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__32615\,
            I => \N__32608\
        );

    \I__6943\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32603\
        );

    \I__6942\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32603\
        );

    \I__6941\ : Odrv4
    port map (
            O => \N__32608\,
            I => \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__32603\,
            I => \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__32598\,
            I => \N__32595\
        );

    \I__6938\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32592\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__32592\,
            I => \b2v_inst6.un2_count_1_axb_6\
        );

    \I__6936\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32586\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__32586\,
            I => \b2v_inst6.count_rst_2\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__32583\,
            I => \N__32579\
        );

    \I__6933\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32574\
        );

    \I__6932\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32574\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__32574\,
            I => \b2v_inst6.count_0_12\
        );

    \I__6930\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32562\
        );

    \I__6929\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32562\
        );

    \I__6928\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32562\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__32562\,
            I => \b2v_inst6.un2_count_1_cry_11_c_RNI8RABZ0\
        );

    \I__6926\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32556\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__32556\,
            I => \b2v_inst6.un2_count_1_axb_12\
        );

    \I__6924\ : InMux
    port map (
            O => \N__32553\,
            I => \N__32550\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__32550\,
            I => \b2v_inst6.un2_count_1_axb_10\
        );

    \I__6922\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32543\
        );

    \I__6921\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32540\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__32543\,
            I => \b2v_inst6.count_0_10\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__32540\,
            I => \b2v_inst6.count_0_10\
        );

    \I__6918\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32529\
        );

    \I__6917\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32529\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__32529\,
            I => \b2v_inst6.count_0_14\
        );

    \I__6915\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32517\
        );

    \I__6914\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32517\
        );

    \I__6913\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32517\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__32517\,
            I => \b2v_inst6.un2_count_1_cry_13_c_RNIR6IOZ0Z5\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__32514\,
            I => \N__32511\
        );

    \I__6910\ : InMux
    port map (
            O => \N__32511\,
            I => \N__32508\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__32508\,
            I => \b2v_inst6.un2_count_1_axb_14\
        );

    \I__6908\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32502\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__32502\,
            I => \b2v_inst6.countZ0Z_14\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__32499\,
            I => \b2v_inst6.count_rst_12_cascade_\
        );

    \I__6905\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32493\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__32493\,
            I => \N__32490\
        );

    \I__6903\ : Odrv4
    port map (
            O => \N__32490\,
            I => \b2v_inst6.count_1_i_a3_12_0\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__32487\,
            I => \b2v_inst6.count_1_i_a3_1_0_cascade_\
        );

    \I__6901\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32478\
        );

    \I__6900\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32478\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__32478\,
            I => \b2v_inst6.count_0_2\
        );

    \I__6898\ : CascadeMux
    port map (
            O => \N__32475\,
            I => \N__32471\
        );

    \I__6897\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32463\
        );

    \I__6896\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32463\
        );

    \I__6895\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32463\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__32463\,
            I => \b2v_inst6.un2_count_1_cry_1_c_RNIN2PZ0Z3\
        );

    \I__6893\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32457\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__32457\,
            I => \b2v_inst6.un2_count_1_axb_2\
        );

    \I__6891\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__32451\,
            I => \b2v_inst6.count_rst_7\
        );

    \I__6889\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32444\
        );

    \I__6888\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32441\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__32444\,
            I => \b2v_inst6.count_0_7\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__32441\,
            I => \b2v_inst6.count_0_7\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__32436\,
            I => \b2v_inst6.countZ0Z_5_cascade_\
        );

    \I__6884\ : CascadeMux
    port map (
            O => \N__32433\,
            I => \b2v_inst6.count_RNICV5H1Z0Z_1_cascade_\
        );

    \I__6883\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32426\
        );

    \I__6882\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32423\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__32426\,
            I => \b2v_inst6.un2_count_1_axb_1\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__32423\,
            I => \b2v_inst6.un2_count_1_axb_1\
        );

    \I__6879\ : CascadeMux
    port map (
            O => \N__32418\,
            I => \b2v_inst6.un2_count_1_axb_1_cascade_\
        );

    \I__6878\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32412\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__32412\,
            I => \b2v_inst6.count_RNICV5H1Z0Z_1\
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__32409\,
            I => \N__32405\
        );

    \I__6875\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32401\
        );

    \I__6874\ : InMux
    port map (
            O => \N__32405\,
            I => \N__32398\
        );

    \I__6873\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32395\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__32401\,
            I => \N__32392\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__32398\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__32395\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__32392\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6868\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32379\
        );

    \I__6867\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32379\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__32379\,
            I => \b2v_inst6.count_0_1\
        );

    \I__6865\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__32373\,
            I => \N__32370\
        );

    \I__6863\ : Odrv12
    port map (
            O => \N__32370\,
            I => \b2v_inst6.count_1_i_a3_4_0\
        );

    \I__6862\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__6860\ : Odrv12
    port map (
            O => \N__32361\,
            I => \b2v_inst6.count_1_i_a3_6_0\
        );

    \I__6859\ : CascadeMux
    port map (
            O => \N__32358\,
            I => \b2v_inst6.count_1_i_a3_3_0_cascade_\
        );

    \I__6858\ : InMux
    port map (
            O => \N__32355\,
            I => \N__32352\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__32352\,
            I => \b2v_inst6.count_1_i_a3_5_0\
        );

    \I__6856\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32343\
        );

    \I__6855\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32343\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__32343\,
            I => \b2v_inst6.count_0_5\
        );

    \I__6853\ : InMux
    port map (
            O => \N__32340\,
            I => \N__32334\
        );

    \I__6852\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32334\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__32334\,
            I => \b2v_inst6.count_rst_9\
        );

    \I__6850\ : CascadeMux
    port map (
            O => \N__32331\,
            I => \N__32327\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__32330\,
            I => \N__32324\
        );

    \I__6848\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32318\
        );

    \I__6847\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32318\
        );

    \I__6846\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32315\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__32318\,
            I => \b2v_inst6.un2_count_1_axb_5\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__32315\,
            I => \b2v_inst6.un2_count_1_axb_5\
        );

    \I__6843\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32298\
        );

    \I__6842\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32289\
        );

    \I__6841\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32286\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__32307\,
            I => \N__32279\
        );

    \I__6839\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32270\
        );

    \I__6838\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32263\
        );

    \I__6837\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32260\
        );

    \I__6836\ : InMux
    port map (
            O => \N__32303\,
            I => \N__32253\
        );

    \I__6835\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32253\
        );

    \I__6834\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32253\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__32298\,
            I => \N__32250\
        );

    \I__6832\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32243\
        );

    \I__6831\ : InMux
    port map (
            O => \N__32296\,
            I => \N__32243\
        );

    \I__6830\ : InMux
    port map (
            O => \N__32295\,
            I => \N__32234\
        );

    \I__6829\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32234\
        );

    \I__6828\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32234\
        );

    \I__6827\ : InMux
    port map (
            O => \N__32292\,
            I => \N__32234\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__32289\,
            I => \N__32229\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__32286\,
            I => \N__32229\
        );

    \I__6824\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32226\
        );

    \I__6823\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32217\
        );

    \I__6822\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32217\
        );

    \I__6821\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32217\
        );

    \I__6820\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32217\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__32278\,
            I => \N__32214\
        );

    \I__6818\ : InMux
    port map (
            O => \N__32277\,
            I => \N__32205\
        );

    \I__6817\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32205\
        );

    \I__6816\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32205\
        );

    \I__6815\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32205\
        );

    \I__6814\ : CascadeMux
    port map (
            O => \N__32273\,
            I => \N__32200\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__32270\,
            I => \N__32193\
        );

    \I__6812\ : InMux
    port map (
            O => \N__32269\,
            I => \N__32186\
        );

    \I__6811\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32186\
        );

    \I__6810\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32186\
        );

    \I__6809\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32177\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__32263\,
            I => \N__32174\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__32260\,
            I => \N__32167\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__32253\,
            I => \N__32167\
        );

    \I__6805\ : Span4Mux_v
    port map (
            O => \N__32250\,
            I => \N__32167\
        );

    \I__6804\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32164\
        );

    \I__6803\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32160\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__32243\,
            I => \N__32157\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__32234\,
            I => \N__32148\
        );

    \I__6800\ : Span4Mux_v
    port map (
            O => \N__32229\,
            I => \N__32148\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__32226\,
            I => \N__32148\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32148\
        );

    \I__6797\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32143\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32140\
        );

    \I__6795\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32125\
        );

    \I__6794\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32125\
        );

    \I__6793\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32125\
        );

    \I__6792\ : InMux
    port map (
            O => \N__32199\,
            I => \N__32125\
        );

    \I__6791\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32125\
        );

    \I__6790\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32125\
        );

    \I__6789\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32125\
        );

    \I__6788\ : Span4Mux_v
    port map (
            O => \N__32193\,
            I => \N__32120\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__32186\,
            I => \N__32120\
        );

    \I__6786\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32107\
        );

    \I__6785\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32107\
        );

    \I__6784\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32107\
        );

    \I__6783\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32107\
        );

    \I__6782\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32107\
        );

    \I__6781\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32107\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32104\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__32174\,
            I => \N__32097\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__32167\,
            I => \N__32097\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32097\
        );

    \I__6776\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32094\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__32160\,
            I => \N__32087\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__32157\,
            I => \N__32087\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__32148\,
            I => \N__32087\
        );

    \I__6772\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32082\
        );

    \I__6771\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32082\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32073\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__32140\,
            I => \N__32073\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32073\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__32120\,
            I => \N__32073\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__32107\,
            I => \N__32070\
        );

    \I__6765\ : Odrv12
    port map (
            O => \N__32104\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6764\ : Odrv4
    port map (
            O => \N__32097\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__32094\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__32087\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__32082\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6760\ : Odrv4
    port map (
            O => \N__32073\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6759\ : Odrv12
    port map (
            O => \N__32070\,
            I => \b2v_inst11.N_2904_i\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__32055\,
            I => \N__32052\
        );

    \I__6757\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32049\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__6755\ : Span12Mux_s1_h
    port map (
            O => \N__32046\,
            I => \N__32043\
        );

    \I__6754\ : Odrv12
    port map (
            O => \N__32043\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_12\
        );

    \I__6753\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__32037\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_7\
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__32034\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\
        );

    \I__6750\ : CascadeMux
    port map (
            O => \N__32031\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_9_cascade_\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__6748\ : InMux
    port map (
            O => \N__32025\,
            I => \N__32022\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__32022\,
            I => \N__32019\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__32016\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_10\
        );

    \I__6744\ : InMux
    port map (
            O => \N__32013\,
            I => \N__32010\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__6741\ : Odrv4
    port map (
            O => \N__32004\,
            I => \b2v_inst11.un1_dutycycle_94_s1_9\
        );

    \I__6740\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31998\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31995\
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__31995\,
            I => \b2v_inst11.un1_dutycycle_94_s0_9\
        );

    \I__6737\ : CascadeMux
    port map (
            O => \N__31992\,
            I => \b2v_inst11.i2_mux_cascade_\
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__31989\,
            I => \N__31980\
        );

    \I__6735\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31977\
        );

    \I__6734\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31974\
        );

    \I__6733\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31971\
        );

    \I__6732\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31966\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__31984\,
            I => \N__31962\
        );

    \I__6730\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31958\
        );

    \I__6729\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31955\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__31977\,
            I => \N__31952\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__31974\,
            I => \N__31949\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__31971\,
            I => \N__31945\
        );

    \I__6725\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31942\
        );

    \I__6724\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31939\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__31966\,
            I => \N__31936\
        );

    \I__6722\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31929\
        );

    \I__6721\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31929\
        );

    \I__6720\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31929\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__31958\,
            I => \N__31926\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__31955\,
            I => \N__31923\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__31952\,
            I => \N__31920\
        );

    \I__6716\ : Span4Mux_h
    port map (
            O => \N__31949\,
            I => \N__31917\
        );

    \I__6715\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31914\
        );

    \I__6714\ : Span4Mux_s3_h
    port map (
            O => \N__31945\,
            I => \N__31903\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__31942\,
            I => \N__31903\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__31939\,
            I => \N__31903\
        );

    \I__6711\ : Span4Mux_s1_v
    port map (
            O => \N__31936\,
            I => \N__31903\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31903\
        );

    \I__6709\ : Span4Mux_s2_h
    port map (
            O => \N__31926\,
            I => \N__31898\
        );

    \I__6708\ : Span4Mux_s2_h
    port map (
            O => \N__31923\,
            I => \N__31898\
        );

    \I__6707\ : Odrv4
    port map (
            O => \N__31920\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__6706\ : Odrv4
    port map (
            O => \N__31917\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__31914\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__6704\ : Odrv4
    port map (
            O => \N__31903\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__31898\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__6702\ : CascadeMux
    port map (
            O => \N__31887\,
            I => \b2v_inst11.un1_N_5_cascade_\
        );

    \I__6701\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31880\
        );

    \I__6700\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31877\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__31880\,
            I => \b2v_inst11.un1_i2_mux_0_0\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__31877\,
            I => \b2v_inst11.un1_i2_mux_0_0\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__31872\,
            I => \N__31869\
        );

    \I__6696\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31866\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31863\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__31863\,
            I => \N__31860\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__31860\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_11\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__31857\,
            I => \N__31854\
        );

    \I__6691\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31851\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__31851\,
            I => \N__31848\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__31848\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_14\
        );

    \I__6688\ : InMux
    port map (
            O => \N__31845\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_s0\
        );

    \I__6687\ : InMux
    port map (
            O => \N__31842\,
            I => \N__31839\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__31839\,
            I => \N__31836\
        );

    \I__6685\ : Span4Mux_s3_v
    port map (
            O => \N__31836\,
            I => \N__31833\
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__31833\,
            I => \b2v_inst11.un1_dutycycle_94_axb_15_s0\
        );

    \I__6683\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31827\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__31827\,
            I => \N__31824\
        );

    \I__6681\ : Odrv12
    port map (
            O => \N__31824\,
            I => \b2v_inst11.un1_dutycycle_94_s1_15\
        );

    \I__6680\ : InMux
    port map (
            O => \N__31821\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14_s0\
        );

    \I__6679\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31815\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__31815\,
            I => \N__31812\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__31812\,
            I => \b2v_inst11.un1_dutycycle_53_axb_12_1\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__31809\,
            I => \N__31806\
        );

    \I__6675\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31803\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31800\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__31800\,
            I => \b2v_inst11.un1_dutycycle_53_3_1\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__31797\,
            I => \b2v_inst11.un1_dutycycle_53_31_cascade_\
        );

    \I__6671\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__31788\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_13\
        );

    \I__6668\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31782\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__31782\,
            I => \b2v_inst11.un1_dutycycle_53_31\
        );

    \I__6666\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31773\
        );

    \I__6665\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31773\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__6663\ : Span12Mux_s3_h
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__6662\ : Odrv12
    port map (
            O => \N__31767\,
            I => \b2v_inst11.un1_dutycycle_53_55_0_tz\
        );

    \I__6661\ : CascadeMux
    port map (
            O => \N__31764\,
            I => \b2v_inst11.un1_dutycycle_53_axb_14_1_cascade_\
        );

    \I__6660\ : CascadeMux
    port map (
            O => \N__31761\,
            I => \b2v_inst11.un1_dutycycle_53_axb_14_cascade_\
        );

    \I__6659\ : CascadeMux
    port map (
            O => \N__31758\,
            I => \N__31755\
        );

    \I__6658\ : InMux
    port map (
            O => \N__31755\,
            I => \N__31752\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__31752\,
            I => \N__31749\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__31749\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_14\
        );

    \I__6655\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__31737\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_9\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__6650\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__6648\ : Odrv4
    port map (
            O => \N__31725\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_6\
        );

    \I__6647\ : InMux
    port map (
            O => \N__31722\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_s0\
        );

    \I__6646\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__31716\,
            I => \b2v_inst11.dutycycle_RNI_10Z0Z_7\
        );

    \I__6644\ : InMux
    port map (
            O => \N__31713\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_s0\
        );

    \I__6643\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__31707\,
            I => \N__31704\
        );

    \I__6641\ : Span4Mux_h
    port map (
            O => \N__31704\,
            I => \N__31701\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__31701\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_8\
        );

    \I__6639\ : InMux
    port map (
            O => \N__31698\,
            I => \bfn_11_14_0_\
        );

    \I__6638\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__31692\,
            I => \N__31689\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__31689\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_9\
        );

    \I__6635\ : InMux
    port map (
            O => \N__31686\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_s0\
        );

    \I__6634\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__6632\ : Odrv12
    port map (
            O => \N__31677\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_10\
        );

    \I__6631\ : InMux
    port map (
            O => \N__31674\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_s0\
        );

    \I__6630\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31668\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31665\
        );

    \I__6628\ : Span4Mux_s1_h
    port map (
            O => \N__31665\,
            I => \N__31662\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__31662\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_11\
        );

    \I__6626\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31656\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N__31653\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__31653\,
            I => \b2v_inst11.un1_dutycycle_94_s0_11\
        );

    \I__6623\ : InMux
    port map (
            O => \N__31650\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10_s0\
        );

    \I__6622\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31644\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__31644\,
            I => \N__31641\
        );

    \I__6620\ : Odrv4
    port map (
            O => \N__31641\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_12\
        );

    \I__6619\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__31635\,
            I => \N__31632\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__31632\,
            I => \b2v_inst11.un1_dutycycle_94_s0_12\
        );

    \I__6616\ : InMux
    port map (
            O => \N__31629\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11_s0\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__31626\,
            I => \N__31623\
        );

    \I__6614\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31617\
        );

    \I__6612\ : Span4Mux_s1_h
    port map (
            O => \N__31617\,
            I => \N__31614\
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__31614\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_13\
        );

    \I__6610\ : InMux
    port map (
            O => \N__31611\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_s0\
        );

    \I__6609\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31605\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31602\
        );

    \I__6607\ : Odrv4
    port map (
            O => \N__31602\,
            I => \b2v_inst11.un1_dutycycle_94_s1_11\
        );

    \I__6606\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31593\
        );

    \I__6605\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31593\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__31593\,
            I => \N__31590\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__31590\,
            I => \N__31587\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__31587\,
            I => \b2v_inst11.dutycycle_rst_6\
        );

    \I__6601\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31578\
        );

    \I__6600\ : CascadeMux
    port map (
            O => \N__31583\,
            I => \N__31574\
        );

    \I__6599\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31571\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__31581\,
            I => \N__31567\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__31578\,
            I => \N__31564\
        );

    \I__6596\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31559\
        );

    \I__6595\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31559\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31549\
        );

    \I__6593\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31544\
        );

    \I__6592\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31544\
        );

    \I__6591\ : Span4Mux_s2_h
    port map (
            O => \N__31564\,
            I => \N__31541\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__31559\,
            I => \N__31538\
        );

    \I__6589\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31535\
        );

    \I__6588\ : CascadeMux
    port map (
            O => \N__31557\,
            I => \N__31529\
        );

    \I__6587\ : CascadeMux
    port map (
            O => \N__31556\,
            I => \N__31524\
        );

    \I__6586\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31515\
        );

    \I__6585\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31515\
        );

    \I__6584\ : InMux
    port map (
            O => \N__31553\,
            I => \N__31515\
        );

    \I__6583\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31515\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__31549\,
            I => \N__31512\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31509\
        );

    \I__6580\ : Span4Mux_v
    port map (
            O => \N__31541\,
            I => \N__31506\
        );

    \I__6579\ : Span12Mux_s7_v
    port map (
            O => \N__31538\,
            I => \N__31501\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__31535\,
            I => \N__31501\
        );

    \I__6577\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31494\
        );

    \I__6576\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31494\
        );

    \I__6575\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31494\
        );

    \I__6574\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31489\
        );

    \I__6573\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31489\
        );

    \I__6572\ : InMux
    port map (
            O => \N__31527\,
            I => \N__31484\
        );

    \I__6571\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31484\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__31515\,
            I => \N__31477\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__31512\,
            I => \N__31477\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__31509\,
            I => \N__31477\
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__31506\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6566\ : Odrv12
    port map (
            O => \N__31501\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__31494\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__31489\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__31484\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__31477\,
            I => \b2v_inst11.dutycycle\
        );

    \I__6561\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31457\
        );

    \I__6560\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31450\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__31462\,
            I => \N__31445\
        );

    \I__6558\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31435\
        );

    \I__6557\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31435\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__31457\,
            I => \N__31432\
        );

    \I__6555\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31429\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__31455\,
            I => \N__31426\
        );

    \I__6553\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31418\
        );

    \I__6552\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31418\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__31450\,
            I => \N__31415\
        );

    \I__6550\ : InMux
    port map (
            O => \N__31449\,
            I => \N__31406\
        );

    \I__6549\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31406\
        );

    \I__6548\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31406\
        );

    \I__6547\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31406\
        );

    \I__6546\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31399\
        );

    \I__6545\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31399\
        );

    \I__6544\ : InMux
    port map (
            O => \N__31441\,
            I => \N__31399\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31396\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__31435\,
            I => \N__31390\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__31432\,
            I => \N__31385\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31385\
        );

    \I__6539\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31382\
        );

    \I__6538\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31375\
        );

    \I__6537\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31375\
        );

    \I__6536\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31375\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__31418\,
            I => \N__31366\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__31415\,
            I => \N__31366\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__31406\,
            I => \N__31366\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__31399\,
            I => \N__31366\
        );

    \I__6531\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31363\
        );

    \I__6530\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31360\
        );

    \I__6529\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31355\
        );

    \I__6528\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31355\
        );

    \I__6527\ : Span4Mux_h
    port map (
            O => \N__31390\,
            I => \N__31352\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__31385\,
            I => \N__31341\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__31382\,
            I => \N__31341\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31341\
        );

    \I__6523\ : Span4Mux_v
    port map (
            O => \N__31366\,
            I => \N__31341\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__31363\,
            I => \N__31341\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__31360\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__31355\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__6519\ : Odrv4
    port map (
            O => \N__31352\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__31341\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__31332\,
            I => \N__31329\
        );

    \I__6516\ : InMux
    port map (
            O => \N__31329\,
            I => \N__31326\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__6514\ : Odrv12
    port map (
            O => \N__31323\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_1\
        );

    \I__6513\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__31317\,
            I => \N__31314\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__31311\,
            I => \N__31308\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__31308\,
            I => \b2v_inst11.un1_dutycycle_94_s0_1\
        );

    \I__6508\ : InMux
    port map (
            O => \N__31305\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_s0\
        );

    \I__6507\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31292\
        );

    \I__6506\ : CascadeMux
    port map (
            O => \N__31301\,
            I => \N__31286\
        );

    \I__6505\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31283\
        );

    \I__6504\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31280\
        );

    \I__6503\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31277\
        );

    \I__6502\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31274\
        );

    \I__6501\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31271\
        );

    \I__6500\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31268\
        );

    \I__6499\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31265\
        );

    \I__6498\ : CascadeMux
    port map (
            O => \N__31291\,
            I => \N__31262\
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__31290\,
            I => \N__31259\
        );

    \I__6496\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31252\
        );

    \I__6495\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31252\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__31283\,
            I => \N__31249\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__31280\,
            I => \N__31246\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31243\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__31274\,
            I => \N__31236\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__31271\,
            I => \N__31236\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__31268\,
            I => \N__31236\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__31265\,
            I => \N__31233\
        );

    \I__6487\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31230\
        );

    \I__6486\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31227\
        );

    \I__6485\ : InMux
    port map (
            O => \N__31258\,
            I => \N__31222\
        );

    \I__6484\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31222\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31219\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__31249\,
            I => \N__31210\
        );

    \I__6481\ : Span4Mux_v
    port map (
            O => \N__31246\,
            I => \N__31210\
        );

    \I__6480\ : Span4Mux_v
    port map (
            O => \N__31243\,
            I => \N__31210\
        );

    \I__6479\ : Span4Mux_v
    port map (
            O => \N__31236\,
            I => \N__31210\
        );

    \I__6478\ : Span4Mux_h
    port map (
            O => \N__31233\,
            I => \N__31207\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__31230\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__31227\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__31222\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__6474\ : Odrv4
    port map (
            O => \N__31219\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__31210\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__31207\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__31194\,
            I => \N__31191\
        );

    \I__6470\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31185\
        );

    \I__6468\ : Span4Mux_s2_h
    port map (
            O => \N__31185\,
            I => \N__31182\
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__31182\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_2\
        );

    \I__6466\ : InMux
    port map (
            O => \N__31179\,
            I => \N__31176\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__31176\,
            I => \N__31173\
        );

    \I__6464\ : Span4Mux_v
    port map (
            O => \N__31173\,
            I => \N__31170\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__6462\ : Odrv4
    port map (
            O => \N__31167\,
            I => \b2v_inst11.un1_dutycycle_94_s0_2\
        );

    \I__6461\ : InMux
    port map (
            O => \N__31164\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_s0\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__6459\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31155\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__31155\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_3\
        );

    \I__6457\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__31149\,
            I => \N__31146\
        );

    \I__6455\ : Odrv4
    port map (
            O => \N__31146\,
            I => \b2v_inst11.un1_dutycycle_94_s0_3\
        );

    \I__6454\ : InMux
    port map (
            O => \N__31143\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2_s0\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__6452\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__6450\ : Odrv12
    port map (
            O => \N__31131\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_4\
        );

    \I__6449\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__31125\,
            I => \N__31122\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__31122\,
            I => \N__31119\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__31119\,
            I => \b2v_inst11.un1_dutycycle_94_s0_4\
        );

    \I__6445\ : InMux
    port map (
            O => \N__31116\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3_s0\
        );

    \I__6444\ : InMux
    port map (
            O => \N__31113\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4_s0\
        );

    \I__6443\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31107\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__31107\,
            I => \N__31104\
        );

    \I__6441\ : Odrv4
    port map (
            O => \N__31104\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_3\
        );

    \I__6440\ : CascadeMux
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__6439\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31092\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__31092\,
            I => \b2v_inst11.un1_dutycycle_94_s1_12\
        );

    \I__6436\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31085\
        );

    \I__6435\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31082\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31077\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31077\
        );

    \I__6432\ : Odrv4
    port map (
            O => \N__31077\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EGZ0Z1\
        );

    \I__6431\ : InMux
    port map (
            O => \N__31074\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10_s1\
        );

    \I__6430\ : InMux
    port map (
            O => \N__31071\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11_s1\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__6428\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31062\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31059\
        );

    \I__6426\ : Span4Mux_s3_h
    port map (
            O => \N__31059\,
            I => \N__31056\
        );

    \I__6425\ : Odrv4
    port map (
            O => \N__31056\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_13\
        );

    \I__6424\ : InMux
    port map (
            O => \N__31053\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_s1\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__6422\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__6420\ : Span4Mux_s2_h
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__31038\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_14\
        );

    \I__6418\ : InMux
    port map (
            O => \N__31035\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_s1\
        );

    \I__6417\ : InMux
    port map (
            O => \N__31032\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14_s1\
        );

    \I__6416\ : CascadeMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__6415\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__31020\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_6\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__6411\ : InMux
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__31008\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_11\
        );

    \I__6408\ : InMux
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__31002\,
            I => \N__30999\
        );

    \I__6406\ : Odrv12
    port map (
            O => \N__30999\,
            I => \b2v_inst11.un1_dutycycle_94_s1_3\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__30996\,
            I => \N__30993\
        );

    \I__6404\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__30990\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_8\
        );

    \I__6402\ : InMux
    port map (
            O => \N__30987\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_s1\
        );

    \I__6401\ : InMux
    port map (
            O => \N__30984\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2_s1\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__30981\,
            I => \N__30978\
        );

    \I__6399\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__30972\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_4\
        );

    \I__6396\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__30963\,
            I => \N__30960\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__30960\,
            I => \N__30957\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__30957\,
            I => \b2v_inst11.un1_dutycycle_94_s1_4\
        );

    \I__6391\ : InMux
    port map (
            O => \N__30954\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3_s1\
        );

    \I__6390\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__30948\,
            I => \N__30942\
        );

    \I__6388\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30939\
        );

    \I__6387\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30936\
        );

    \I__6386\ : IoInMux
    port map (
            O => \N__30945\,
            I => \N__30933\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__30942\,
            I => \N__30930\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30925\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__30936\,
            I => \N__30925\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30922\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__30930\,
            I => \N__30917\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__30925\,
            I => \N__30917\
        );

    \I__6379\ : Span4Mux_s1_h
    port map (
            O => \N__30922\,
            I => \N__30914\
        );

    \I__6378\ : Sp12to4
    port map (
            O => \N__30917\,
            I => \N__30911\
        );

    \I__6377\ : Span4Mux_v
    port map (
            O => \N__30914\,
            I => \N__30908\
        );

    \I__6376\ : Odrv12
    port map (
            O => \N__30911\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__30908\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6374\ : InMux
    port map (
            O => \N__30903\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4_s1\
        );

    \I__6373\ : InMux
    port map (
            O => \N__30900\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_s1\
        );

    \I__6372\ : CascadeMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__6371\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30891\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__6369\ : Span4Mux_s2_h
    port map (
            O => \N__30888\,
            I => \N__30885\
        );

    \I__6368\ : Odrv4
    port map (
            O => \N__30885\,
            I => \b2v_inst11.dutycycle_RNI_9Z0Z_7\
        );

    \I__6367\ : InMux
    port map (
            O => \N__30882\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_s1\
        );

    \I__6366\ : InMux
    port map (
            O => \N__30879\,
            I => \bfn_11_10_0_\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__30876\,
            I => \N__30873\
        );

    \I__6364\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30867\
        );

    \I__6362\ : Odrv12
    port map (
            O => \N__30867\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_9\
        );

    \I__6361\ : InMux
    port map (
            O => \N__30864\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_s1\
        );

    \I__6360\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30855\
        );

    \I__6358\ : Odrv12
    port map (
            O => \N__30855\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_10\
        );

    \I__6357\ : InMux
    port map (
            O => \N__30852\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_s1\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \b2v_inst11.count_clk_en_cascade_\
        );

    \I__6355\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30842\
        );

    \I__6354\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30839\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__30842\,
            I => \N__30836\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__30839\,
            I => \N__30833\
        );

    \I__6351\ : Odrv12
    port map (
            O => \N__30836\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__6350\ : Odrv4
    port map (
            O => \N__30833\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__6349\ : CascadeMux
    port map (
            O => \N__30828\,
            I => \N__30825\
        );

    \I__6348\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30821\
        );

    \I__6347\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30818\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__30821\,
            I => \N__30815\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__30818\,
            I => \N__30812\
        );

    \I__6344\ : Span4Mux_s3_h
    port map (
            O => \N__30815\,
            I => \N__30809\
        );

    \I__6343\ : Span4Mux_v
    port map (
            O => \N__30812\,
            I => \N__30806\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__30809\,
            I => \b2v_inst11.N_417\
        );

    \I__6341\ : Odrv4
    port map (
            O => \N__30806\,
            I => \b2v_inst11.N_417\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__30801\,
            I => \N__30796\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__30800\,
            I => \N__30793\
        );

    \I__6338\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30783\
        );

    \I__6337\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30783\
        );

    \I__6336\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30783\
        );

    \I__6335\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30783\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__30783\,
            I => \N__30779\
        );

    \I__6333\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__6332\ : Odrv12
    port map (
            O => \N__30779\,
            I => \b2v_inst11.func_state_RNID7Q51Z0Z_0\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__30776\,
            I => \b2v_inst11.func_state_RNID7Q51Z0Z_0\
        );

    \I__6330\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30762\
        );

    \I__6329\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30762\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__30769\,
            I => \N__30758\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30755\
        );

    \I__6326\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30750\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__30762\,
            I => \N__30744\
        );

    \I__6324\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30741\
        );

    \I__6323\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30732\
        );

    \I__6322\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30732\
        );

    \I__6321\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30732\
        );

    \I__6320\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30732\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__30750\,
            I => \N__30729\
        );

    \I__6318\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30722\
        );

    \I__6317\ : InMux
    port map (
            O => \N__30748\,
            I => \N__30722\
        );

    \I__6316\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30722\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__30744\,
            I => \N__30719\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__30741\,
            I => \N__30714\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__30732\,
            I => \N__30714\
        );

    \I__6312\ : Odrv12
    port map (
            O => \N__30729\,
            I => \b2v_inst11.count_off_RNI_1Z0Z_1\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__30722\,
            I => \b2v_inst11.count_off_RNI_1Z0Z_1\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__30719\,
            I => \b2v_inst11.count_off_RNI_1Z0Z_1\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__30714\,
            I => \b2v_inst11.count_off_RNI_1Z0Z_1\
        );

    \I__6308\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__30702\,
            I => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0\
        );

    \I__6306\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30693\
        );

    \I__6305\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30693\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__30693\,
            I => \N__30690\
        );

    \I__6303\ : Odrv12
    port map (
            O => \N__30690\,
            I => \b2v_inst11.func_state_RNI6M5R2Z0Z_1\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__30687\,
            I => \N__30684\
        );

    \I__6301\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30672\
        );

    \I__6300\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30672\
        );

    \I__6299\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30672\
        );

    \I__6298\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30672\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30669\
        );

    \I__6296\ : Span4Mux_s1_h
    port map (
            O => \N__30669\,
            I => \N__30666\
        );

    \I__6295\ : Odrv4
    port map (
            O => \N__30666\,
            I => \b2v_inst11.func_state_RNIJGA54Z0Z_1\
        );

    \I__6294\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30657\
        );

    \I__6293\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30657\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__30657\,
            I => \N__30654\
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__30654\,
            I => \b2v_inst11.count_clk_1_14\
        );

    \I__6290\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30648\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__30648\,
            I => \b2v_inst11.count_clk_0_14\
        );

    \I__6288\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30638\
        );

    \I__6287\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30638\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__30643\,
            I => \N__30630\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__30638\,
            I => \N__30624\
        );

    \I__6284\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30621\
        );

    \I__6283\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30616\
        );

    \I__6282\ : InMux
    port map (
            O => \N__30635\,
            I => \N__30616\
        );

    \I__6281\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30613\
        );

    \I__6280\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30610\
        );

    \I__6279\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30605\
        );

    \I__6278\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30605\
        );

    \I__6277\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30600\
        );

    \I__6276\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30600\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__30624\,
            I => \N__30595\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__30621\,
            I => \N__30595\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__30616\,
            I => \N__30592\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__30613\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__30610\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__30605\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__30600\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__30595\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__30592\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__30579\,
            I => \b2v_inst11.N_2904_i_cascade_\
        );

    \I__6265\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30573\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__6263\ : Span4Mux_v
    port map (
            O => \N__30570\,
            I => \N__30567\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__30567\,
            I => \N__30564\
        );

    \I__6261\ : Odrv4
    port map (
            O => \N__30564\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_1\
        );

    \I__6260\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30558\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__30558\,
            I => \N__30555\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__30555\,
            I => \b2v_inst11.un1_dutycycle_94_s1_1\
        );

    \I__6257\ : InMux
    port map (
            O => \N__30552\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_s1\
        );

    \I__6256\ : CascadeMux
    port map (
            O => \N__30549\,
            I => \N__30546\
        );

    \I__6255\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30543\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__6253\ : Span4Mux_s2_h
    port map (
            O => \N__30540\,
            I => \N__30537\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__30537\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_2\
        );

    \I__6251\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30531\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__30531\,
            I => \N__30528\
        );

    \I__6249\ : Span4Mux_h
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__30525\,
            I => \b2v_inst11.un1_dutycycle_94_s1_2\
        );

    \I__6247\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30515\
        );

    \I__6246\ : InMux
    port map (
            O => \N__30521\,
            I => \N__30515\
        );

    \I__6245\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30512\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__30515\,
            I => \N__30509\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__30512\,
            I => \N__30506\
        );

    \I__6242\ : Span4Mux_v
    port map (
            O => \N__30509\,
            I => \N__30503\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__30506\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__30503\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__6239\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30492\
        );

    \I__6238\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30492\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__30489\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\
        );

    \I__6235\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__30483\,
            I => \b2v_inst11.count_clk_0_8\
        );

    \I__6233\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30471\
        );

    \I__6232\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30471\
        );

    \I__6231\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30471\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__30471\,
            I => \N__30467\
        );

    \I__6229\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30464\
        );

    \I__6228\ : Span4Mux_h
    port map (
            O => \N__30467\,
            I => \N__30461\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__30464\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__30461\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__6225\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30450\
        );

    \I__6224\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30450\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__30450\,
            I => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\
        );

    \I__6222\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30444\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__30444\,
            I => \b2v_inst11.count_clk_0_9\
        );

    \I__6220\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30431\
        );

    \I__6219\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30431\
        );

    \I__6218\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30425\
        );

    \I__6217\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30422\
        );

    \I__6216\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30417\
        );

    \I__6215\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30417\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__30431\,
            I => \N__30414\
        );

    \I__6213\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30411\
        );

    \I__6212\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30406\
        );

    \I__6211\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30406\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__30425\,
            I => \N__30403\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__30422\,
            I => \N__30392\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__30417\,
            I => \N__30392\
        );

    \I__6207\ : Span4Mux_v
    port map (
            O => \N__30414\,
            I => \N__30392\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30392\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30392\
        );

    \I__6204\ : Span4Mux_v
    port map (
            O => \N__30403\,
            I => \N__30389\
        );

    \I__6203\ : Span4Mux_v
    port map (
            O => \N__30392\,
            I => \N__30386\
        );

    \I__6202\ : Odrv4
    port map (
            O => \N__30389\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__6201\ : Odrv4
    port map (
            O => \N__30386\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__30381\,
            I => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0_cascade_\
        );

    \I__6199\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30374\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__30377\,
            I => \N__30371\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30367\
        );

    \I__6196\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30364\
        );

    \I__6195\ : InMux
    port map (
            O => \N__30370\,
            I => \N__30361\
        );

    \I__6194\ : Span4Mux_s2_h
    port map (
            O => \N__30367\,
            I => \N__30358\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__30364\,
            I => \b2v_inst11.N_369\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__30361\,
            I => \b2v_inst11.N_369\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__30358\,
            I => \b2v_inst11.N_369\
        );

    \I__6190\ : InMux
    port map (
            O => \N__30351\,
            I => \bfn_11_6_0_\
        );

    \I__6189\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__30342\,
            I => \b2v_inst11.un1_count_clk_2_axb_10\
        );

    \I__6186\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30330\
        );

    \I__6185\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30330\
        );

    \I__6184\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30330\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__30330\,
            I => \N__30327\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__30327\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\
        );

    \I__6181\ : InMux
    port map (
            O => \N__30324\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\
        );

    \I__6180\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__6178\ : Span4Mux_s3_h
    port map (
            O => \N__30315\,
            I => \N__30312\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__30312\,
            I => \b2v_inst11.un1_count_clk_2_axb_11\
        );

    \I__6176\ : InMux
    port map (
            O => \N__30309\,
            I => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\
        );

    \I__6175\ : InMux
    port map (
            O => \N__30306\,
            I => \b2v_inst11.un1_count_clk_2_cry_11\
        );

    \I__6174\ : InMux
    port map (
            O => \N__30303\,
            I => \b2v_inst11.un1_count_clk_2_cry_12\
        );

    \I__6173\ : InMux
    port map (
            O => \N__30300\,
            I => \b2v_inst11.un1_count_clk_2_cry_13\
        );

    \I__6172\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30291\
        );

    \I__6171\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30291\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__30291\,
            I => \N__30276\
        );

    \I__6169\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30267\
        );

    \I__6168\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30267\
        );

    \I__6167\ : InMux
    port map (
            O => \N__30288\,
            I => \N__30267\
        );

    \I__6166\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30267\
        );

    \I__6165\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30255\
        );

    \I__6164\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30255\
        );

    \I__6163\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30255\
        );

    \I__6162\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30255\
        );

    \I__6161\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30243\
        );

    \I__6160\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30243\
        );

    \I__6159\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30243\
        );

    \I__6158\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30243\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__30276\,
            I => \N__30240\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30237\
        );

    \I__6155\ : InMux
    port map (
            O => \N__30266\,
            I => \N__30230\
        );

    \I__6154\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30230\
        );

    \I__6153\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30230\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__30255\,
            I => \N__30227\
        );

    \I__6151\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30220\
        );

    \I__6150\ : InMux
    port map (
            O => \N__30253\,
            I => \N__30220\
        );

    \I__6149\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30220\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__30243\,
            I => \N__30211\
        );

    \I__6147\ : Span4Mux_s0_h
    port map (
            O => \N__30240\,
            I => \N__30211\
        );

    \I__6146\ : Span4Mux_v
    port map (
            O => \N__30237\,
            I => \N__30211\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__30230\,
            I => \N__30211\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__30227\,
            I => \b2v_inst11.func_state_RNIIGCET1_0_1\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__30220\,
            I => \b2v_inst11.func_state_RNIIGCET1_0_1\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__30211\,
            I => \b2v_inst11.func_state_RNIIGCET1_0_1\
        );

    \I__6141\ : InMux
    port map (
            O => \N__30204\,
            I => \b2v_inst11.un1_count_clk_2_cry_14\
        );

    \I__6140\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30196\
        );

    \I__6139\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30193\
        );

    \I__6138\ : InMux
    port map (
            O => \N__30199\,
            I => \N__30190\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__30196\,
            I => \N__30187\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30184\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__30190\,
            I => \N__30179\
        );

    \I__6134\ : Span4Mux_v
    port map (
            O => \N__30187\,
            I => \N__30179\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__30184\,
            I => \b2v_inst11.count_clk_1_11\
        );

    \I__6132\ : Odrv4
    port map (
            O => \N__30179\,
            I => \b2v_inst11.count_clk_1_11\
        );

    \I__6131\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30170\
        );

    \I__6130\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30167\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__30170\,
            I => \N__30164\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__30167\,
            I => \N__30161\
        );

    \I__6127\ : Span4Mux_h
    port map (
            O => \N__30164\,
            I => \N__30158\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__30161\,
            I => \b2v_inst11.count_clk_0_11\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__30158\,
            I => \b2v_inst11.count_clk_0_11\
        );

    \I__6124\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30143\
        );

    \I__6123\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30143\
        );

    \I__6122\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30143\
        );

    \I__6121\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30140\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__30143\,
            I => \N__30137\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30134\
        );

    \I__6118\ : Span4Mux_h
    port map (
            O => \N__30137\,
            I => \N__30129\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__30134\,
            I => \N__30129\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__30129\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__6115\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30120\
        );

    \I__6114\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30120\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__30120\,
            I => \b2v_inst11.count_clk_0_10\
        );

    \I__6112\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30110\
        );

    \I__6110\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30107\
        );

    \I__6109\ : Span4Mux_s2_h
    port map (
            O => \N__30110\,
            I => \N__30104\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__30107\,
            I => \b2v_inst11.un1_count_clk_2_axb_1\
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__30104\,
            I => \b2v_inst11.un1_count_clk_2_axb_1\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__30099\,
            I => \N__30096\
        );

    \I__6105\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30091\
        );

    \I__6104\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30088\
        );

    \I__6103\ : CascadeMux
    port map (
            O => \N__30094\,
            I => \N__30085\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30080\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__30088\,
            I => \N__30077\
        );

    \I__6100\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30070\
        );

    \I__6099\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30070\
        );

    \I__6098\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30070\
        );

    \I__6097\ : Span4Mux_s2_h
    port map (
            O => \N__30080\,
            I => \N__30067\
        );

    \I__6096\ : Odrv12
    port map (
            O => \N__30077\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__30070\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__30067\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__6093\ : InMux
    port map (
            O => \N__30060\,
            I => \b2v_inst11.un1_count_clk_2_cry_1\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__30057\,
            I => \N__30054\
        );

    \I__6091\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30051\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__30051\,
            I => \N__30048\
        );

    \I__6089\ : Odrv12
    port map (
            O => \N__30048\,
            I => \b2v_inst11.un1_count_clk_2_axb_3\
        );

    \I__6088\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30036\
        );

    \I__6087\ : InMux
    port map (
            O => \N__30044\,
            I => \N__30036\
        );

    \I__6086\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30036\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__30036\,
            I => \N__30033\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__30033\,
            I => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\
        );

    \I__6083\ : InMux
    port map (
            O => \N__30030\,
            I => \b2v_inst11.un1_count_clk_2_cry_2\
        );

    \I__6082\ : InMux
    port map (
            O => \N__30027\,
            I => \b2v_inst11.un1_count_clk_2_cry_3\
        );

    \I__6081\ : InMux
    port map (
            O => \N__30024\,
            I => \b2v_inst11.un1_count_clk_2_cry_4\
        );

    \I__6080\ : InMux
    port map (
            O => \N__30021\,
            I => \b2v_inst11.un1_count_clk_2_cry_5\
        );

    \I__6079\ : InMux
    port map (
            O => \N__30018\,
            I => \b2v_inst11.un1_count_clk_2_cry_6\
        );

    \I__6078\ : InMux
    port map (
            O => \N__30015\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\
        );

    \I__6077\ : InMux
    port map (
            O => \N__30012\,
            I => \b2v_inst6.un2_count_1_cry_14\
        );

    \I__6076\ : InMux
    port map (
            O => \N__30009\,
            I => \N__30006\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__30006\,
            I => \b2v_inst6.un2_count_1_axb_13\
        );

    \I__6074\ : InMux
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__30000\,
            I => \b2v_inst11.count_clkZ0Z_10\
        );

    \I__6072\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29994\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__29994\,
            I => \b2v_inst11.count_clkZ0Z_12\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__29991\,
            I => \b2v_inst11.count_clkZ0Z_13_cascade_\
        );

    \I__6069\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29985\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__29985\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__29982\,
            I => \b2v_inst11.un2_count_clk_17_0_o2_4_cascade_\
        );

    \I__6066\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29967\
        );

    \I__6065\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29967\
        );

    \I__6064\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29967\
        );

    \I__6063\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29967\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__29967\,
            I => \N__29964\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__29964\,
            I => \N__29961\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__29961\,
            I => \b2v_inst11.N_175\
        );

    \I__6059\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29954\
        );

    \I__6058\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29951\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__29954\,
            I => \b2v_inst6.un2_count_1_axb_7\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__29951\,
            I => \b2v_inst6.un2_count_1_axb_7\
        );

    \I__6055\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29940\
        );

    \I__6054\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29940\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__29940\,
            I => \b2v_inst6.un2_count_1_cry_6_THRU_CO\
        );

    \I__6052\ : InMux
    port map (
            O => \N__29937\,
            I => \b2v_inst6.un2_count_1_cry_6\
        );

    \I__6051\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29931\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29927\
        );

    \I__6049\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29924\
        );

    \I__6048\ : Span4Mux_s2_h
    port map (
            O => \N__29927\,
            I => \N__29921\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__29924\,
            I => \b2v_inst6.un2_count_1_axb_8\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__29921\,
            I => \b2v_inst6.un2_count_1_axb_8\
        );

    \I__6045\ : CascadeMux
    port map (
            O => \N__29916\,
            I => \N__29913\
        );

    \I__6044\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29907\
        );

    \I__6043\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29907\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__29907\,
            I => \N__29904\
        );

    \I__6041\ : Span4Mux_s1_v
    port map (
            O => \N__29904\,
            I => \N__29901\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__29901\,
            I => \b2v_inst6.un2_count_1_cry_7_THRU_CO\
        );

    \I__6039\ : InMux
    port map (
            O => \N__29898\,
            I => \b2v_inst6.un2_count_1_cry_7\
        );

    \I__6038\ : InMux
    port map (
            O => \N__29895\,
            I => \N__29891\
        );

    \I__6037\ : InMux
    port map (
            O => \N__29894\,
            I => \N__29888\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__29891\,
            I => \N__29885\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29880\
        );

    \I__6034\ : Span4Mux_v
    port map (
            O => \N__29885\,
            I => \N__29880\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__29880\,
            I => \b2v_inst6.un2_count_1_axb_9\
        );

    \I__6032\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29871\
        );

    \I__6031\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29871\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29868\
        );

    \I__6029\ : Span4Mux_s2_v
    port map (
            O => \N__29868\,
            I => \N__29865\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__29865\,
            I => \b2v_inst6.un2_count_1_cry_8_THRU_CO\
        );

    \I__6027\ : InMux
    port map (
            O => \N__29862\,
            I => \bfn_11_3_0_\
        );

    \I__6026\ : InMux
    port map (
            O => \N__29859\,
            I => \b2v_inst6.un2_count_1_cry_9\
        );

    \I__6025\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29850\
        );

    \I__6024\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29850\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__29850\,
            I => \N__29847\
        );

    \I__6022\ : Odrv4
    port map (
            O => \N__29847\,
            I => \b2v_inst6.un2_count_1_cry_10_THRU_CO\
        );

    \I__6021\ : InMux
    port map (
            O => \N__29844\,
            I => \b2v_inst6.un2_count_1_cry_10\
        );

    \I__6020\ : InMux
    port map (
            O => \N__29841\,
            I => \b2v_inst6.un2_count_1_cry_11\
        );

    \I__6019\ : InMux
    port map (
            O => \N__29838\,
            I => \b2v_inst6.un2_count_1_cry_12\
        );

    \I__6018\ : InMux
    port map (
            O => \N__29835\,
            I => \b2v_inst6.un2_count_1_cry_13\
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__29832\,
            I => \b2v_inst6.count_rst_3_cascade_\
        );

    \I__6016\ : CascadeMux
    port map (
            O => \N__29829\,
            I => \b2v_inst6.countZ0Z_11_cascade_\
        );

    \I__6015\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29823\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__29823\,
            I => \b2v_inst6.count_0_11\
        );

    \I__6013\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29810\
        );

    \I__6012\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29797\
        );

    \I__6011\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29797\
        );

    \I__6010\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29797\
        );

    \I__6009\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29797\
        );

    \I__6008\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29797\
        );

    \I__6007\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29797\
        );

    \I__6006\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29790\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__29810\,
            I => \N__29787\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__29797\,
            I => \N__29784\
        );

    \I__6003\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29770\
        );

    \I__6002\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29770\
        );

    \I__6001\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29770\
        );

    \I__6000\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29770\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__29790\,
            I => \N__29763\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29763\
        );

    \I__5997\ : Span4Mux_s1_v
    port map (
            O => \N__29784\,
            I => \N__29763\
        );

    \I__5996\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29754\
        );

    \I__5995\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29754\
        );

    \I__5994\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29754\
        );

    \I__5993\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29754\
        );

    \I__5992\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29751\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__29770\,
            I => \b2v_inst6.N_394\
        );

    \I__5990\ : Odrv4
    port map (
            O => \N__29763\,
            I => \b2v_inst6.N_394\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__29754\,
            I => \b2v_inst6.N_394\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__29751\,
            I => \b2v_inst6.N_394\
        );

    \I__5987\ : InMux
    port map (
            O => \N__29742\,
            I => \b2v_inst6.un2_count_1_cry_1\
        );

    \I__5986\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29735\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__29735\,
            I => \N__29729\
        );

    \I__5983\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29726\
        );

    \I__5982\ : Span4Mux_s3_h
    port map (
            O => \N__29729\,
            I => \N__29723\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__29726\,
            I => \b2v_inst6.un2_count_1_axb_3\
        );

    \I__5980\ : Odrv4
    port map (
            O => \N__29723\,
            I => \b2v_inst6.un2_count_1_axb_3\
        );

    \I__5979\ : InMux
    port map (
            O => \N__29718\,
            I => \N__29712\
        );

    \I__5978\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29712\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__5976\ : Span4Mux_s1_v
    port map (
            O => \N__29709\,
            I => \N__29706\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__29706\,
            I => \b2v_inst6.un2_count_1_cry_2_THRU_CO\
        );

    \I__5974\ : InMux
    port map (
            O => \N__29703\,
            I => \b2v_inst6.un2_count_1_cry_2\
        );

    \I__5973\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29695\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__29699\,
            I => \N__29692\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__29698\,
            I => \N__29689\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29686\
        );

    \I__5969\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29681\
        );

    \I__5968\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29681\
        );

    \I__5967\ : Span4Mux_v
    port map (
            O => \N__29686\,
            I => \N__29678\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__29681\,
            I => \b2v_inst6.un2_count_1_axb_4\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__29678\,
            I => \b2v_inst6.un2_count_1_axb_4\
        );

    \I__5964\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29667\
        );

    \I__5963\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29667\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__29667\,
            I => \N__29664\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__29664\,
            I => \N__29661\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__29661\,
            I => \b2v_inst6.un2_count_1_cry_3_THRU_CO\
        );

    \I__5959\ : InMux
    port map (
            O => \N__29658\,
            I => \b2v_inst6.un2_count_1_cry_3\
        );

    \I__5958\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29649\
        );

    \I__5957\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29649\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__29649\,
            I => \b2v_inst6.un2_count_1_cry_4_THRU_CO\
        );

    \I__5955\ : InMux
    port map (
            O => \N__29646\,
            I => \b2v_inst6.un2_count_1_cry_4\
        );

    \I__5954\ : InMux
    port map (
            O => \N__29643\,
            I => \b2v_inst6.un2_count_1_cry_5\
        );

    \I__5953\ : CascadeMux
    port map (
            O => \N__29640\,
            I => \b2v_inst11.N_11_cascade_\
        );

    \I__5952\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__29634\,
            I => \b2v_inst11.N_35_0\
        );

    \I__5950\ : CascadeMux
    port map (
            O => \N__29631\,
            I => \b2v_inst11.N_13_cascade_\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__29628\,
            I => \N__29624\
        );

    \I__5948\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29619\
        );

    \I__5947\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29619\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__29619\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_11\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__29616\,
            I => \N__29613\
        );

    \I__5944\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__29610\,
            I => \b2v_inst11.g0_6_a5_1_0\
        );

    \I__5942\ : CascadeMux
    port map (
            O => \N__29607\,
            I => \b2v_inst6.count_rst_7_cascade_\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__29604\,
            I => \b2v_inst6.un2_count_1_axb_7_cascade_\
        );

    \I__5940\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__29598\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_6\
        );

    \I__5938\ : CascadeMux
    port map (
            O => \N__29595\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_\
        );

    \I__5937\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29589\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__29589\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_11\
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__29586\,
            I => \N__29583\
        );

    \I__5934\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29580\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__29580\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_15\
        );

    \I__5932\ : CascadeMux
    port map (
            O => \N__29577\,
            I => \N__29574\
        );

    \I__5931\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29571\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__29571\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_14\
        );

    \I__5929\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29562\
        );

    \I__5928\ : InMux
    port map (
            O => \N__29567\,
            I => \N__29562\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__29562\,
            I => \b2v_inst11.un1_dutycycle_53_44_0_0\
        );

    \I__5926\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29556\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__29556\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_8\
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__29553\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_\
        );

    \I__5923\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__5921\ : Span4Mux_s1_v
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__29541\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_7\
        );

    \I__5919\ : CascadeMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__5918\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29532\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__29532\,
            I => \b2v_inst11.un1_dutycycle_53_axb_10\
        );

    \I__5916\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29522\
        );

    \I__5914\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29519\
        );

    \I__5913\ : Odrv4
    port map (
            O => \N__29522\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_7\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__29519\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_7\
        );

    \I__5911\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29511\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__29511\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_7\
        );

    \I__5909\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29504\
        );

    \I__5908\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29501\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__29504\,
            I => \N__29498\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__29501\,
            I => \b2v_inst11.CO2_THRU_CO\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__29498\,
            I => \b2v_inst11.CO2_THRU_CO\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__5903\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29487\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__5901\ : Odrv4
    port map (
            O => \N__29484\,
            I => \b2v_inst11.mult1_un54_sum_axb_6_i_l_fx\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__5899\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29471\
        );

    \I__5898\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29471\
        );

    \I__5897\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29468\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29465\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__29468\,
            I => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\
        );

    \I__5894\ : Odrv4
    port map (
            O => \N__29465\,
            I => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__5892\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29451\
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__29451\,
            I => \b2v_inst11.mult1_un54_sum_axb_5_i_l_ofx\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__29448\,
            I => \N__29443\
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__29447\,
            I => \N__29438\
        );

    \I__5887\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29435\
        );

    \I__5886\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29432\
        );

    \I__5885\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29425\
        );

    \I__5884\ : InMux
    port map (
            O => \N__29441\,
            I => \N__29425\
        );

    \I__5883\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29425\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__29435\,
            I => \N__29422\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__29432\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__29425\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__29422\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0\
        );

    \I__5878\ : CascadeMux
    port map (
            O => \N__29415\,
            I => \N__29410\
        );

    \I__5877\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29406\
        );

    \I__5876\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29399\
        );

    \I__5875\ : InMux
    port map (
            O => \N__29410\,
            I => \N__29399\
        );

    \I__5874\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29399\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__29406\,
            I => \b2v_inst11.mult1_un40_sum_i_2\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__29399\,
            I => \b2v_inst11.mult1_un40_sum_i_2\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__5870\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29388\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__29388\,
            I => \N__29385\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__29385\,
            I => \b2v_inst11.mult1_un47_sum1_3\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__29382\,
            I => \b2v_inst11.un1_dutycycle_53_axb_12_cascade_\
        );

    \I__5866\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29376\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__29376\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_15\
        );

    \I__5864\ : CascadeMux
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__5863\ : InMux
    port map (
            O => \N__29370\,
            I => \N__29367\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__29367\,
            I => \b2v_inst11.dutycycle_eena_9\
        );

    \I__5861\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29358\
        );

    \I__5860\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29358\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__29358\,
            I => \b2v_inst11.dutycycleZ1Z_12\
        );

    \I__5858\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29349\
        );

    \I__5857\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29349\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__29349\,
            I => \b2v_inst11.dutycycleZ1Z_11\
        );

    \I__5855\ : InMux
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__29343\,
            I => \b2v_inst11.dutycycle_eena_7\
        );

    \I__5853\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__29337\,
            I => \b2v_inst11.N_6_0\
        );

    \I__5851\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \b2v_inst11.N_8_cascade_\
        );

    \I__5850\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__29328\,
            I => \N__29324\
        );

    \I__5848\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29321\
        );

    \I__5847\ : Span4Mux_h
    port map (
            O => \N__29324\,
            I => \N__29318\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__29321\,
            I => \b2v_inst11.N_355\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__29318\,
            I => \b2v_inst11.N_355\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__29313\,
            I => \b2v_inst11.g0_6_a5_0_0_cascade_\
        );

    \I__5843\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__29307\,
            I => \b2v_inst11.g0_6_a5_2_1\
        );

    \I__5841\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29301\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__5839\ : Span4Mux_v
    port map (
            O => \N__29298\,
            I => \N__29294\
        );

    \I__5838\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29291\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__29294\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__29291\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__29286\,
            I => \b2v_inst11.dutycycle_eena_9_cascade_\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__29283\,
            I => \b2v_inst11.dutycycle_eena_7_cascade_\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__29280\,
            I => \N__29272\
        );

    \I__5832\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29263\
        );

    \I__5831\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29263\
        );

    \I__5830\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29263\
        );

    \I__5829\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29263\
        );

    \I__5828\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29258\
        );

    \I__5827\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29258\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29253\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__29258\,
            I => \N__29253\
        );

    \I__5824\ : Span4Mux_h
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__29250\,
            I => \b2v_inst11.N_2943_i\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__5821\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29236\
        );

    \I__5820\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29236\
        );

    \I__5819\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29233\
        );

    \I__5818\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29230\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29225\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29225\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__29230\,
            I => \N__29221\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__29225\,
            I => \N__29218\
        );

    \I__5813\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29215\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__29221\,
            I => \b2v_inst11.func_state_RNIDQ4A1Z0Z_1\
        );

    \I__5811\ : Odrv4
    port map (
            O => \N__29218\,
            I => \b2v_inst11.func_state_RNIDQ4A1Z0Z_1\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__29215\,
            I => \b2v_inst11.func_state_RNIDQ4A1Z0Z_1\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__29208\,
            I => \b2v_inst11.N_360_cascade_\
        );

    \I__5808\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29202\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__29202\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\
        );

    \I__5806\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29193\
        );

    \I__5805\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29193\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__29193\,
            I => \b2v_inst11.N_234_N\
        );

    \I__5803\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29187\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__29187\,
            I => \N__29184\
        );

    \I__5801\ : Span4Mux_h
    port map (
            O => \N__29184\,
            I => \N__29181\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__29181\,
            I => \b2v_inst11.N_309\
        );

    \I__5799\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29175\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__29175\,
            I => \N__29172\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__29172\,
            I => \b2v_inst11.un1_dutycycle_96_0_a3_1\
        );

    \I__5796\ : CascadeMux
    port map (
            O => \N__29169\,
            I => \N__29166\
        );

    \I__5795\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29159\
        );

    \I__5793\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29156\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__29159\,
            I => \b2v_inst11.dutycycle_eena_0\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__29156\,
            I => \b2v_inst11.dutycycle_eena_0\
        );

    \I__5790\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29146\
        );

    \I__5789\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29141\
        );

    \I__5788\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29141\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29138\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29135\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__29138\,
            I => \b2v_inst11.un1_clk_100khz_25_and_i_0_1_0\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__29135\,
            I => \b2v_inst11.un1_clk_100khz_25_and_i_0_1_0\
        );

    \I__5783\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__29127\,
            I => \b2v_inst11.N_186_i\
        );

    \I__5781\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29121\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__29121\,
            I => \b2v_inst11.N_117_f0_1\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29113\
        );

    \I__5778\ : IoInMux
    port map (
            O => \N__29117\,
            I => \N__29109\
        );

    \I__5777\ : IoInMux
    port map (
            O => \N__29116\,
            I => \N__29104\
        );

    \I__5776\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29099\
        );

    \I__5775\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29099\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__29109\,
            I => \N__29096\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__29108\,
            I => \N__29093\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__29107\,
            I => \N__29090\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__29104\,
            I => \N__29084\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__29099\,
            I => \N__29081\
        );

    \I__5769\ : IoSpan4Mux
    port map (
            O => \N__29096\,
            I => \N__29078\
        );

    \I__5768\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29075\
        );

    \I__5767\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29068\
        );

    \I__5766\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29068\
        );

    \I__5765\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29068\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__29087\,
            I => \N__29065\
        );

    \I__5763\ : Span4Mux_s2_h
    port map (
            O => \N__29084\,
            I => \N__29062\
        );

    \I__5762\ : Span4Mux_h
    port map (
            O => \N__29081\,
            I => \N__29059\
        );

    \I__5761\ : Span4Mux_s2_h
    port map (
            O => \N__29078\,
            I => \N__29056\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29051\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29051\
        );

    \I__5758\ : InMux
    port map (
            O => \N__29065\,
            I => \N__29048\
        );

    \I__5757\ : Span4Mux_h
    port map (
            O => \N__29062\,
            I => \N__29043\
        );

    \I__5756\ : Span4Mux_v
    port map (
            O => \N__29059\,
            I => \N__29043\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__29056\,
            I => \N__29038\
        );

    \I__5754\ : Span4Mux_h
    port map (
            O => \N__29051\,
            I => \N__29038\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__29048\,
            I => v5s_enn
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__29043\,
            I => v5s_enn
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__29038\,
            I => v5s_enn
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__29031\,
            I => \b2v_inst11.N_117_f0_1_cascade_\
        );

    \I__5749\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29022\
        );

    \I__5748\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29022\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__29022\,
            I => \b2v_inst11.dutycycle_eena\
        );

    \I__5746\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29013\
        );

    \I__5745\ : InMux
    port map (
            O => \N__29018\,
            I => \N__29013\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__29013\,
            I => \b2v_inst11.dutycycleZ1Z_2\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__29010\,
            I => \N__29006\
        );

    \I__5742\ : InMux
    port map (
            O => \N__29009\,
            I => \N__29003\
        );

    \I__5741\ : InMux
    port map (
            O => \N__29006\,
            I => \N__29000\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__29003\,
            I => \N__28995\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__29000\,
            I => \N__28995\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__28995\,
            I => \N__28992\
        );

    \I__5737\ : Odrv4
    port map (
            O => \N__28992\,
            I => \b2v_inst11.N_73\
        );

    \I__5736\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28983\
        );

    \I__5735\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28983\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__28983\,
            I => \b2v_inst11.dutycycle_eena_1\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28977\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28974\
        );

    \I__5731\ : Span4Mux_h
    port map (
            O => \N__28974\,
            I => \N__28971\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__28971\,
            I => \b2v_inst11.N_159\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__28968\,
            I => \b2v_inst11.dutycycleZ0Z_1_cascade_\
        );

    \I__5728\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28961\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__28964\,
            I => \N__28957\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__28961\,
            I => \N__28953\
        );

    \I__5725\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28946\
        );

    \I__5724\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28946\
        );

    \I__5723\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28946\
        );

    \I__5722\ : Span4Mux_h
    port map (
            O => \N__28953\,
            I => \N__28943\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__28946\,
            I => \b2v_inst11.N_363\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__28943\,
            I => \b2v_inst11.N_363\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__28938\,
            I => \b2v_inst11.dutycycle_1_0_1_cascade_\
        );

    \I__5718\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28929\
        );

    \I__5717\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28929\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__28926\,
            I => \b2v_inst11.dutycycleZ1Z_1\
        );

    \I__5714\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__28920\,
            I => \b2v_inst11.dutycycle_1_0_0\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__5711\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28908\
        );

    \I__5710\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28908\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__28908\,
            I => \b2v_inst11.dutycycleZ1Z_0\
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__28905\,
            I => \b2v_inst11.dutycycle_1_0_0_cascade_\
        );

    \I__5707\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28896\
        );

    \I__5706\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28896\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__28896\,
            I => \b2v_inst11.dutycycle_RNI_8Z0Z_0\
        );

    \I__5704\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28889\
        );

    \I__5703\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28886\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__28889\,
            I => \N__28880\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28880\
        );

    \I__5700\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28877\
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__28880\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_2\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__28877\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_2\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__28872\,
            I => \N__28868\
        );

    \I__5696\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28863\
        );

    \I__5695\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28863\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28855\
        );

    \I__5693\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28852\
        );

    \I__5692\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28849\
        );

    \I__5691\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28842\
        );

    \I__5690\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28842\
        );

    \I__5689\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28842\
        );

    \I__5688\ : Span4Mux_h
    port map (
            O => \N__28855\,
            I => \N__28839\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__28852\,
            I => \b2v_inst11.N_19_i\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__28849\,
            I => \b2v_inst11.N_19_i\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__28842\,
            I => \b2v_inst11.N_19_i\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__28839\,
            I => \b2v_inst11.N_19_i\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__28830\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_0_cascade_\
        );

    \I__5682\ : InMux
    port map (
            O => \N__28827\,
            I => \N__28824\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__28824\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__28821\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__28818\,
            I => \b2v_inst11.N_186_i_cascade_\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__28815\,
            I => \N__28811\
        );

    \I__5677\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28801\
        );

    \I__5676\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28801\
        );

    \I__5675\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28801\
        );

    \I__5674\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28797\
        );

    \I__5673\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28791\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28787\
        );

    \I__5671\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28784\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28781\
        );

    \I__5669\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28774\
        );

    \I__5668\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28774\
        );

    \I__5667\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28774\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__28791\,
            I => \N__28771\
        );

    \I__5665\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28766\
        );

    \I__5664\ : Span4Mux_h
    port map (
            O => \N__28787\,
            I => \N__28763\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28754\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__28781\,
            I => \N__28754\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__28774\,
            I => \N__28754\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__28771\,
            I => \N__28754\
        );

    \I__5659\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28749\
        );

    \I__5658\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28749\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__28766\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__28763\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__28754\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__28749\,
            I => \curr_state_RNID8DP1_0_0\
        );

    \I__5653\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__28737\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0_0\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__28734\,
            I => \N__28730\
        );

    \I__5650\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28725\
        );

    \I__5649\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28725\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__28725\,
            I => \b2v_inst11.N_160_i\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__28722\,
            I => \b2v_inst11.N_160_i_cascade_\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__28719\,
            I => \N__28715\
        );

    \I__5645\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28711\
        );

    \I__5644\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28706\
        );

    \I__5643\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28706\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__28711\,
            I => \N__28702\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__28706\,
            I => \N__28699\
        );

    \I__5640\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28696\
        );

    \I__5639\ : Span4Mux_v
    port map (
            O => \N__28702\,
            I => \N__28693\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__28699\,
            I => \N__28690\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__28696\,
            I => \N__28687\
        );

    \I__5636\ : Odrv4
    port map (
            O => \N__28693\,
            I => \b2v_inst11.func_state_RNI5DLRZ0Z_0\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__28690\,
            I => \b2v_inst11.func_state_RNI5DLRZ0Z_0\
        );

    \I__5634\ : Odrv4
    port map (
            O => \N__28687\,
            I => \b2v_inst11.func_state_RNI5DLRZ0Z_0\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__28680\,
            I => \N__28675\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__28679\,
            I => \N__28672\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__28678\,
            I => \N__28667\
        );

    \I__5630\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28663\
        );

    \I__5629\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28658\
        );

    \I__5628\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28658\
        );

    \I__5627\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28651\
        );

    \I__5626\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28651\
        );

    \I__5625\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28651\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28646\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28646\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28643\
        );

    \I__5621\ : Span4Mux_h
    port map (
            O => \N__28646\,
            I => \N__28640\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__28643\,
            I => \N__28637\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__28640\,
            I => \b2v_inst11.N_366\
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__28637\,
            I => \b2v_inst11.N_366\
        );

    \I__5617\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28623\
        );

    \I__5616\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28623\
        );

    \I__5615\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28618\
        );

    \I__5614\ : InMux
    port map (
            O => \N__28629\,
            I => \N__28618\
        );

    \I__5613\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28615\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__28623\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_0\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__28618\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_0\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__28615\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_0\
        );

    \I__5609\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__28605\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_313_N\
        );

    \I__5607\ : CascadeMux
    port map (
            O => \N__28602\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2BZ0_cascade_\
        );

    \I__5606\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__28596\,
            I => \b2v_inst11.dutycycle_1_0_1\
        );

    \I__5604\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__28590\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__5602\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28584\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28581\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__28581\,
            I => \N__28576\
        );

    \I__5599\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28573\
        );

    \I__5598\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28570\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__28576\,
            I => \b2v_inst11.count_clk_RNIG510TZ0Z_5\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__28573\,
            I => \b2v_inst11.count_clk_RNIG510TZ0Z_5\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__28570\,
            I => \b2v_inst11.count_clk_RNIG510TZ0Z_5\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__28563\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\
        );

    \I__5593\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__28557\,
            I => \b2v_inst11.un1_func_state25_6_0_1\
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__28554\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__28551\,
            I => \N__28540\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__28550\,
            I => \N__28537\
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__28549\,
            I => \N__28534\
        );

    \I__5587\ : CEMux
    port map (
            O => \N__28548\,
            I => \N__28528\
        );

    \I__5586\ : CEMux
    port map (
            O => \N__28547\,
            I => \N__28521\
        );

    \I__5585\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28512\
        );

    \I__5584\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28512\
        );

    \I__5583\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28512\
        );

    \I__5582\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28512\
        );

    \I__5581\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28503\
        );

    \I__5580\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28503\
        );

    \I__5579\ : InMux
    port map (
            O => \N__28534\,
            I => \N__28503\
        );

    \I__5578\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28503\
        );

    \I__5577\ : CEMux
    port map (
            O => \N__28532\,
            I => \N__28495\
        );

    \I__5576\ : CEMux
    port map (
            O => \N__28531\,
            I => \N__28492\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__28528\,
            I => \N__28489\
        );

    \I__5574\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28482\
        );

    \I__5573\ : InMux
    port map (
            O => \N__28526\,
            I => \N__28482\
        );

    \I__5572\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28482\
        );

    \I__5571\ : CEMux
    port map (
            O => \N__28524\,
            I => \N__28479\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__28521\,
            I => \N__28472\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__28512\,
            I => \N__28472\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__28503\,
            I => \N__28472\
        );

    \I__5567\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28469\
        );

    \I__5566\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28464\
        );

    \I__5565\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28464\
        );

    \I__5564\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28459\
        );

    \I__5563\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28459\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28456\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28453\
        );

    \I__5560\ : Span4Mux_v
    port map (
            O => \N__28489\,
            I => \N__28450\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__28482\,
            I => \N__28447\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28436\
        );

    \I__5557\ : Span4Mux_v
    port map (
            O => \N__28472\,
            I => \N__28436\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28436\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__28464\,
            I => \N__28436\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28436\
        );

    \I__5553\ : Span4Mux_h
    port map (
            O => \N__28456\,
            I => \N__28433\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__28453\,
            I => \N__28428\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__28450\,
            I => \N__28428\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__28447\,
            I => \N__28425\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__28436\,
            I => \N__28422\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__28433\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__28428\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__28425\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__28422\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__28413\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__28410\,
            I => \N__28384\
        );

    \I__5542\ : InMux
    port map (
            O => \N__28409\,
            I => \N__28379\
        );

    \I__5541\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28372\
        );

    \I__5540\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28372\
        );

    \I__5539\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28372\
        );

    \I__5538\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28365\
        );

    \I__5537\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28365\
        );

    \I__5536\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28365\
        );

    \I__5535\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28362\
        );

    \I__5534\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28353\
        );

    \I__5533\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28353\
        );

    \I__5532\ : InMux
    port map (
            O => \N__28399\,
            I => \N__28353\
        );

    \I__5531\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28353\
        );

    \I__5530\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28344\
        );

    \I__5529\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28344\
        );

    \I__5528\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28344\
        );

    \I__5527\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28340\
        );

    \I__5526\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28331\
        );

    \I__5525\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28331\
        );

    \I__5524\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28331\
        );

    \I__5523\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28331\
        );

    \I__5522\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28321\
        );

    \I__5521\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28314\
        );

    \I__5520\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28314\
        );

    \I__5519\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28311\
        );

    \I__5518\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28306\
        );

    \I__5517\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28306\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__28379\,
            I => \N__28295\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__28372\,
            I => \N__28295\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__28365\,
            I => \N__28295\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__28362\,
            I => \N__28295\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__28353\,
            I => \N__28295\
        );

    \I__5511\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28290\
        );

    \I__5510\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28290\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__28344\,
            I => \N__28287\
        );

    \I__5508\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28284\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28279\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28279\
        );

    \I__5505\ : InMux
    port map (
            O => \N__28330\,
            I => \N__28274\
        );

    \I__5504\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28274\
        );

    \I__5503\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28267\
        );

    \I__5502\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28267\
        );

    \I__5501\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28267\
        );

    \I__5500\ : CascadeMux
    port map (
            O => \N__28325\,
            I => \N__28264\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__28324\,
            I => \N__28261\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__28321\,
            I => \N__28254\
        );

    \I__5497\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28249\
        );

    \I__5496\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28249\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__28314\,
            I => \N__28242\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__28311\,
            I => \N__28242\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__28306\,
            I => \N__28242\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__28295\,
            I => \N__28235\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28235\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__28287\,
            I => \N__28226\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__28284\,
            I => \N__28226\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__28279\,
            I => \N__28226\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28226\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__28267\,
            I => \N__28223\
        );

    \I__5485\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28220\
        );

    \I__5484\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28215\
        );

    \I__5483\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28215\
        );

    \I__5482\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28212\
        );

    \I__5481\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28209\
        );

    \I__5480\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28206\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__28254\,
            I => \N__28203\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__28249\,
            I => \N__28200\
        );

    \I__5477\ : Span12Mux_s6_v
    port map (
            O => \N__28242\,
            I => \N__28197\
        );

    \I__5476\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28192\
        );

    \I__5475\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28192\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__28235\,
            I => \N__28185\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__28226\,
            I => \N__28185\
        );

    \I__5472\ : Span4Mux_h
    port map (
            O => \N__28223\,
            I => \N__28185\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28180\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__28215\,
            I => \N__28180\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__28212\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__28209\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__28206\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5466\ : Odrv4
    port map (
            O => \N__28203\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5465\ : Odrv4
    port map (
            O => \N__28200\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5464\ : Odrv12
    port map (
            O => \N__28197\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__28192\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__28185\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__28180\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__28161\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6_cascade_\
        );

    \I__5459\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28154\
        );

    \I__5458\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28151\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__28154\,
            I => \b2v_inst11.N_382_N\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__28151\,
            I => \b2v_inst11.N_382_N\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \N__28139\
        );

    \I__5454\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28136\
        );

    \I__5453\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28133\
        );

    \I__5452\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28130\
        );

    \I__5451\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28125\
        );

    \I__5450\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28125\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__28136\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__28133\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__28130\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__28125\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__5445\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28108\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__28115\,
            I => \N__28104\
        );

    \I__5443\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28097\
        );

    \I__5442\ : InMux
    port map (
            O => \N__28113\,
            I => \N__28097\
        );

    \I__5441\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28097\
        );

    \I__5440\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28094\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__28108\,
            I => \N__28091\
        );

    \I__5438\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28086\
        );

    \I__5437\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28086\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__28097\,
            I => \N__28082\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28079\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__28091\,
            I => \N__28073\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__28086\,
            I => \N__28073\
        );

    \I__5432\ : InMux
    port map (
            O => \N__28085\,
            I => \N__28070\
        );

    \I__5431\ : Span4Mux_v
    port map (
            O => \N__28082\,
            I => \N__28067\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__28079\,
            I => \N__28064\
        );

    \I__5429\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28061\
        );

    \I__5428\ : Odrv4
    port map (
            O => \N__28073\,
            I => \RSMRSTn_0\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__28070\,
            I => \RSMRSTn_0\
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__28067\,
            I => \RSMRSTn_0\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__28064\,
            I => \RSMRSTn_0\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__28061\,
            I => \RSMRSTn_0\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__28050\,
            I => \b2v_inst11.g0_4_sx_cascade_\
        );

    \I__5422\ : InMux
    port map (
            O => \N__28047\,
            I => \N__28044\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__28044\,
            I => \b2v_inst11.N_428\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__28041\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__28038\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_\
        );

    \I__5418\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28032\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__28032\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0\
        );

    \I__5416\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28023\
        );

    \I__5415\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28023\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__28023\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\
        );

    \I__5413\ : CascadeMux
    port map (
            O => \N__28020\,
            I => \b2v_inst11.func_state_1_m2_am_1_0_cascade_\
        );

    \I__5412\ : InMux
    port map (
            O => \N__28017\,
            I => \N__28014\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__28014\,
            I => \N__28011\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__28011\,
            I => \N__28008\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__28008\,
            I => \b2v_inst11.func_state_RNINCPR4Z0Z_0\
        );

    \I__5408\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27998\
        );

    \I__5407\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27998\
        );

    \I__5406\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27995\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__27998\,
            I => \b2v_inst11.N_382\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__27995\,
            I => \b2v_inst11.N_382\
        );

    \I__5403\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27987\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__27987\,
            I => \b2v_inst11.N_315\
        );

    \I__5401\ : IoInMux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__27981\,
            I => \N__27978\
        );

    \I__5399\ : Span4Mux_s3_h
    port map (
            O => \N__27978\,
            I => \N__27975\
        );

    \I__5398\ : Span4Mux_h
    port map (
            O => \N__27975\,
            I => \N__27972\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__27972\,
            I => \N__27969\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__27969\,
            I => vccst_en
        );

    \I__5395\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27963\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__27963\,
            I => \b2v_inst11.count_clk_RNIZ0Z_1\
        );

    \I__5393\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27951\
        );

    \I__5392\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27951\
        );

    \I__5391\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27951\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__27951\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__5389\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27939\
        );

    \I__5388\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27939\
        );

    \I__5387\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27939\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__27939\,
            I => \b2v_inst11.N_379\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__27936\,
            I => \b2v_inst11.count_clkZ0Z_3_cascade_\
        );

    \I__5384\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__27930\,
            I => \b2v_inst11.N_190\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__27927\,
            I => \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\
        );

    \I__5381\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27921\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__27921\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__5379\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27915\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__27915\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__27912\,
            I => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5Z0Z_0_cascade_\
        );

    \I__5376\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27903\
        );

    \I__5375\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27903\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__27903\,
            I => \b2v_inst11.count_clk_0_3\
        );

    \I__5373\ : InMux
    port map (
            O => \N__27900\,
            I => \N__27894\
        );

    \I__5372\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27894\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__27894\,
            I => \b2v_inst6.N_276_0\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__27891\,
            I => \b2v_inst6.curr_state_RNIKIRD1Z0Z_0_cascade_\
        );

    \I__5369\ : CascadeMux
    port map (
            O => \N__27888\,
            I => \N__27884\
        );

    \I__5368\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27879\
        );

    \I__5367\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27879\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__27879\,
            I => \b2v_inst6.delayed_vccin_vccinaux_ok_0\
        );

    \I__5365\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27869\
        );

    \I__5364\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27869\
        );

    \I__5363\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27866\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__27869\,
            I => \b2v_inst6.N_2992_i\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__27866\,
            I => \b2v_inst6.N_2992_i\
        );

    \I__5360\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27855\
        );

    \I__5359\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27848\
        );

    \I__5358\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27848\
        );

    \I__5357\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27848\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__27855\,
            I => \b2v_inst6.N_3011_i\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__27848\,
            I => \b2v_inst6.N_3011_i\
        );

    \I__5354\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27834\
        );

    \I__5353\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27834\
        );

    \I__5352\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27834\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27831\
        );

    \I__5350\ : Odrv4
    port map (
            O => \N__27831\,
            I => \b2v_inst6.N_192\
        );

    \I__5349\ : CascadeMux
    port map (
            O => \N__27828\,
            I => \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__5348\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \b2v_inst11.count_clkZ0Z_0_cascade_\
        );

    \I__5347\ : CascadeMux
    port map (
            O => \N__27822\,
            I => \b2v_inst11.count_clk_RNIZ0Z_1_cascade_\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__27819\,
            I => \b2v_inst11.un1_count_clk_2_axb_1_cascade_\
        );

    \I__5345\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27813\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__27813\,
            I => \b2v_inst11.count_clk_0_0\
        );

    \I__5343\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27804\
        );

    \I__5342\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27804\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__27804\,
            I => \b2v_inst11.count_clk_0_1\
        );

    \I__5340\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27798\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__27798\,
            I => \b2v_inst6.curr_state_1_0\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__27795\,
            I => \b2v_inst6.curr_state_7_0_cascade_\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__27792\,
            I => \b2v_inst6.count_RNICV5H1Z0Z_0_cascade_\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__27789\,
            I => \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\
        );

    \I__5335\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__27783\,
            I => \N__27779\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__27782\,
            I => \N__27774\
        );

    \I__5332\ : Span4Mux_h
    port map (
            O => \N__27779\,
            I => \N__27771\
        );

    \I__5331\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27766\
        );

    \I__5330\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27766\
        );

    \I__5329\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27763\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__27771\,
            I => \N__27754\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__27766\,
            I => \N__27754\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27754\
        );

    \I__5325\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27749\
        );

    \I__5324\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27749\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__27754\,
            I => \N__27744\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27744\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__27744\,
            I => \N__27741\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__27741\,
            I => \N_222\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__27738\,
            I => \b2v_inst6.N_2992_i_cascade_\
        );

    \I__5318\ : CascadeMux
    port map (
            O => \N__27735\,
            I => \N__27727\
        );

    \I__5317\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27718\
        );

    \I__5316\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27718\
        );

    \I__5315\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27718\
        );

    \I__5314\ : InMux
    port map (
            O => \N__27731\,
            I => \N__27718\
        );

    \I__5313\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27715\
        );

    \I__5312\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27712\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__27718\,
            I => \SYNTHESIZED_WIRE_8\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__27715\,
            I => \SYNTHESIZED_WIRE_8\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__27712\,
            I => \SYNTHESIZED_WIRE_8\
        );

    \I__5308\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__27702\,
            I => \N__27699\
        );

    \I__5306\ : IoSpan4Mux
    port map (
            O => \N__27699\,
            I => \N__27696\
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__27696\,
            I => v5s_ok
        );

    \I__5304\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__27690\,
            I => \N__27687\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__5300\ : Span4Mux_v
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__27678\,
            I => v33s_ok
        );

    \I__5298\ : IoInMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__5296\ : Span4Mux_s2_v
    port map (
            O => \N__27669\,
            I => \N__27665\
        );

    \I__5295\ : IoInMux
    port map (
            O => \N__27668\,
            I => \N__27662\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__27665\,
            I => \N__27659\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__27662\,
            I => \N__27656\
        );

    \I__5292\ : Span4Mux_v
    port map (
            O => \N__27659\,
            I => \N__27653\
        );

    \I__5291\ : Span4Mux_s3_h
    port map (
            O => \N__27656\,
            I => \N__27650\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__27653\,
            I => vccinaux_en
        );

    \I__5289\ : Odrv4
    port map (
            O => \N__27650\,
            I => vccinaux_en
        );

    \I__5288\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27642\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27637\
        );

    \I__5286\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27632\
        );

    \I__5285\ : InMux
    port map (
            O => \N__27640\,
            I => \N__27632\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__27637\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__27632\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__5282\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27622\
        );

    \I__5281\ : InMux
    port map (
            O => \N__27626\,
            I => \N__27619\
        );

    \I__5280\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27616\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__27622\,
            I => \b2v_inst6.curr_state_RNIKIRD1Z0Z_0\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__27619\,
            I => \b2v_inst6.curr_state_RNIKIRD1Z0Z_0\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__27616\,
            I => \b2v_inst6.curr_state_RNIKIRD1Z0Z_0\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__27609\,
            I => \b2v_inst6.un2_count_1_axb_9_cascade_\
        );

    \I__5275\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27600\
        );

    \I__5274\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27600\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__27600\,
            I => \b2v_inst6.count_rst_6\
        );

    \I__5272\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27591\
        );

    \I__5271\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27591\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__27591\,
            I => \b2v_inst6.count_rst_5\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__27588\,
            I => \b2v_inst6.countZ0Z_8_cascade_\
        );

    \I__5268\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27579\
        );

    \I__5267\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27579\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__27579\,
            I => \b2v_inst6.count_0_9\
        );

    \I__5265\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27570\
        );

    \I__5264\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27570\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__27570\,
            I => \b2v_inst6.count_0_8\
        );

    \I__5262\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27559\
        );

    \I__5261\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27552\
        );

    \I__5260\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27552\
        );

    \I__5259\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27552\
        );

    \I__5258\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27547\
        );

    \I__5257\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27547\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27530\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__27552\,
            I => \N__27527\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__27547\,
            I => \N__27524\
        );

    \I__5253\ : CEMux
    port map (
            O => \N__27546\,
            I => \N__27489\
        );

    \I__5252\ : CEMux
    port map (
            O => \N__27545\,
            I => \N__27489\
        );

    \I__5251\ : CEMux
    port map (
            O => \N__27544\,
            I => \N__27489\
        );

    \I__5250\ : CEMux
    port map (
            O => \N__27543\,
            I => \N__27489\
        );

    \I__5249\ : CEMux
    port map (
            O => \N__27542\,
            I => \N__27489\
        );

    \I__5248\ : CEMux
    port map (
            O => \N__27541\,
            I => \N__27489\
        );

    \I__5247\ : CEMux
    port map (
            O => \N__27540\,
            I => \N__27489\
        );

    \I__5246\ : CEMux
    port map (
            O => \N__27539\,
            I => \N__27489\
        );

    \I__5245\ : CEMux
    port map (
            O => \N__27538\,
            I => \N__27489\
        );

    \I__5244\ : CEMux
    port map (
            O => \N__27537\,
            I => \N__27489\
        );

    \I__5243\ : CEMux
    port map (
            O => \N__27536\,
            I => \N__27489\
        );

    \I__5242\ : CEMux
    port map (
            O => \N__27535\,
            I => \N__27489\
        );

    \I__5241\ : CEMux
    port map (
            O => \N__27534\,
            I => \N__27489\
        );

    \I__5240\ : CEMux
    port map (
            O => \N__27533\,
            I => \N__27489\
        );

    \I__5239\ : Glb2LocalMux
    port map (
            O => \N__27530\,
            I => \N__27489\
        );

    \I__5238\ : Glb2LocalMux
    port map (
            O => \N__27527\,
            I => \N__27489\
        );

    \I__5237\ : Glb2LocalMux
    port map (
            O => \N__27524\,
            I => \N__27489\
        );

    \I__5236\ : GlobalMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__5235\ : gio2CtrlBuf
    port map (
            O => \N__27486\,
            I => \N_607_g\
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \b2v_inst6.N_394_cascade_\
        );

    \I__5233\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__27474\,
            I => \b2v_inst6.curr_state_1_1\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__27471\,
            I => \b2v_inst6.m6_i_a3_cascade_\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__27468\,
            I => \N__27462\
        );

    \I__5228\ : InMux
    port map (
            O => \N__27467\,
            I => \N__27457\
        );

    \I__5227\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27457\
        );

    \I__5226\ : InMux
    port map (
            O => \N__27465\,
            I => \N__27452\
        );

    \I__5225\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27452\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__27457\,
            I => \N__27449\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__27452\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__27449\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__27444\,
            I => \b2v_inst6.curr_stateZ0Z_1_cascade_\
        );

    \I__5220\ : InMux
    port map (
            O => \N__27441\,
            I => \b2v_inst11.CO2\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \N__27434\
        );

    \I__5218\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27431\
        );

    \I__5217\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27428\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__27431\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__27428\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__5214\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27420\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__27420\,
            I => \b2v_inst11.mult1_un61_sum_i\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__27417\,
            I => \N__27414\
        );

    \I__5211\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__27411\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_13\
        );

    \I__5209\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27404\
        );

    \I__5208\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27401\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__27404\,
            I => \N__27398\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__27401\,
            I => \b2v_inst11.mult1_un47_sum_6\
        );

    \I__5205\ : Odrv4
    port map (
            O => \N__27398\,
            I => \b2v_inst11.mult1_un47_sum_6\
        );

    \I__5204\ : CascadeMux
    port map (
            O => \N__27393\,
            I => \N__27390\
        );

    \I__5203\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27386\
        );

    \I__5202\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27383\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__27386\,
            I => \N__27380\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__27383\,
            I => \b2v_inst11.mult1_un89_sum\
        );

    \I__5199\ : Odrv12
    port map (
            O => \N__27380\,
            I => \b2v_inst11.mult1_un89_sum\
        );

    \I__5198\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27372\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__27372\,
            I => \N__27369\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__27369\,
            I => \b2v_inst11.mult1_un89_sum_i\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__27366\,
            I => \b2v_inst6.un2_count_1_axb_8_cascade_\
        );

    \I__5194\ : InMux
    port map (
            O => \N__27363\,
            I => \bfn_8_15_0_\
        );

    \I__5193\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27356\
        );

    \I__5192\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27353\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__27356\,
            I => \N__27348\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__27353\,
            I => \N__27348\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__27345\,
            I => \b2v_inst11.mult1_un82_sum\
        );

    \I__5187\ : InMux
    port map (
            O => \N__27342\,
            I => \b2v_inst11.un1_dutycycle_53_cry_8\
        );

    \I__5186\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27336\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__27336\,
            I => \N__27332\
        );

    \I__5184\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27329\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__27332\,
            I => \N__27326\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27323\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__27326\,
            I => \b2v_inst11.mult1_un75_sum\
        );

    \I__5180\ : Odrv4
    port map (
            O => \N__27323\,
            I => \b2v_inst11.mult1_un75_sum\
        );

    \I__5179\ : InMux
    port map (
            O => \N__27318\,
            I => \b2v_inst11.un1_dutycycle_53_cry_9\
        );

    \I__5178\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27312\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__27312\,
            I => \N__27308\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__27311\,
            I => \N__27305\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__27308\,
            I => \N__27302\
        );

    \I__5174\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27299\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__27302\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__27299\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__5171\ : InMux
    port map (
            O => \N__27294\,
            I => \b2v_inst11.un1_dutycycle_53_cry_10\
        );

    \I__5170\ : InMux
    port map (
            O => \N__27291\,
            I => \b2v_inst11.un1_dutycycle_53_cry_11\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__27288\,
            I => \N__27285\
        );

    \I__5168\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27281\
        );

    \I__5167\ : CascadeMux
    port map (
            O => \N__27284\,
            I => \N__27278\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27275\
        );

    \I__5165\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27272\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__27275\,
            I => \b2v_inst11.mult1_un47_sum_1\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__27272\,
            I => \b2v_inst11.mult1_un47_sum_1\
        );

    \I__5162\ : InMux
    port map (
            O => \N__27267\,
            I => \b2v_inst11.un1_dutycycle_53_cry_12\
        );

    \I__5161\ : InMux
    port map (
            O => \N__27264\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13\
        );

    \I__5160\ : InMux
    port map (
            O => \N__27261\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14\
        );

    \I__5159\ : InMux
    port map (
            O => \N__27258\,
            I => \bfn_8_16_0_\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__5157\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__27249\,
            I => \N__27245\
        );

    \I__5155\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27242\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__27245\,
            I => \N__27239\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__27242\,
            I => \b2v_inst11.un1_dutycycle_53_axb_0\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__27239\,
            I => \b2v_inst11.un1_dutycycle_53_axb_0\
        );

    \I__5151\ : CascadeMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__5150\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__5148\ : Odrv12
    port map (
            O => \N__27225\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_0\
        );

    \I__5147\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27218\
        );

    \I__5146\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27215\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__27218\,
            I => \N__27212\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__27215\,
            I => \N__27209\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__27212\,
            I => \N__27206\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__27209\,
            I => \N__27203\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__27206\,
            I => \N__27200\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__27203\,
            I => \b2v_inst11.mult1_un138_sum\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__27200\,
            I => \b2v_inst11.mult1_un138_sum\
        );

    \I__5138\ : InMux
    port map (
            O => \N__27195\,
            I => \b2v_inst11.un1_dutycycle_53_cry_0\
        );

    \I__5137\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__27189\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_2\
        );

    \I__5135\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27182\
        );

    \I__5134\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27179\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__27182\,
            I => \N__27176\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27173\
        );

    \I__5131\ : Span4Mux_s2_v
    port map (
            O => \N__27176\,
            I => \N__27170\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__27173\,
            I => \b2v_inst11.mult1_un131_sum\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__27170\,
            I => \b2v_inst11.mult1_un131_sum\
        );

    \I__5128\ : InMux
    port map (
            O => \N__27165\,
            I => \b2v_inst11.un1_dutycycle_53_cry_1\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__27162\,
            I => \N__27159\
        );

    \I__5126\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__27156\,
            I => \N__27153\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__27150\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_2\
        );

    \I__5122\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27143\
        );

    \I__5121\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27140\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__27143\,
            I => \N__27137\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__27140\,
            I => \N__27134\
        );

    \I__5118\ : Span4Mux_v
    port map (
            O => \N__27137\,
            I => \N__27129\
        );

    \I__5117\ : Span4Mux_s2_v
    port map (
            O => \N__27134\,
            I => \N__27129\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__27129\,
            I => \b2v_inst11.mult1_un124_sum\
        );

    \I__5115\ : InMux
    port map (
            O => \N__27126\,
            I => \b2v_inst11.un1_dutycycle_53_cry_2\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__5113\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__27117\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5\
        );

    \I__5111\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27111\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__27111\,
            I => \N__27107\
        );

    \I__5109\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27104\
        );

    \I__5108\ : Span4Mux_s2_v
    port map (
            O => \N__27107\,
            I => \N__27101\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__27104\,
            I => \N__27098\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__27101\,
            I => \b2v_inst11.mult1_un117_sum\
        );

    \I__5105\ : Odrv12
    port map (
            O => \N__27098\,
            I => \b2v_inst11.mult1_un117_sum\
        );

    \I__5104\ : InMux
    port map (
            O => \N__27093\,
            I => \b2v_inst11.un1_dutycycle_53_cry_3\
        );

    \I__5103\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__27087\,
            I => \N__27083\
        );

    \I__5101\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27080\
        );

    \I__5100\ : Span4Mux_v
    port map (
            O => \N__27083\,
            I => \N__27075\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__27080\,
            I => \N__27075\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__27075\,
            I => \b2v_inst11.mult1_un110_sum\
        );

    \I__5097\ : InMux
    port map (
            O => \N__27072\,
            I => \b2v_inst11.un1_dutycycle_53_cry_4\
        );

    \I__5096\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27065\
        );

    \I__5095\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27062\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27059\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__27062\,
            I => \N__27056\
        );

    \I__5092\ : Span4Mux_s3_h
    port map (
            O => \N__27059\,
            I => \N__27053\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__27056\,
            I => \N__27050\
        );

    \I__5090\ : Span4Mux_h
    port map (
            O => \N__27053\,
            I => \N__27047\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__27050\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__27047\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__5087\ : InMux
    port map (
            O => \N__27042\,
            I => \b2v_inst11.un1_dutycycle_53_cry_5\
        );

    \I__5086\ : InMux
    port map (
            O => \N__27039\,
            I => \N__27035\
        );

    \I__5085\ : InMux
    port map (
            O => \N__27038\,
            I => \N__27032\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__27035\,
            I => \N__27029\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__27032\,
            I => \N__27026\
        );

    \I__5082\ : Span4Mux_v
    port map (
            O => \N__27029\,
            I => \N__27021\
        );

    \I__5081\ : Span4Mux_s2_v
    port map (
            O => \N__27026\,
            I => \N__27021\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__27021\,
            I => \b2v_inst11.mult1_un96_sum\
        );

    \I__5079\ : InMux
    port map (
            O => \N__27018\,
            I => \b2v_inst11.un1_dutycycle_53_cry_6\
        );

    \I__5078\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27009\
        );

    \I__5077\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27009\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__27009\,
            I => \b2v_inst11.dutycycle_RNI_10Z0Z_0\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__27006\,
            I => \b2v_inst11.dutycycle_RNIPKS23Z0Z_4_cascade_\
        );

    \I__5074\ : InMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__27000\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08UZ0\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__26997\,
            I => \N__26992\
        );

    \I__5071\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26985\
        );

    \I__5070\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26985\
        );

    \I__5069\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26985\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__26985\,
            I => \b2v_inst11.dutycycleZ1Z_4\
        );

    \I__5067\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26976\
        );

    \I__5066\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26976\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__26976\,
            I => \b2v_inst11.dutycycle_RNI5AV24Z0Z_4\
        );

    \I__5064\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26970\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__26970\,
            I => \b2v_inst11.dutycycle_RNIPKS23Z0Z_4\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__26967\,
            I => \b2v_inst11.dutycycleZ0Z_6_cascade_\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__26964\,
            I => \b2v_inst11.un1_i3_mux_cascade_\
        );

    \I__5060\ : InMux
    port map (
            O => \N__26961\,
            I => \N__26958\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__26958\,
            I => \b2v_inst11.d_i3_mux\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__26955\,
            I => \b2v_inst11.un1_dutycycle_172_m4_rn_0_cascade_\
        );

    \I__5057\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26949\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__26949\,
            I => \b2v_inst11.un1_dutycycle_172_m4\
        );

    \I__5055\ : InMux
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__26943\,
            I => \b2v_inst11.N_3057_0\
        );

    \I__5053\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26934\
        );

    \I__5052\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26934\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__26934\,
            I => \b2v_inst11.g1_0_0_0\
        );

    \I__5050\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__26928\,
            I => \b2v_inst11.N_3055_0_0\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__26925\,
            I => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_1_cascade_\
        );

    \I__5047\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__26919\,
            I => \b2v_inst11.g0_0_1\
        );

    \I__5045\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26910\
        );

    \I__5044\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26910\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__26910\,
            I => \b2v_inst11.g1_0_1_0\
        );

    \I__5042\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__26904\,
            I => \b2v_inst11.g0_3_2\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__26901\,
            I => \b2v_inst11.g2_1_0_1_cascade_\
        );

    \I__5039\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__26895\,
            I => \b2v_inst11.g2_1_0\
        );

    \I__5037\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__26889\,
            I => \b2v_inst11.dutycycle_RNI_9Z0Z_0\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \b2v_inst11.un1_dutycycle_172_m3_d_ns_1_0_cascade_\
        );

    \I__5034\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__26880\,
            I => \b2v_inst11.g1_1\
        );

    \I__5032\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26874\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__26874\,
            I => \b2v_inst11.dutycycle_RNIDQ4A1Z0Z_5\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__26871\,
            I => \b2v_inst11.un1_dutycycle_172_m4_rn_1_cascade_\
        );

    \I__5029\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__26865\,
            I => \b2v_inst11.dutycycle_RNI_11Z0Z_0\
        );

    \I__5027\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26856\
        );

    \I__5026\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26856\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__26856\,
            I => \N__26851\
        );

    \I__5024\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26848\
        );

    \I__5023\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26845\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__26851\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_5\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__26848\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_5\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__26845\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_5\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__26838\,
            I => \b2v_inst11.dutycycleZ1Z_5_cascade_\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__26835\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_5_cascade_\
        );

    \I__5017\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__26826\,
            I => \b2v_inst11.N_293\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__5013\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26814\
        );

    \I__5012\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26814\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__26814\,
            I => \N__26810\
        );

    \I__5010\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26807\
        );

    \I__5009\ : Span4Mux_h
    port map (
            O => \N__26810\,
            I => \N__26804\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__26807\,
            I => \b2v_inst11.N_365\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__26804\,
            I => \b2v_inst11.N_365\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__26799\,
            I => \b2v_inst11.N_159_cascade_\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__26796\,
            I => \b2v_inst11.func_state_1_m2_0_cascade_\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__26793\,
            I => \b2v_inst11.func_stateZ0Z_0_cascade_\
        );

    \I__5003\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__26787\,
            I => \b2v_inst11.func_state_1_m2_0\
        );

    \I__5001\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__26778\,
            I => \N__26770\
        );

    \I__4998\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26767\
        );

    \I__4997\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26762\
        );

    \I__4996\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26762\
        );

    \I__4995\ : InMux
    port map (
            O => \N__26774\,
            I => \N__26757\
        );

    \I__4994\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26757\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__26770\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__26767\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__26762\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__26757\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__4989\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26742\
        );

    \I__4988\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26742\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__26742\,
            I => \b2v_inst11.func_stateZ1Z_0\
        );

    \I__4986\ : CascadeMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__4985\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26725\
        );

    \I__4984\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26725\
        );

    \I__4983\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26725\
        );

    \I__4982\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26720\
        );

    \I__4981\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26720\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__26725\,
            I => \b2v_inst11.count_clk_en_0\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__26720\,
            I => \b2v_inst11.count_clk_en_0\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__26715\,
            I => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1_cascade_\
        );

    \I__4977\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__26709\,
            I => \b2v_inst11.un1_dutycycle_53_axb_3_1\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__26706\,
            I => \N__26703\
        );

    \I__4974\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__26700\,
            I => \b2v_inst11.d_N_5\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__4971\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26682\
        );

    \I__4970\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26682\
        );

    \I__4969\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26682\
        );

    \I__4968\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26682\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__26682\,
            I => \N__26677\
        );

    \I__4966\ : InMux
    port map (
            O => \N__26681\,
            I => \N__26674\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__26680\,
            I => \N__26666\
        );

    \I__4964\ : Span4Mux_h
    port map (
            O => \N__26677\,
            I => \N__26661\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__26674\,
            I => \N__26661\
        );

    \I__4962\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26658\
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__26672\,
            I => \N__26655\
        );

    \I__4960\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26645\
        );

    \I__4959\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26645\
        );

    \I__4958\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26645\
        );

    \I__4957\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26645\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__26661\,
            I => \N__26640\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__26658\,
            I => \N__26640\
        );

    \I__4954\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26635\
        );

    \I__4953\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26635\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__26645\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__26640\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__26635\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4949\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26622\
        );

    \I__4948\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26622\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__26622\,
            I => \b2v_inst11.func_state_1_ss0_i_0_o3_0\
        );

    \I__4946\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__26616\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_331_N\
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__26613\,
            I => \b2v_inst11.un1_func_state25_6_0_a3_0_1_cascade_\
        );

    \I__4943\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__26604\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_332_N\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__4939\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26594\
        );

    \I__4938\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26591\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__26594\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__26591\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__26586\,
            I => \b2v_inst11.N_337_cascade_\
        );

    \I__4934\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__26580\,
            I => \b2v_inst11.func_state_1_m2s2_i_1\
        );

    \I__4932\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__26574\,
            I => \b2v_inst11.N_76\
        );

    \I__4930\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26568\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__26568\,
            I => \b2v_inst11.func_state_RNI6IFF4_0Z0Z_1\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__26565\,
            I => \b2v_inst11.N_428_cascade_\
        );

    \I__4927\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26559\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__26559\,
            I => \b2v_inst11.count_clk_RNITV5AUZ0Z_7\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__26556\,
            I => \N__26549\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__26555\,
            I => \N__26544\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__26554\,
            I => \N__26541\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__26553\,
            I => \N__26538\
        );

    \I__4921\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26517\
        );

    \I__4920\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26517\
        );

    \I__4919\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26506\
        );

    \I__4918\ : InMux
    port map (
            O => \N__26547\,
            I => \N__26506\
        );

    \I__4917\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26506\
        );

    \I__4916\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26506\
        );

    \I__4915\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26506\
        );

    \I__4914\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26489\
        );

    \I__4913\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26489\
        );

    \I__4912\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26489\
        );

    \I__4911\ : InMux
    port map (
            O => \N__26534\,
            I => \N__26489\
        );

    \I__4910\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26489\
        );

    \I__4909\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26489\
        );

    \I__4908\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26489\
        );

    \I__4907\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26489\
        );

    \I__4906\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26474\
        );

    \I__4905\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26474\
        );

    \I__4904\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26474\
        );

    \I__4903\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26474\
        );

    \I__4902\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26474\
        );

    \I__4901\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26474\
        );

    \I__4900\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26474\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__26522\,
            I => \N__26468\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__26517\,
            I => \N__26461\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__26506\,
            I => \N__26461\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__26489\,
            I => \N__26452\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__26474\,
            I => \N__26452\
        );

    \I__4894\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26439\
        );

    \I__4893\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26439\
        );

    \I__4892\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26439\
        );

    \I__4891\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26439\
        );

    \I__4890\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26439\
        );

    \I__4889\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26439\
        );

    \I__4888\ : Span4Mux_h
    port map (
            O => \N__26461\,
            I => \N__26436\
        );

    \I__4887\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26427\
        );

    \I__4886\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26427\
        );

    \I__4885\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26427\
        );

    \I__4884\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26427\
        );

    \I__4883\ : Span4Mux_h
    port map (
            O => \N__26452\,
            I => \N__26424\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__26439\,
            I => \N__26421\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__26436\,
            I => \b2v_inst11.count_clk_RNILG61T1Z0Z_5\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__26427\,
            I => \b2v_inst11.count_clk_RNILG61T1Z0Z_5\
        );

    \I__4879\ : Odrv4
    port map (
            O => \N__26424\,
            I => \b2v_inst11.count_clk_RNILG61T1Z0Z_5\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__26421\,
            I => \b2v_inst11.count_clk_RNILG61T1Z0Z_5\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__26412\,
            I => \b2v_inst11.un1_func_state25_4_i_a2_sxZ0_cascade_\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__26409\,
            I => \rsmrstn_cascade_\
        );

    \I__4875\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26403\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__26403\,
            I => \N__26400\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__26400\,
            I => \N__26397\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__26397\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_0_2\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__26394\,
            I => \N__26391\
        );

    \I__4870\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26388\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26385\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__26385\,
            I => \N__26382\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__26382\,
            I => \N__26379\
        );

    \I__4866\ : Sp12to4
    port map (
            O => \N__26379\,
            I => \N__26376\
        );

    \I__4865\ : Odrv12
    port map (
            O => \N__26376\,
            I => vr_ready_vccin
        );

    \I__4864\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \b2v_inst6.N_192_cascade_\
        );

    \I__4863\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \b2v_inst6.N_241_cascade_\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \b2v_inst11.count_clk_RNIG8KAHZ0Z_7_cascade_\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__26364\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_\
        );

    \I__4860\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26358\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__26358\,
            I => \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__26355\,
            I => \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1_cascade_\
        );

    \I__4857\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26346\
        );

    \I__4856\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26346\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__26346\,
            I => \b2v_inst5.count_1_10\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__26343\,
            I => \b2v_inst5.count_rst_4_cascade_\
        );

    \I__4853\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__4851\ : Span4Mux_v
    port map (
            O => \N__26334\,
            I => \N__26331\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__26331\,
            I => \b2v_inst5.un12_clk_100khz_4\
        );

    \I__4849\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26325\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__26325\,
            I => \b2v_inst5.un12_clk_100khz_11\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__26322\,
            I => \b2v_inst5.un12_clk_100khz_5_cascade_\
        );

    \I__4846\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26316\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__26316\,
            I => \b2v_inst5.un12_clk_100khz_12\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__26313\,
            I => \b2v_inst5.N_1_i_cascade_\
        );

    \I__4843\ : CEMux
    port map (
            O => \N__26310\,
            I => \N__26307\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26303\
        );

    \I__4841\ : CEMux
    port map (
            O => \N__26306\,
            I => \N__26300\
        );

    \I__4840\ : Span4Mux_s0_v
    port map (
            O => \N__26303\,
            I => \N__26295\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__26300\,
            I => \N__26295\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__26295\,
            I => \N__26291\
        );

    \I__4837\ : CEMux
    port map (
            O => \N__26294\,
            I => \N__26288\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__26291\,
            I => \N__26282\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26282\
        );

    \I__4834\ : CEMux
    port map (
            O => \N__26287\,
            I => \N__26279\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__26282\,
            I => \N__26271\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__26279\,
            I => \N__26271\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__26278\,
            I => \N__26267\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__26277\,
            I => \N__26259\
        );

    \I__4829\ : CEMux
    port map (
            O => \N__26276\,
            I => \N__26247\
        );

    \I__4828\ : Span4Mux_v
    port map (
            O => \N__26271\,
            I => \N__26244\
        );

    \I__4827\ : CEMux
    port map (
            O => \N__26270\,
            I => \N__26233\
        );

    \I__4826\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26233\
        );

    \I__4825\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26233\
        );

    \I__4824\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26233\
        );

    \I__4823\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26233\
        );

    \I__4822\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26224\
        );

    \I__4821\ : InMux
    port map (
            O => \N__26262\,
            I => \N__26224\
        );

    \I__4820\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26224\
        );

    \I__4819\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26224\
        );

    \I__4818\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26216\
        );

    \I__4817\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26216\
        );

    \I__4816\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26209\
        );

    \I__4815\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26209\
        );

    \I__4814\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26209\
        );

    \I__4813\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26202\
        );

    \I__4812\ : InMux
    port map (
            O => \N__26251\,
            I => \N__26202\
        );

    \I__4811\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26202\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26193\
        );

    \I__4809\ : Span4Mux_s0_v
    port map (
            O => \N__26244\,
            I => \N__26193\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__26233\,
            I => \N__26193\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26193\
        );

    \I__4806\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26190\
        );

    \I__4805\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26185\
        );

    \I__4804\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26185\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__26216\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__26209\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__26202\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__26193\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__26190\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__26185\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__26172\,
            I => \N__26169\
        );

    \I__4796\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26166\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__26166\,
            I => \b2v_inst5.count_1_9\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__26163\,
            I => \N__26159\
        );

    \I__4793\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26156\
        );

    \I__4792\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26152\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N__26149\
        );

    \I__4790\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26146\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__26152\,
            I => \N__26143\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__26149\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__26146\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__26143\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__4785\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26132\
        );

    \I__4784\ : InMux
    port map (
            O => \N__26135\,
            I => \N__26129\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26126\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__26129\,
            I => \N__26123\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__26126\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__4780\ : Odrv12
    port map (
            O => \N__26123\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__4779\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26115\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26112\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__26112\,
            I => \b2v_inst5.count_rst_1\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__26109\,
            I => \N__26105\
        );

    \I__4775\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26091\
        );

    \I__4774\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26091\
        );

    \I__4773\ : InMux
    port map (
            O => \N__26104\,
            I => \N__26091\
        );

    \I__4772\ : InMux
    port map (
            O => \N__26103\,
            I => \N__26091\
        );

    \I__4771\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26091\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__26091\,
            I => \N__26082\
        );

    \I__4769\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26078\
        );

    \I__4768\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26075\
        );

    \I__4767\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26070\
        );

    \I__4766\ : InMux
    port map (
            O => \N__26087\,
            I => \N__26070\
        );

    \I__4765\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26065\
        );

    \I__4764\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26065\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__26082\,
            I => \N__26062\
        );

    \I__4762\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26059\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__26078\,
            I => \b2v_inst5.N_1_i\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__26075\,
            I => \b2v_inst5.N_1_i\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__26070\,
            I => \b2v_inst5.N_1_i\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__26065\,
            I => \b2v_inst5.N_1_i\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__26062\,
            I => \b2v_inst5.N_1_i\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__26059\,
            I => \b2v_inst5.N_1_i\
        );

    \I__4755\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26042\
        );

    \I__4754\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26039\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__26042\,
            I => \N__26036\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__26039\,
            I => \N__26031\
        );

    \I__4751\ : Span4Mux_s3_v
    port map (
            O => \N__26036\,
            I => \N__26031\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__26031\,
            I => \b2v_inst5.un2_count_1_cry_8_THRU_CO\
        );

    \I__4749\ : InMux
    port map (
            O => \N__26028\,
            I => \N__26024\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__26027\,
            I => \N__26021\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__4746\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26013\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__26018\,
            I => \N__26010\
        );

    \I__4744\ : InMux
    port map (
            O => \N__26017\,
            I => \N__26005\
        );

    \I__4743\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26005\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__26013\,
            I => \b2v_inst5.countZ0Z_9\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__26010\,
            I => \b2v_inst5.countZ0Z_9\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__26005\,
            I => \b2v_inst5.countZ0Z_9\
        );

    \I__4739\ : SRMux
    port map (
            O => \N__25998\,
            I => \N__25995\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__25995\,
            I => \N__25992\
        );

    \I__4737\ : Span4Mux_v
    port map (
            O => \N__25992\,
            I => \N__25985\
        );

    \I__4736\ : SRMux
    port map (
            O => \N__25991\,
            I => \N__25982\
        );

    \I__4735\ : SRMux
    port map (
            O => \N__25990\,
            I => \N__25971\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__25989\,
            I => \N__25967\
        );

    \I__4733\ : SRMux
    port map (
            O => \N__25988\,
            I => \N__25955\
        );

    \I__4732\ : Span4Mux_h
    port map (
            O => \N__25985\,
            I => \N__25950\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__25982\,
            I => \N__25950\
        );

    \I__4730\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25947\
        );

    \I__4729\ : SRMux
    port map (
            O => \N__25980\,
            I => \N__25944\
        );

    \I__4728\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25937\
        );

    \I__4727\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25937\
        );

    \I__4726\ : SRMux
    port map (
            O => \N__25977\,
            I => \N__25937\
        );

    \I__4725\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25934\
        );

    \I__4724\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25929\
        );

    \I__4723\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25929\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__25971\,
            I => \N__25926\
        );

    \I__4721\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25915\
        );

    \I__4720\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25915\
        );

    \I__4719\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25915\
        );

    \I__4718\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25915\
        );

    \I__4717\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25915\
        );

    \I__4716\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25904\
        );

    \I__4715\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25904\
        );

    \I__4714\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25904\
        );

    \I__4713\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25904\
        );

    \I__4712\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25904\
        );

    \I__4711\ : CascadeMux
    port map (
            O => \N__25958\,
            I => \N__25899\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__25955\,
            I => \N__25893\
        );

    \I__4709\ : Span4Mux_h
    port map (
            O => \N__25950\,
            I => \N__25884\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25884\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__25944\,
            I => \N__25884\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__25937\,
            I => \N__25884\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__25934\,
            I => \N__25879\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__25929\,
            I => \N__25876\
        );

    \I__4703\ : Span4Mux_s1_v
    port map (
            O => \N__25926\,
            I => \N__25869\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25869\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__25904\,
            I => \N__25869\
        );

    \I__4700\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25858\
        );

    \I__4699\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25858\
        );

    \I__4698\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25858\
        );

    \I__4697\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25858\
        );

    \I__4696\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25858\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__25896\,
            I => \N__25850\
        );

    \I__4694\ : Span4Mux_s1_v
    port map (
            O => \N__25893\,
            I => \N__25846\
        );

    \I__4693\ : Span4Mux_v
    port map (
            O => \N__25884\,
            I => \N__25843\
        );

    \I__4692\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25840\
        );

    \I__4691\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25837\
        );

    \I__4690\ : Span4Mux_s2_v
    port map (
            O => \N__25879\,
            I => \N__25832\
        );

    \I__4689\ : Span4Mux_h
    port map (
            O => \N__25876\,
            I => \N__25832\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__25869\,
            I => \N__25827\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25827\
        );

    \I__4686\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25816\
        );

    \I__4685\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25816\
        );

    \I__4684\ : InMux
    port map (
            O => \N__25855\,
            I => \N__25816\
        );

    \I__4683\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25816\
        );

    \I__4682\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25816\
        );

    \I__4681\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25811\
        );

    \I__4680\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25811\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__25846\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__25843\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__25840\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__25837\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__25832\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__25827\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__25816\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__25811\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__4671\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25791\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__25791\,
            I => \b2v_inst5.count_rst_5\
        );

    \I__4669\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25785\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__25785\,
            I => \N__25782\
        );

    \I__4667\ : Sp12to4
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__4666\ : Span12Mux_v
    port map (
            O => \N__25779\,
            I => \N__25776\
        );

    \I__4665\ : Odrv12
    port map (
            O => \N__25776\,
            I => v33a_ok
        );

    \I__4664\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25770\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__25770\,
            I => \N__25767\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__25767\,
            I => \N__25764\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__25764\,
            I => vccst_cpu_ok
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__25761\,
            I => \N__25758\
        );

    \I__4659\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25755\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__4656\ : Sp12to4
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__4655\ : Span12Mux_s11_v
    port map (
            O => \N__25746\,
            I => \N__25743\
        );

    \I__4654\ : Odrv12
    port map (
            O => \N__25743\,
            I => v1p8a_ok
        );

    \I__4653\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__4651\ : Span12Mux_s4_v
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__4650\ : Odrv12
    port map (
            O => \N__25731\,
            I => v5a_ok
        );

    \I__4649\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25725\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__25725\,
            I => \N__25722\
        );

    \I__4647\ : Span4Mux_v
    port map (
            O => \N__25722\,
            I => \N__25719\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__25719\,
            I => \N__25716\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__25716\,
            I => vr_ready_vccinaux
        );

    \I__4644\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25704\
        );

    \I__4643\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25704\
        );

    \I__4642\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25704\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__4640\ : Span4Mux_s3_v
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__4639\ : Odrv4
    port map (
            O => \N__25698\,
            I => \b2v_inst5.count_rst_3\
        );

    \I__4638\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25691\
        );

    \I__4637\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25688\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__25691\,
            I => \b2v_inst5.count_1_11\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__25688\,
            I => \b2v_inst5.count_1_11\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__25683\,
            I => \b2v_inst5.countZ0Z_7_cascade_\
        );

    \I__4633\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25674\
        );

    \I__4632\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25674\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__25674\,
            I => \N__25671\
        );

    \I__4630\ : Span4Mux_s2_v
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__25668\,
            I => \b2v_inst5.un2_count_1_cry_1_c_RNIMEQZ0Z9\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__25665\,
            I => \N__25662\
        );

    \I__4627\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__25659\,
            I => \b2v_inst5.count_1_2\
        );

    \I__4625\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25652\
        );

    \I__4624\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25649\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__25652\,
            I => \N__25646\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__25649\,
            I => \N__25643\
        );

    \I__4621\ : Span4Mux_h
    port map (
            O => \N__25646\,
            I => \N__25640\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__25643\,
            I => \b2v_inst5.countZ0Z_2\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__25640\,
            I => \b2v_inst5.countZ0Z_2\
        );

    \I__4618\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25628\
        );

    \I__4616\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25625\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__25628\,
            I => \N__25622\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__25625\,
            I => \N__25619\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__25622\,
            I => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__25619\,
            I => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__4610\ : InMux
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__25608\,
            I => \b2v_inst5.count_1_3\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__25605\,
            I => \b2v_inst5.un2_count_1_axb_10_cascade_\
        );

    \I__4607\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__25599\,
            I => \b2v_inst5.un12_clk_100khz_9\
        );

    \I__4605\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25592\
        );

    \I__4604\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__25592\,
            I => \b2v_inst5.countZ0Z_5\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__25589\,
            I => \b2v_inst5.countZ0Z_5\
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__4600\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25578\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__25578\,
            I => \b2v_inst5.un12_clk_100khz_1\
        );

    \I__4598\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__25572\,
            I => \N__25568\
        );

    \I__4596\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25565\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__25568\,
            I => \b2v_inst5.countZ0Z_6\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__25565\,
            I => \b2v_inst5.countZ0Z_6\
        );

    \I__4593\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__25557\,
            I => \N__25553\
        );

    \I__4591\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25550\
        );

    \I__4590\ : Span4Mux_h
    port map (
            O => \N__25553\,
            I => \N__25547\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__25550\,
            I => \b2v_inst5.un2_count_1_axb_10\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__25547\,
            I => \b2v_inst5.un2_count_1_axb_10\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__25542\,
            I => \N__25538\
        );

    \I__4586\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25533\
        );

    \I__4585\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25533\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__25527\,
            I => \b2v_inst5.un2_count_1_cry_9_THRU_CO\
        );

    \I__4581\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__25521\,
            I => \b2v_inst5.count_rst_4\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__25518\,
            I => \b2v_inst6.count_rst_10_cascade_\
        );

    \I__4578\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__25512\,
            I => \b2v_inst6.count_rst_11\
        );

    \I__4576\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25503\
        );

    \I__4575\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25503\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__25503\,
            I => \b2v_inst6.count_0_3\
        );

    \I__4573\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__25497\,
            I => \b2v_inst6.count_rst_10\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__25494\,
            I => \b2v_inst6.countZ0Z_3_cascade_\
        );

    \I__4570\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25485\
        );

    \I__4569\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25485\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__25485\,
            I => \b2v_inst6.count_0_4\
        );

    \I__4567\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25479\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__25473\,
            I => \b2v_inst5.un2_count_1_axb_11\
        );

    \I__4563\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__25467\,
            I => \b2v_inst5.count_1_7\
        );

    \I__4561\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25458\
        );

    \I__4560\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25458\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__4558\ : Span4Mux_s2_v
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__25452\,
            I => \b2v_inst5.un2_count_1_cry_6_c_RNIROVZ0Z9\
        );

    \I__4556\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__4554\ : Span4Mux_h
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__25440\,
            I => \b2v_inst5.countZ0Z_7\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__25437\,
            I => \N__25434\
        );

    \I__4551\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__25431\,
            I => \b2v_inst11.mult1_un68_sum_cry_4_s\
        );

    \I__4549\ : InMux
    port map (
            O => \N__25428\,
            I => \b2v_inst11.mult1_un68_sum_cry_3\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__4547\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__25419\,
            I => \b2v_inst11.mult1_un61_sum_cry_4_s\
        );

    \I__4545\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__25413\,
            I => \b2v_inst11.mult1_un68_sum_cry_5_s\
        );

    \I__4543\ : InMux
    port map (
            O => \N__25410\,
            I => \b2v_inst11.mult1_un68_sum_cry_4\
        );

    \I__4542\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__25404\,
            I => \b2v_inst11.mult1_un61_sum_cry_5_s\
        );

    \I__4540\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__25398\,
            I => \b2v_inst11.mult1_un68_sum_cry_6_s\
        );

    \I__4538\ : InMux
    port map (
            O => \N__25395\,
            I => \b2v_inst11.mult1_un68_sum_cry_5\
        );

    \I__4537\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__25389\,
            I => \b2v_inst11.mult1_un61_sum_cry_6_s\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__4534\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__25380\,
            I => \b2v_inst11.mult1_un75_sum_axb_8\
        );

    \I__4532\ : InMux
    port map (
            O => \N__25377\,
            I => \b2v_inst11.mult1_un68_sum_cry_6\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__4530\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25368\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__25368\,
            I => \b2v_inst11.mult1_un68_sum_axb_8\
        );

    \I__4528\ : InMux
    port map (
            O => \N__25365\,
            I => \b2v_inst11.mult1_un68_sum_cry_7\
        );

    \I__4527\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__4525\ : Span4Mux_s2_h
    port map (
            O => \N__25356\,
            I => \N__25352\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__25355\,
            I => \N__25348\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__25352\,
            I => \N__25343\
        );

    \I__4522\ : InMux
    port map (
            O => \N__25351\,
            I => \N__25340\
        );

    \I__4521\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25333\
        );

    \I__4520\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25333\
        );

    \I__4519\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25333\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__25343\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__25340\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__25333\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__4515\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25322\
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \N__25318\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25313\
        );

    \I__4512\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25310\
        );

    \I__4511\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25303\
        );

    \I__4510\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25303\
        );

    \I__4509\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25303\
        );

    \I__4508\ : Odrv12
    port map (
            O => \N__25313\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__25310\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__25303\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__25296\,
            I => \N__25292\
        );

    \I__4504\ : CascadeMux
    port map (
            O => \N__25295\,
            I => \N__25288\
        );

    \I__4503\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25281\
        );

    \I__4502\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25281\
        );

    \I__4501\ : InMux
    port map (
            O => \N__25288\,
            I => \N__25281\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__25281\,
            I => \b2v_inst11.mult1_un61_sum_i_0_8\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__25278\,
            I => \b2v_inst6.count_rst_11_cascade_\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__25275\,
            I => \b2v_inst6.un2_count_1_axb_3_cascade_\
        );

    \I__4497\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__25269\,
            I => \b2v_inst11.mult1_un54_sum_cry_3_s\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__25266\,
            I => \N__25263\
        );

    \I__4494\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25256\
        );

    \I__4493\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25256\
        );

    \I__4492\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25253\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__25256\,
            I => \b2v_inst11.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__25253\,
            I => \b2v_inst11.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__4489\ : InMux
    port map (
            O => \N__25248\,
            I => \b2v_inst11.mult1_un61_sum_cry_3\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__4487\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__25239\,
            I => \b2v_inst11.mult1_un54_sum_cry_4_s\
        );

    \I__4485\ : InMux
    port map (
            O => \N__25236\,
            I => \b2v_inst11.mult1_un61_sum_cry_4\
        );

    \I__4484\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25230\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__25230\,
            I => \b2v_inst11.mult1_un54_sum_cry_5_s\
        );

    \I__4482\ : InMux
    port map (
            O => \N__25227\,
            I => \b2v_inst11.mult1_un61_sum_cry_5\
        );

    \I__4481\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__25221\,
            I => \b2v_inst11.mult1_un54_sum_cry_6_s\
        );

    \I__4479\ : InMux
    port map (
            O => \N__25218\,
            I => \b2v_inst11.mult1_un61_sum_cry_6\
        );

    \I__4478\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25212\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__25212\,
            I => \b2v_inst11.mult1_un54_sum_cry_6_THRU_CO\
        );

    \I__4476\ : InMux
    port map (
            O => \N__25209\,
            I => \b2v_inst11.mult1_un61_sum_cry_7\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__25206\,
            I => \N__25202\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__25205\,
            I => \N__25199\
        );

    \I__4473\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25188\
        );

    \I__4472\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25188\
        );

    \I__4471\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25188\
        );

    \I__4470\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25188\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__25188\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__4467\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__25179\,
            I => \b2v_inst11.mult1_un54_sum_i_8\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__25176\,
            I => \N__25173\
        );

    \I__4464\ : InMux
    port map (
            O => \N__25173\,
            I => \N__25170\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__25170\,
            I => \b2v_inst11.mult1_un68_sum_cry_3_s\
        );

    \I__4462\ : InMux
    port map (
            O => \N__25167\,
            I => \b2v_inst11.mult1_un68_sum_cry_2\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__4460\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__25158\,
            I => \b2v_inst11.mult1_un61_sum_cry_3_s\
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__25155\,
            I => \N__25152\
        );

    \I__4457\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25149\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__25149\,
            I => \b2v_inst11.mult1_un54_sum_s_3_sf\
        );

    \I__4455\ : InMux
    port map (
            O => \N__25146\,
            I => \b2v_inst11.mult1_un54_sum_cry_2\
        );

    \I__4454\ : InMux
    port map (
            O => \N__25143\,
            I => \b2v_inst11.mult1_un54_sum_cry_3\
        );

    \I__4453\ : InMux
    port map (
            O => \N__25140\,
            I => \b2v_inst11.mult1_un54_sum_cry_4\
        );

    \I__4452\ : InMux
    port map (
            O => \N__25137\,
            I => \b2v_inst11.mult1_un54_sum_cry_5\
        );

    \I__4451\ : InMux
    port map (
            O => \N__25134\,
            I => \b2v_inst11.mult1_un54_sum_cry_6\
        );

    \I__4450\ : InMux
    port map (
            O => \N__25131\,
            I => \b2v_inst11.mult1_un54_sum_cry_7\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__4448\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__25119\,
            I => \b2v_inst11.mult1_un47_sum_i_1\
        );

    \I__4445\ : InMux
    port map (
            O => \N__25116\,
            I => \b2v_inst11.mult1_un61_sum_cry_2\
        );

    \I__4444\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__25110\,
            I => \b2v_inst11.g0_3_2_0\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__25107\,
            I => \b2v_inst11.un2_count_clk_17_0_a2_1_4_cascade_\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__25104\,
            I => \b2v_inst11.N_363_cascade_\
        );

    \I__4440\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__25095\,
            I => \b2v_inst11.mult1_un145_sum_i\
        );

    \I__4437\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25086\
        );

    \I__4435\ : Odrv12
    port map (
            O => \N__25086\,
            I => \b2v_inst11.mult1_un131_sum_i\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__25083\,
            I => \b2v_inst11.N_3055_0_cascade_\
        );

    \I__4433\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25077\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__25077\,
            I => \b2v_inst11.dutycycle_RNI_14Z0Z_0\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__25074\,
            I => \b2v_inst11.un1_dutycycle_172_m3_0_cascade_\
        );

    \I__4430\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__25068\,
            I => \b2v_inst11.un1_dutycycle_172_0\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__25065\,
            I => \b2v_inst11.N_19_i_cascade_\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__25062\,
            I => \b2v_inst11.un1_dutycycle_172_m0_ns_1_cascade_\
        );

    \I__4426\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__25056\,
            I => \b2v_inst11.un1_dutycycle_172_m0\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__25053\,
            I => \b2v_inst11.g0_4_1_cascade_\
        );

    \I__4423\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25047\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__25047\,
            I => \b2v_inst11.N_293_0\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__25044\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVKZ0_cascade_\
        );

    \I__4420\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__25038\,
            I => \b2v_inst11.N_236\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__25035\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\
        );

    \I__4417\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25029\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__25029\,
            I => \b2v_inst11.N_295\
        );

    \I__4415\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__25023\,
            I => \b2v_inst11.mult1_un152_sum_i\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__25020\,
            I => \v5s_enn_cascade_\
        );

    \I__4412\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__25014\,
            I => \N__25009\
        );

    \I__4410\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25006\
        );

    \I__4409\ : CascadeMux
    port map (
            O => \N__25012\,
            I => \N__25003\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__25009\,
            I => \N__24999\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24996\
        );

    \I__4406\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24991\
        );

    \I__4405\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24991\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__24999\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__24996\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__24991\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__4401\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__24981\,
            I => \b2v_inst20.un4_counter_0_and\
        );

    \I__4399\ : InMux
    port map (
            O => \N__24978\,
            I => \N__24975\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__4397\ : Odrv12
    port map (
            O => \N__24972\,
            I => \b2v_inst20.counter_1_cry_1_THRU_CO\
        );

    \I__4396\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24965\
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__24968\,
            I => \N__24962\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__24965\,
            I => \N__24958\
        );

    \I__4393\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24953\
        );

    \I__4392\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24953\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__24958\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__24953\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__4389\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__24945\,
            I => \N__24942\
        );

    \I__4387\ : Odrv12
    port map (
            O => \N__24942\,
            I => \b2v_inst20.counter_1_cry_2_THRU_CO\
        );

    \I__4386\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24935\
        );

    \I__4385\ : CascadeMux
    port map (
            O => \N__24938\,
            I => \N__24931\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__24935\,
            I => \N__24928\
        );

    \I__4383\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24923\
        );

    \I__4382\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24923\
        );

    \I__4381\ : Odrv12
    port map (
            O => \N__24928\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__24923\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__4379\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24915\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__4377\ : Odrv12
    port map (
            O => \N__24912\,
            I => \b2v_inst20.counter_1_cry_3_THRU_CO\
        );

    \I__4376\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__24906\,
            I => \N__24901\
        );

    \I__4374\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24896\
        );

    \I__4373\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24896\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__24901\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__24896\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__24891\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_1_cascade_\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__24888\,
            I => \N__24885\
        );

    \I__4368\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__24882\,
            I => \b2v_inst11.func_state_1_m2_1\
        );

    \I__4366\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24873\
        );

    \I__4365\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24873\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__24873\,
            I => \b2v_inst11.func_stateZ0Z_1\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__24870\,
            I => \b2v_inst11.un1_clk_100khz_51_and_i_a3_0_1_cascade_\
        );

    \I__4362\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__4360\ : Span4Mux_v
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__24858\,
            I => \N__24855\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__24852\,
            I => vpp_ok
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__24849\,
            I => \VCCST_EN_i_0_o3_0_cascade_\
        );

    \I__4355\ : IoInMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__4353\ : IoSpan4Mux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__4352\ : Span4Mux_s2_h
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__4351\ : Span4Mux_h
    port map (
            O => \N__24834\,
            I => \N__24831\
        );

    \I__4350\ : Span4Mux_v
    port map (
            O => \N__24831\,
            I => \N__24828\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__24828\,
            I => vddq_en
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__24825\,
            I => \b2v_inst11.count_clk_en_0_xZ0Z1_cascade_\
        );

    \I__4347\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__24819\,
            I => \N__24816\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__24816\,
            I => \b2v_inst11.N_335\
        );

    \I__4344\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24810\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__4342\ : Span4Mux_v
    port map (
            O => \N__24807\,
            I => \N__24803\
        );

    \I__4341\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24800\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__24803\,
            I => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__24800\,
            I => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\
        );

    \I__4338\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__24786\,
            I => \b2v_inst11.count_off_0_9\
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__24783\,
            I => \b2v_inst11.N_76_cascade_\
        );

    \I__4333\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24777\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__24777\,
            I => \b2v_inst11.func_state_RNICMPB4Z0Z_0\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__24774\,
            I => \b2v_inst11.func_state_1_m2_1_cascade_\
        );

    \I__4330\ : CascadeMux
    port map (
            O => \N__24771\,
            I => \b2v_inst11.func_state_cascade_\
        );

    \I__4329\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24765\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__24765\,
            I => \b2v_inst11.N_339\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__24762\,
            I => \b2v_inst11.N_339_cascade_\
        );

    \I__4326\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__24756\,
            I => \b2v_inst11.func_state_RNI6IFF4Z0Z_1\
        );

    \I__4324\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__24747\,
            I => \N__24744\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__24744\,
            I => \b2v_inst36.DSW_PWROK_0\
        );

    \I__4320\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24738\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__24738\,
            I => \b2v_inst36.curr_state_RNI3E27Z0Z_0\
        );

    \I__4318\ : IoInMux
    port map (
            O => \N__24735\,
            I => \N__24732\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__24732\,
            I => \N__24729\
        );

    \I__4316\ : Span4Mux_s2_h
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__24723\,
            I => dsw_pwrok
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__24720\,
            I => \curr_state_RNID8DP1_0_0_cascade_\
        );

    \I__4312\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24708\
        );

    \I__4311\ : InMux
    port map (
            O => \N__24716\,
            I => \N__24708\
        );

    \I__4310\ : InMux
    port map (
            O => \N__24715\,
            I => \N__24708\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__24708\,
            I => \N_413\
        );

    \I__4308\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__24702\,
            I => \b2v_inst5.curr_state_0_0\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__24699\,
            I => \N__24695\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__24698\,
            I => \N__24691\
        );

    \I__4304\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24684\
        );

    \I__4303\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24684\
        );

    \I__4302\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24684\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__24684\,
            I => \b2v_inst5.curr_stateZ0Z_0\
        );

    \I__4300\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24674\
        );

    \I__4299\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__4298\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24671\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__24674\,
            I => \b2v_inst5.N_2856_i\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__24671\,
            I => \b2v_inst5.N_2856_i\
        );

    \I__4295\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24659\
        );

    \I__4294\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24650\
        );

    \I__4293\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24650\
        );

    \I__4292\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24650\
        );

    \I__4291\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24650\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__24659\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__24650\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__24645\,
            I => \b2v_inst5.N_2856_i_cascade_\
        );

    \I__4287\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24639\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__24639\,
            I => \N__24636\
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__24636\,
            I => \b2v_inst11.count_off_0_7\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__24633\,
            I => \N__24629\
        );

    \I__4283\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24626\
        );

    \I__4282\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24623\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__24626\,
            I => \N__24620\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__24623\,
            I => \N__24617\
        );

    \I__4279\ : Span4Mux_h
    port map (
            O => \N__24620\,
            I => \N__24614\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__24617\,
            I => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__24614\,
            I => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__24609\,
            I => \N__24606\
        );

    \I__4275\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24602\
        );

    \I__4274\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24599\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__24602\,
            I => \N__24596\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__24599\,
            I => \b2v_inst11.count_offZ0Z_7\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__24596\,
            I => \b2v_inst11.count_offZ0Z_7\
        );

    \I__4270\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24588\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__4268\ : Span4Mux_h
    port map (
            O => \N__24585\,
            I => \N__24582\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__24582\,
            I => \b2v_inst11.un34_clk_100khz_11\
        );

    \I__4266\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24576\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__24576\,
            I => \b2v_inst11.un34_clk_100khz_9\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__4263\ : InMux
    port map (
            O => \N__24570\,
            I => \N__24567\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__24561\,
            I => \b2v_inst11.un34_clk_100khz_10\
        );

    \I__4259\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__24555\,
            I => \b2v_inst11.un34_clk_100khz_8\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__24552\,
            I => \b2v_inst11.count_off_RNI_1Z0Z_1_cascade_\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__24549\,
            I => \b2v_inst11.func_state_1_m0_0_0_1_cascade_\
        );

    \I__4255\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24540\
        );

    \I__4254\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24540\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__24537\,
            I => \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__24534\,
            I => \N__24531\
        );

    \I__4250\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24528\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__24528\,
            I => \b2v_inst11.count_off_0_8\
        );

    \I__4248\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24522\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__24522\,
            I => \N__24518\
        );

    \I__4246\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24515\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__24518\,
            I => \b2v_inst11.count_offZ0Z_8\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__24515\,
            I => \b2v_inst11.count_offZ0Z_8\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__24510\,
            I => \b2v_inst5.curr_stateZ0Z_1_cascade_\
        );

    \I__4242\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24501\
        );

    \I__4241\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24501\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__24501\,
            I => \b2v_inst5.count_1_0\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__4238\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24489\
        );

    \I__4237\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24489\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__24489\,
            I => \b2v_inst5.count_rst_14\
        );

    \I__4235\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24479\
        );

    \I__4234\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24479\
        );

    \I__4233\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24476\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__24479\,
            I => \b2v_inst5.count_i_0\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__24476\,
            I => \b2v_inst5.count_i_0\
        );

    \I__4230\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__24468\,
            I => \b2v_inst5.curr_stateZ0Z_1\
        );

    \I__4228\ : InMux
    port map (
            O => \N__24465\,
            I => \N__24462\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__24462\,
            I => \N__24459\
        );

    \I__4226\ : Odrv12
    port map (
            O => \N__24459\,
            I => \b2v_inst5.count_1_15\
        );

    \I__4225\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24453\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__24453\,
            I => \N__24450\
        );

    \I__4223\ : Span4Mux_s0_v
    port map (
            O => \N__24450\,
            I => \N__24446\
        );

    \I__4222\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24443\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__24446\,
            I => \b2v_inst5.count_rst\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__24443\,
            I => \b2v_inst5.count_rst\
        );

    \I__4219\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24435\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__24435\,
            I => \N__24431\
        );

    \I__4217\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24428\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__24431\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__24428\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__24423\,
            I => \b2v_inst5.curr_stateZ0Z_0_cascade_\
        );

    \I__4213\ : InMux
    port map (
            O => \N__24420\,
            I => \N__24414\
        );

    \I__4212\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24414\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__24414\,
            I => \b2v_inst5.N_51\
        );

    \I__4210\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24408\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__24408\,
            I => \b2v_inst5.m4_0\
        );

    \I__4208\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24399\
        );

    \I__4207\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24399\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__24399\,
            I => \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__4204\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__24390\,
            I => \b2v_inst5.count_1_12\
        );

    \I__4202\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__24384\,
            I => \b2v_inst5.count_1_14\
        );

    \I__4200\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24375\
        );

    \I__4199\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24375\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__24375\,
            I => \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\
        );

    \I__4197\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24369\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__24369\,
            I => \b2v_inst5.countZ0Z_14\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__24366\,
            I => \b2v_inst5.countZ0Z_14_cascade_\
        );

    \I__4194\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24359\
        );

    \I__4193\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24356\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__24359\,
            I => \b2v_inst5.countZ0Z_12\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__24356\,
            I => \b2v_inst5.countZ0Z_12\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__24351\,
            I => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_\
        );

    \I__4189\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__24345\,
            I => \b2v_inst5.un2_count_1_axb_0\
        );

    \I__4187\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24339\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__24339\,
            I => \b2v_inst5.curr_state_0_1\
        );

    \I__4185\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24330\
        );

    \I__4184\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24330\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__24330\,
            I => \b2v_inst5.un2_count_1_cry_4_c_RNIPKTZ0Z9\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__24327\,
            I => \N__24324\
        );

    \I__4181\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__24321\,
            I => \b2v_inst5.count_1_5\
        );

    \I__4179\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24314\
        );

    \I__4178\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24311\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__24314\,
            I => \b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__24311\,
            I => \b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__24306\,
            I => \N__24303\
        );

    \I__4174\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24300\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__24300\,
            I => \b2v_inst5.count_1_6\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__24297\,
            I => \b2v_inst5.countZ0Z_13_cascade_\
        );

    \I__4171\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24291\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__24291\,
            I => \b2v_inst5.count_1_13\
        );

    \I__4169\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__24285\,
            I => \b2v_inst5.countZ0Z_3\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__24282\,
            I => \b2v_inst5.countZ0Z_3_cascade_\
        );

    \I__4166\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24272\
        );

    \I__4164\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24269\
        );

    \I__4163\ : Odrv4
    port map (
            O => \N__24272\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__24269\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__4161\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24258\
        );

    \I__4160\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24258\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24255\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__24255\,
            I => \b2v_inst5.un2_count_1_cry_0_c_RNILCPZ0Z9\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__24252\,
            I => \N__24249\
        );

    \I__4156\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__24246\,
            I => \b2v_inst5.count_1_1\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__4153\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24237\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__24237\,
            I => \b2v_inst11.mult1_un75_sum_cry_4_s\
        );

    \I__4151\ : InMux
    port map (
            O => \N__24234\,
            I => \b2v_inst11.mult1_un75_sum_cry_3\
        );

    \I__4150\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24228\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__24228\,
            I => \b2v_inst11.mult1_un75_sum_cry_5_s\
        );

    \I__4148\ : InMux
    port map (
            O => \N__24225\,
            I => \b2v_inst11.mult1_un75_sum_cry_4\
        );

    \I__4147\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24219\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__24219\,
            I => \b2v_inst11.mult1_un75_sum_cry_6_s\
        );

    \I__4145\ : InMux
    port map (
            O => \N__24216\,
            I => \b2v_inst11.mult1_un75_sum_cry_5\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__24213\,
            I => \N__24210\
        );

    \I__4143\ : InMux
    port map (
            O => \N__24210\,
            I => \N__24207\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__24207\,
            I => \b2v_inst11.mult1_un82_sum_axb_8\
        );

    \I__4141\ : InMux
    port map (
            O => \N__24204\,
            I => \b2v_inst11.mult1_un75_sum_cry_6\
        );

    \I__4140\ : InMux
    port map (
            O => \N__24201\,
            I => \b2v_inst11.mult1_un75_sum_cry_7\
        );

    \I__4139\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24195\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__24195\,
            I => \N__24191\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__24194\,
            I => \N__24187\
        );

    \I__4136\ : Span4Mux_s3_h
    port map (
            O => \N__24191\,
            I => \N__24182\
        );

    \I__4135\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24179\
        );

    \I__4134\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24172\
        );

    \I__4133\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24172\
        );

    \I__4132\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24172\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__24182\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__24179\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__24172\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24161\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__24164\,
            I => \N__24157\
        );

    \I__4126\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24150\
        );

    \I__4125\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24150\
        );

    \I__4124\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24150\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__24150\,
            I => \b2v_inst11.mult1_un68_sum_i_0_8\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__24147\,
            I => \N__24144\
        );

    \I__4121\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__24141\,
            I => \b2v_inst11.mult1_un82_sum_cry_4_s\
        );

    \I__4119\ : InMux
    port map (
            O => \N__24138\,
            I => \b2v_inst11.mult1_un82_sum_cry_3\
        );

    \I__4118\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__24132\,
            I => \b2v_inst11.mult1_un82_sum_cry_5_s\
        );

    \I__4116\ : InMux
    port map (
            O => \N__24129\,
            I => \b2v_inst11.mult1_un82_sum_cry_4\
        );

    \I__4115\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24123\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__24123\,
            I => \b2v_inst11.mult1_un82_sum_cry_6_s\
        );

    \I__4113\ : InMux
    port map (
            O => \N__24120\,
            I => \b2v_inst11.mult1_un82_sum_cry_5\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__24117\,
            I => \N__24114\
        );

    \I__4111\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24111\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__24111\,
            I => \b2v_inst11.mult1_un89_sum_axb_8\
        );

    \I__4109\ : InMux
    port map (
            O => \N__24108\,
            I => \b2v_inst11.mult1_un82_sum_cry_6\
        );

    \I__4108\ : InMux
    port map (
            O => \N__24105\,
            I => \b2v_inst11.mult1_un82_sum_cry_7\
        );

    \I__4107\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24099\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__24099\,
            I => \N__24095\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__24098\,
            I => \N__24091\
        );

    \I__4104\ : Span4Mux_s2_v
    port map (
            O => \N__24095\,
            I => \N__24086\
        );

    \I__4103\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24083\
        );

    \I__4102\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24076\
        );

    \I__4101\ : InMux
    port map (
            O => \N__24090\,
            I => \N__24076\
        );

    \I__4100\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24076\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__24086\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__24083\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__24076\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__24069\,
            I => \N__24065\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__24068\,
            I => \N__24061\
        );

    \I__4094\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24054\
        );

    \I__4093\ : InMux
    port map (
            O => \N__24064\,
            I => \N__24054\
        );

    \I__4092\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24054\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__24054\,
            I => \b2v_inst11.mult1_un75_sum_i_0_8\
        );

    \I__4090\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24048\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24045\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__24045\,
            I => \b2v_inst11.mult1_un68_sum_i\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__24042\,
            I => \N__24039\
        );

    \I__4086\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24036\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__24036\,
            I => \b2v_inst11.mult1_un75_sum_cry_3_s\
        );

    \I__4084\ : InMux
    port map (
            O => \N__24033\,
            I => \b2v_inst11.mult1_un75_sum_cry_2\
        );

    \I__4083\ : InMux
    port map (
            O => \N__24030\,
            I => \b2v_inst11.mult1_un152_sum_cry_7\
        );

    \I__4082\ : InMux
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__24021\
        );

    \I__4080\ : Span4Mux_s2_h
    port map (
            O => \N__24021\,
            I => \N__24017\
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__24020\,
            I => \N__24013\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__24017\,
            I => \N__24009\
        );

    \I__4077\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24004\
        );

    \I__4076\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24004\
        );

    \I__4075\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24001\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__24009\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__24004\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__24001\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__23994\,
            I => \b2v_inst11.mult1_un152_sum_s_8_cascade_\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__23991\,
            I => \N__23987\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__23990\,
            I => \N__23983\
        );

    \I__4068\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23976\
        );

    \I__4067\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23976\
        );

    \I__4066\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23976\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__23976\,
            I => \b2v_inst11.mult1_un152_sum_i_0_8\
        );

    \I__4064\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23970\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23967\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__23967\,
            I => \b2v_inst11.mult1_un82_sum_i\
        );

    \I__4061\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__23961\,
            I => \N__23958\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__23958\,
            I => \N__23955\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__23955\,
            I => \b2v_inst11.mult1_un96_sum_i\
        );

    \I__4057\ : IoInMux
    port map (
            O => \N__23952\,
            I => \N__23949\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__23949\,
            I => \N__23946\
        );

    \I__4055\ : Span4Mux_s3_h
    port map (
            O => \N__23946\,
            I => \N__23942\
        );

    \I__4054\ : IoInMux
    port map (
            O => \N__23945\,
            I => \N__23938\
        );

    \I__4053\ : Span4Mux_v
    port map (
            O => \N__23942\,
            I => \N__23935\
        );

    \I__4052\ : IoInMux
    port map (
            O => \N__23941\,
            I => \N__23932\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__23938\,
            I => \N__23929\
        );

    \I__4050\ : Sp12to4
    port map (
            O => \N__23935\,
            I => \N__23926\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__23932\,
            I => \N__23923\
        );

    \I__4048\ : IoSpan4Mux
    port map (
            O => \N__23929\,
            I => \N__23920\
        );

    \I__4047\ : Span12Mux_s5_h
    port map (
            O => \N__23926\,
            I => \N__23915\
        );

    \I__4046\ : Span12Mux_s5_v
    port map (
            O => \N__23923\,
            I => \N__23915\
        );

    \I__4045\ : Sp12to4
    port map (
            O => \N__23920\,
            I => \N__23912\
        );

    \I__4044\ : Odrv12
    port map (
            O => \N__23915\,
            I => pch_pwrok
        );

    \I__4043\ : Odrv12
    port map (
            O => \N__23912\,
            I => pch_pwrok
        );

    \I__4042\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23904\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23901\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__23901\,
            I => \b2v_inst11.mult1_un75_sum_i\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__23898\,
            I => \N__23895\
        );

    \I__4038\ : InMux
    port map (
            O => \N__23895\,
            I => \N__23892\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__23892\,
            I => \b2v_inst11.mult1_un82_sum_cry_3_s\
        );

    \I__4036\ : InMux
    port map (
            O => \N__23889\,
            I => \b2v_inst11.mult1_un82_sum_cry_2\
        );

    \I__4035\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23882\
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__23885\,
            I => \N__23879\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23874\
        );

    \I__4032\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23866\
        );

    \I__4031\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23866\
        );

    \I__4030\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23866\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__23874\,
            I => \N__23863\
        );

    \I__4028\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23860\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__23866\,
            I => \N__23857\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__23863\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__23860\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__4024\ : Odrv4
    port map (
            O => \N__23857\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__4023\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23847\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__23847\,
            I => \N__23844\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__23844\,
            I => \b2v_inst11.mult1_un159_sum_i\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__23841\,
            I => \N__23838\
        );

    \I__4019\ : InMux
    port map (
            O => \N__23838\,
            I => \N__23835\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__23835\,
            I => \b2v_inst11.mult1_un145_sum_i_0_8\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__23832\,
            I => \N__23829\
        );

    \I__4016\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23826\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__23826\,
            I => \b2v_inst11.mult1_un152_sum_cry_3_s\
        );

    \I__4014\ : InMux
    port map (
            O => \N__23823\,
            I => \b2v_inst11.mult1_un152_sum_cry_2\
        );

    \I__4013\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23816\
        );

    \I__4012\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23813\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23810\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__23813\,
            I => \b2v_inst11.mult1_un145_sum_cry_3_s\
        );

    \I__4009\ : Odrv12
    port map (
            O => \N__23810\,
            I => \b2v_inst11.mult1_un145_sum_cry_3_s\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__23805\,
            I => \N__23802\
        );

    \I__4007\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23799\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__23799\,
            I => \b2v_inst11.mult1_un152_sum_axb_4_l_fx\
        );

    \I__4005\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23793\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__23793\,
            I => \b2v_inst11.mult1_un152_sum_cry_4_s\
        );

    \I__4003\ : InMux
    port map (
            O => \N__23790\,
            I => \b2v_inst11.mult1_un152_sum_cry_3\
        );

    \I__4002\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__23781\,
            I => \b2v_inst11.mult1_un145_sum_cry_4_s\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__23778\,
            I => \N__23775\
        );

    \I__3998\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23772\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__23772\,
            I => \b2v_inst11.mult1_un152_sum_cry_5_s\
        );

    \I__3996\ : InMux
    port map (
            O => \N__23769\,
            I => \b2v_inst11.mult1_un152_sum_cry_4\
        );

    \I__3995\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23762\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__23765\,
            I => \N__23758\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__23762\,
            I => \N__23755\
        );

    \I__3992\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23750\
        );

    \I__3991\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23750\
        );

    \I__3990\ : Span4Mux_v
    port map (
            O => \N__23755\,
            I => \N__23741\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__23750\,
            I => \N__23741\
        );

    \I__3988\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23738\
        );

    \I__3987\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23735\
        );

    \I__3986\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23730\
        );

    \I__3985\ : InMux
    port map (
            O => \N__23746\,
            I => \N__23730\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__23741\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__23738\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__23735\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__23730\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__23721\,
            I => \N__23718\
        );

    \I__3979\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23715\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23712\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__23712\,
            I => \b2v_inst11.mult1_un145_sum_cry_5_s\
        );

    \I__3976\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23706\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__23706\,
            I => \b2v_inst11.mult1_un152_sum_cry_6_s\
        );

    \I__3974\ : InMux
    port map (
            O => \N__23703\,
            I => \b2v_inst11.mult1_un152_sum_cry_5\
        );

    \I__3973\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23696\
        );

    \I__3972\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23693\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__23696\,
            I => \N__23690\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__23693\,
            I => \b2v_inst11.mult1_un145_sum_cry_6_s\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__23690\,
            I => \b2v_inst11.mult1_un145_sum_cry_6_s\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__3967\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__23679\,
            I => \b2v_inst11.mult1_un152_sum_axb_7_l_fx\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__3964\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__23670\,
            I => \b2v_inst11.mult1_un159_sum_axb_7\
        );

    \I__3962\ : InMux
    port map (
            O => \N__23667\,
            I => \b2v_inst11.mult1_un152_sum_cry_6\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__3960\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23658\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__23655\,
            I => \b2v_inst11.mult1_un152_sum_axb_8\
        );

    \I__3957\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23648\
        );

    \I__3956\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23645\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__23648\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__23645\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__3953\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23636\
        );

    \I__3952\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23633\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__23636\,
            I => \N__23630\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__23633\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__23630\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__3947\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23618\
        );

    \I__3946\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23615\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23612\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__23615\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__23612\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__3942\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23603\
        );

    \I__3941\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23600\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23597\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__23600\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__23597\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__3937\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23589\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__23589\,
            I => \b2v_inst20.un4_counter_6_and\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__3934\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23580\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__23580\,
            I => \N__23577\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__23577\,
            I => \b2v_inst11.mult1_un159_sum_cry_2_s\
        );

    \I__3931\ : InMux
    port map (
            O => \N__23574\,
            I => \b2v_inst11.mult1_un159_sum_cry_1\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__23571\,
            I => \N__23568\
        );

    \I__3929\ : InMux
    port map (
            O => \N__23568\,
            I => \N__23565\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23562\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__23562\,
            I => \b2v_inst11.mult1_un159_sum_cry_3_s\
        );

    \I__3926\ : InMux
    port map (
            O => \N__23559\,
            I => \b2v_inst11.mult1_un159_sum_cry_2\
        );

    \I__3925\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23553\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__23553\,
            I => \N__23550\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__23550\,
            I => \b2v_inst11.mult1_un159_sum_cry_4_s\
        );

    \I__3922\ : InMux
    port map (
            O => \N__23547\,
            I => \b2v_inst11.mult1_un159_sum_cry_3\
        );

    \I__3921\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23541\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__23541\,
            I => \N__23538\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__23538\,
            I => \b2v_inst11.mult1_un159_sum_cry_5_s\
        );

    \I__3918\ : InMux
    port map (
            O => \N__23535\,
            I => \b2v_inst11.mult1_un159_sum_cry_4\
        );

    \I__3917\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23529\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__23526\,
            I => \b2v_inst11.mult1_un166_sum_axb_6\
        );

    \I__3914\ : InMux
    port map (
            O => \N__23523\,
            I => \b2v_inst11.mult1_un159_sum_cry_5\
        );

    \I__3913\ : InMux
    port map (
            O => \N__23520\,
            I => \b2v_inst11.mult1_un159_sum_cry_6\
        );

    \I__3912\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23514\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23511\
        );

    \I__3910\ : Span4Mux_h
    port map (
            O => \N__23511\,
            I => \N__23508\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__23508\,
            I => \b2v_inst20.un4_counter_5_and\
        );

    \I__3908\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23502\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__23502\,
            I => \b2v_inst20.un4_counter_7_and\
        );

    \I__3906\ : InMux
    port map (
            O => \N__23499\,
            I => \bfn_6_10_0_\
        );

    \I__3905\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23492\
        );

    \I__3904\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23489\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__23492\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__23489\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__3901\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23480\
        );

    \I__3900\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23477\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__23480\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__23477\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__23472\,
            I => \N__23468\
        );

    \I__3896\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23465\
        );

    \I__3895\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23462\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__23465\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__23462\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__3892\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23453\
        );

    \I__3891\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__23453\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__23450\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__3888\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23442\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__23442\,
            I => \b2v_inst20.un4_counter_4_and\
        );

    \I__3886\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23435\
        );

    \I__3885\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23432\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__23435\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__23432\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__3882\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23423\
        );

    \I__3881\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23420\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__23423\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__23420\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__23415\,
            I => \N__23411\
        );

    \I__3877\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23408\
        );

    \I__3876\ : InMux
    port map (
            O => \N__23411\,
            I => \N__23405\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__23408\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__23405\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__3873\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23396\
        );

    \I__3872\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23393\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__23396\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__23393\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__3869\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__23385\,
            I => \b2v_inst20.un4_counter_3_and\
        );

    \I__3867\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23379\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__23379\,
            I => \b2v_inst11.count_off_0_5\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__3864\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23367\
        );

    \I__3863\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23367\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__23364\,
            I => \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__23361\,
            I => \N__23357\
        );

    \I__3859\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__3858\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23351\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23346\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__23351\,
            I => \N__23346\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__23346\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__3854\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__23340\,
            I => \b2v_inst11.count_off_0_6\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__23337\,
            I => \N__23334\
        );

    \I__3851\ : InMux
    port map (
            O => \N__23334\,
            I => \N__23330\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__23333\,
            I => \N__23327\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23324\
        );

    \I__3848\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23321\
        );

    \I__3847\ : Span4Mux_v
    port map (
            O => \N__23324\,
            I => \N__23318\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23315\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__23318\,
            I => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__23315\,
            I => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__3842\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23303\
        );

    \I__3841\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23300\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23297\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23294\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__23297\,
            I => \N__23291\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__23294\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__23291\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__3835\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23283\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__23283\,
            I => \N__23280\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__23280\,
            I => \b2v_inst20.un4_counter_1_and\
        );

    \I__3832\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__3830\ : Span4Mux_v
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__23268\,
            I => \b2v_inst20.un4_counter_2_and\
        );

    \I__3828\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__23259\,
            I => \b2v_inst20.counter_1_cry_4_THRU_CO\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__3824\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23245\
        );

    \I__3822\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23240\
        );

    \I__3821\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23240\
        );

    \I__3820\ : Odrv4
    port map (
            O => \N__23245\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__23240\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3818\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23232\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__23232\,
            I => \N__23229\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__23229\,
            I => \b2v_inst20.counter_1_cry_5_THRU_CO\
        );

    \I__3815\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23222\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__23225\,
            I => \N__23218\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__23222\,
            I => \N__23215\
        );

    \I__3812\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23210\
        );

    \I__3811\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23210\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__23215\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__23210\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__23205\,
            I => \N__23202\
        );

    \I__3807\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23198\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \N__23195\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__23198\,
            I => \N__23192\
        );

    \I__3804\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23189\
        );

    \I__3803\ : Span4Mux_v
    port map (
            O => \N__23192\,
            I => \N__23186\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__23189\,
            I => \N__23183\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__23186\,
            I => \b2v_inst11.count_offZ0Z_3\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__23183\,
            I => \b2v_inst11.count_offZ0Z_3\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__23178\,
            I => \N__23175\
        );

    \I__3798\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23172\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23169\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__23169\,
            I => \N__23164\
        );

    \I__3795\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23159\
        );

    \I__3794\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23159\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__23164\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__23159\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3791\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23134\
        );

    \I__3790\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23134\
        );

    \I__3789\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23134\
        );

    \I__3788\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23134\
        );

    \I__3787\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23134\
        );

    \I__3786\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23134\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__23148\,
            I => \N__23131\
        );

    \I__3784\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23128\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__23134\,
            I => \N__23125\
        );

    \I__3782\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23122\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23119\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__23125\,
            I => \N__23114\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23114\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__23119\,
            I => \N__23111\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__23111\,
            I => \N__23105\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__23108\,
            I => \N__23102\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__23105\,
            I => \N__23099\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__23102\,
            I => \N__23096\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__23099\,
            I => v33dsw_ok
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__23096\,
            I => v33dsw_ok
        );

    \I__3770\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23087\
        );

    \I__3769\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23083\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__23087\,
            I => \N__23079\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__23086\,
            I => \N__23076\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__23083\,
            I => \N__23073\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__23082\,
            I => \N__23069\
        );

    \I__3764\ : Span4Mux_h
    port map (
            O => \N__23079\,
            I => \N__23064\
        );

    \I__3763\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23061\
        );

    \I__3762\ : Span4Mux_s3_h
    port map (
            O => \N__23073\,
            I => \N__23058\
        );

    \I__3761\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23049\
        );

    \I__3760\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23049\
        );

    \I__3759\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23049\
        );

    \I__3758\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23049\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__23064\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__23061\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__23058\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__23049\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__3753\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__23037\,
            I => \N__23033\
        );

    \I__3751\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23030\
        );

    \I__3750\ : Span4Mux_v
    port map (
            O => \N__23033\,
            I => \N__23026\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__23030\,
            I => \N__23023\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__23029\,
            I => \N__23017\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__23026\,
            I => \N__23013\
        );

    \I__3746\ : Span4Mux_s3_h
    port map (
            O => \N__23023\,
            I => \N__23010\
        );

    \I__3745\ : InMux
    port map (
            O => \N__23022\,
            I => \N__22999\
        );

    \I__3744\ : InMux
    port map (
            O => \N__23021\,
            I => \N__22999\
        );

    \I__3743\ : InMux
    port map (
            O => \N__23020\,
            I => \N__22999\
        );

    \I__3742\ : InMux
    port map (
            O => \N__23017\,
            I => \N__22999\
        );

    \I__3741\ : InMux
    port map (
            O => \N__23016\,
            I => \N__22999\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__23013\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__23010\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__22999\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__22992\,
            I => \N__22989\
        );

    \I__3736\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22985\
        );

    \I__3735\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22982\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22979\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__22982\,
            I => \b2v_inst11.count_offZ0Z_4\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__22979\,
            I => \b2v_inst11.count_offZ0Z_4\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__22974\,
            I => \N__22971\
        );

    \I__3730\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22965\
        );

    \I__3729\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22965\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22962\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__22962\,
            I => \N__22959\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__22959\,
            I => \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\
        );

    \I__3725\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22953\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__22953\,
            I => \b2v_inst11.count_off_0_4\
        );

    \I__3723\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22946\
        );

    \I__3722\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22943\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__22946\,
            I => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__22943\,
            I => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\
        );

    \I__3719\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__22935\,
            I => \N__22932\
        );

    \I__3717\ : Odrv12
    port map (
            O => \N__22932\,
            I => \b2v_inst11.count_off_0_15\
        );

    \I__3716\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__22926\,
            I => \b2v_inst11.count_off_0_2\
        );

    \I__3714\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22917\
        );

    \I__3713\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22917\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__22917\,
            I => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__22914\,
            I => \N__22911\
        );

    \I__3710\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__22908\,
            I => \b2v_inst11.count_off_0_0\
        );

    \I__3708\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22902\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__22902\,
            I => \N__22896\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__22901\,
            I => \N__22893\
        );

    \I__3705\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22888\
        );

    \I__3704\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22888\
        );

    \I__3703\ : Span4Mux_h
    port map (
            O => \N__22896\,
            I => \N__22885\
        );

    \I__3702\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22882\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__22888\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__3700\ : Odrv4
    port map (
            O => \N__22885\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__22882\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \b2v_inst11.count_offZ0Z_0_cascade_\
        );

    \I__3697\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__22869\,
            I => \b2v_inst11.count_off_RNIZ0Z_1\
        );

    \I__3695\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__22863\,
            I => \b2v_inst11.count_off_0_1\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__22860\,
            I => \b2v_inst11.count_off_RNIZ0Z_1_cascade_\
        );

    \I__3692\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22853\
        );

    \I__3691\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22850\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__22853\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__22850\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__22845\,
            I => \b2v_inst11.count_offZ0Z_1_cascade_\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__22842\,
            I => \N__22838\
        );

    \I__3686\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22835\
        );

    \I__3685\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22832\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__22835\,
            I => \b2v_inst11.count_offZ0Z_2\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__22832\,
            I => \b2v_inst11.count_offZ0Z_2\
        );

    \I__3682\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22823\
        );

    \I__3681\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22820\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22817\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__22820\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__22817\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__3677\ : InMux
    port map (
            O => \N__22812\,
            I => \b2v_inst5.un2_count_1_cry_14\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__22809\,
            I => \b2v_inst5.countZ0Z_4_cascade_\
        );

    \I__3675\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__22803\,
            I => \b2v_inst5.count_rst_6\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__22800\,
            I => \b2v_inst5.count_rst_6_cascade_\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__22797\,
            I => \N__22793\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__22796\,
            I => \N__22790\
        );

    \I__3670\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22787\
        );

    \I__3669\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22784\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__22787\,
            I => \b2v_inst5.un2_count_1_axb_8\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__22784\,
            I => \b2v_inst5.un2_count_1_axb_8\
        );

    \I__3666\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22773\
        );

    \I__3665\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22773\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__22773\,
            I => \b2v_inst5.un2_count_1_cry_7_THRU_CO\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__22770\,
            I => \b2v_inst5.un2_count_1_axb_8_cascade_\
        );

    \I__3662\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22761\
        );

    \I__3661\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22761\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__22761\,
            I => \b2v_inst5.count_1_8\
        );

    \I__3659\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22755\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__22755\,
            I => \b2v_inst5.count_rst_10\
        );

    \I__3657\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22746\
        );

    \I__3656\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22746\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__22743\,
            I => \b2v_inst5.un2_count_1_cry_3_THRU_CO\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__22740\,
            I => \N__22736\
        );

    \I__3652\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22732\
        );

    \I__3651\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22727\
        );

    \I__3650\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22727\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22724\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__22727\,
            I => \b2v_inst5.countZ0Z_4\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__22724\,
            I => \b2v_inst5.countZ0Z_4\
        );

    \I__3646\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__22716\,
            I => \b2v_inst5.count_1_4\
        );

    \I__3644\ : InMux
    port map (
            O => \N__22713\,
            I => \b2v_inst5.un2_count_1_cry_5\
        );

    \I__3643\ : InMux
    port map (
            O => \N__22710\,
            I => \b2v_inst5.un2_count_1_cry_6\
        );

    \I__3642\ : InMux
    port map (
            O => \N__22707\,
            I => \bfn_6_4_0_\
        );

    \I__3641\ : InMux
    port map (
            O => \N__22704\,
            I => \b2v_inst5.un2_count_1_cry_8\
        );

    \I__3640\ : InMux
    port map (
            O => \N__22701\,
            I => \b2v_inst5.un2_count_1_cry_9\
        );

    \I__3639\ : InMux
    port map (
            O => \N__22698\,
            I => \b2v_inst5.un2_count_1_cry_10\
        );

    \I__3638\ : InMux
    port map (
            O => \N__22695\,
            I => \b2v_inst5.un2_count_1_cry_11\
        );

    \I__3637\ : InMux
    port map (
            O => \N__22692\,
            I => \b2v_inst5.un2_count_1_cry_12\
        );

    \I__3636\ : InMux
    port map (
            O => \N__22689\,
            I => \b2v_inst5.un2_count_1_cry_13\
        );

    \I__3635\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22682\
        );

    \I__3634\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22679\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__22682\,
            I => \b2v_inst200.count_1_6\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__22679\,
            I => \b2v_inst200.count_1_6\
        );

    \I__3631\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22671\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__22671\,
            I => \b2v_inst200.count_3_6\
        );

    \I__3629\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22664\
        );

    \I__3628\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22661\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__22664\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__22661\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__3625\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__22653\,
            I => \b2v_inst200.count_3_7\
        );

    \I__3623\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22646\
        );

    \I__3622\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22643\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22640\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__22643\,
            I => \b2v_inst200.count_1_10\
        );

    \I__3619\ : Odrv4
    port map (
            O => \N__22640\,
            I => \b2v_inst200.count_1_10\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__22635\,
            I => \N__22632\
        );

    \I__3617\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22629\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__22629\,
            I => \b2v_inst200.count_3_10\
        );

    \I__3615\ : InMux
    port map (
            O => \N__22626\,
            I => \N__22590\
        );

    \I__3614\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22590\
        );

    \I__3613\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22590\
        );

    \I__3612\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22590\
        );

    \I__3611\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22590\
        );

    \I__3610\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22579\
        );

    \I__3609\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22579\
        );

    \I__3608\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22579\
        );

    \I__3607\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22579\
        );

    \I__3606\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22579\
        );

    \I__3605\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22574\
        );

    \I__3604\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22574\
        );

    \I__3603\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22565\
        );

    \I__3602\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22565\
        );

    \I__3601\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22565\
        );

    \I__3600\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22565\
        );

    \I__3599\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22552\
        );

    \I__3598\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22552\
        );

    \I__3597\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22552\
        );

    \I__3596\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22552\
        );

    \I__3595\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22552\
        );

    \I__3594\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22552\
        );

    \I__3593\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22543\
        );

    \I__3592\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22543\
        );

    \I__3591\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22543\
        );

    \I__3590\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22543\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22534\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__22579\,
            I => \N__22531\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__22574\,
            I => \N__22528\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22525\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__22552\,
            I => \N__22522\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22519\
        );

    \I__3583\ : CEMux
    port map (
            O => \N__22542\,
            I => \N__22494\
        );

    \I__3582\ : CEMux
    port map (
            O => \N__22541\,
            I => \N__22494\
        );

    \I__3581\ : CEMux
    port map (
            O => \N__22540\,
            I => \N__22494\
        );

    \I__3580\ : CEMux
    port map (
            O => \N__22539\,
            I => \N__22494\
        );

    \I__3579\ : CEMux
    port map (
            O => \N__22538\,
            I => \N__22494\
        );

    \I__3578\ : CEMux
    port map (
            O => \N__22537\,
            I => \N__22494\
        );

    \I__3577\ : Glb2LocalMux
    port map (
            O => \N__22534\,
            I => \N__22494\
        );

    \I__3576\ : Glb2LocalMux
    port map (
            O => \N__22531\,
            I => \N__22494\
        );

    \I__3575\ : Glb2LocalMux
    port map (
            O => \N__22528\,
            I => \N__22494\
        );

    \I__3574\ : Glb2LocalMux
    port map (
            O => \N__22525\,
            I => \N__22494\
        );

    \I__3573\ : Glb2LocalMux
    port map (
            O => \N__22522\,
            I => \N__22494\
        );

    \I__3572\ : Glb2LocalMux
    port map (
            O => \N__22519\,
            I => \N__22494\
        );

    \I__3571\ : GlobalMux
    port map (
            O => \N__22494\,
            I => \N__22491\
        );

    \I__3570\ : gio2CtrlBuf
    port map (
            O => \N__22491\,
            I => \b2v_inst200.count_en_g\
        );

    \I__3569\ : InMux
    port map (
            O => \N__22488\,
            I => \b2v_inst5.un2_count_1_cry_0\
        );

    \I__3568\ : InMux
    port map (
            O => \N__22485\,
            I => \b2v_inst5.un2_count_1_cry_1\
        );

    \I__3567\ : InMux
    port map (
            O => \N__22482\,
            I => \b2v_inst5.un2_count_1_cry_2\
        );

    \I__3566\ : InMux
    port map (
            O => \N__22479\,
            I => \b2v_inst5.un2_count_1_cry_3\
        );

    \I__3565\ : InMux
    port map (
            O => \N__22476\,
            I => \b2v_inst5.un2_count_1_cry_4\
        );

    \I__3564\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22467\
        );

    \I__3563\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22467\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__22467\,
            I => \b2v_inst200.count_3_15\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__3560\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22454\
        );

    \I__3558\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22451\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__22454\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__22451\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__3555\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22437\
        );

    \I__3554\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22437\
        );

    \I__3553\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22437\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__22434\,
            I => \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71\
        );

    \I__3550\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22426\
        );

    \I__3549\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22421\
        );

    \I__3548\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22421\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__22426\,
            I => \b2v_inst200.count_1_8\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__22421\,
            I => \b2v_inst200.count_1_8\
        );

    \I__3545\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22412\
        );

    \I__3544\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22409\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__22412\,
            I => \b2v_inst200.count_3_8\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__22409\,
            I => \b2v_inst200.count_3_8\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__22404\,
            I => \N__22400\
        );

    \I__3540\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22397\
        );

    \I__3539\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22394\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22391\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__22394\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__22391\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__3535\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22380\
        );

    \I__3533\ : Span4Mux_h
    port map (
            O => \N__22380\,
            I => \N__22377\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__22377\,
            I => \b2v_inst200.un25_clk_100khz_14\
        );

    \I__3531\ : InMux
    port map (
            O => \N__22374\,
            I => \N__22371\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__22371\,
            I => \b2v_inst200.un25_clk_100khz_6\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__22368\,
            I => \b2v_inst200.un25_clk_100khz_7_cascade_\
        );

    \I__3528\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22362\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__22362\,
            I => \N__22359\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__22359\,
            I => \b2v_inst200.un25_clk_100khz_13\
        );

    \I__3525\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22351\
        );

    \I__3524\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22348\
        );

    \I__3523\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22345\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__22351\,
            I => \N__22336\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__22348\,
            I => \N__22333\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__22345\,
            I => \N__22330\
        );

    \I__3519\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22325\
        );

    \I__3518\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22325\
        );

    \I__3517\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22320\
        );

    \I__3516\ : InMux
    port map (
            O => \N__22341\,
            I => \N__22320\
        );

    \I__3515\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22315\
        );

    \I__3514\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22315\
        );

    \I__3513\ : Span4Mux_v
    port map (
            O => \N__22336\,
            I => \N__22309\
        );

    \I__3512\ : Span4Mux_h
    port map (
            O => \N__22333\,
            I => \N__22309\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__22330\,
            I => \N__22300\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22300\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22300\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__22315\,
            I => \N__22300\
        );

    \I__3507\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22297\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__22309\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__22300\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__22297\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__22290\,
            I => \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_\
        );

    \I__3502\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22279\
        );

    \I__3501\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22276\
        );

    \I__3500\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22273\
        );

    \I__3499\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22266\
        );

    \I__3498\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22266\
        );

    \I__3497\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22266\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__22279\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__22276\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__22273\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__22266\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__3492\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__22254\,
            I => \b2v_inst200.count_3_0\
        );

    \I__3490\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22247\
        );

    \I__3489\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22244\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__22247\,
            I => \b2v_inst200.count_1_11\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__22244\,
            I => \b2v_inst200.count_1_11\
        );

    \I__3486\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__22236\,
            I => \N__22233\
        );

    \I__3484\ : Span4Mux_h
    port map (
            O => \N__22233\,
            I => \N__22230\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__22230\,
            I => \b2v_inst200.count_3_11\
        );

    \I__3482\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22223\
        );

    \I__3481\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22220\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__22223\,
            I => \N__22217\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__22220\,
            I => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__22217\,
            I => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\
        );

    \I__3477\ : InMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__22209\,
            I => \b2v_inst200.count_3_14\
        );

    \I__3475\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22202\
        );

    \I__3474\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22199\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22196\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__22199\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__22196\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__3470\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22188\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__22188\,
            I => \N__22185\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__22185\,
            I => \N__22182\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__22182\,
            I => \b2v_inst200.count_3_2\
        );

    \I__3466\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22175\
        );

    \I__3465\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22172\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22169\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__22172\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__22169\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__3461\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22161\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__22161\,
            I => \N__22158\
        );

    \I__3459\ : Span4Mux_v
    port map (
            O => \N__22158\,
            I => \N__22155\
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__22155\,
            I => \b2v_inst200.count_3_4\
        );

    \I__3457\ : InMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__22149\,
            I => \b2v_inst11.mult1_un89_sum_cry_5_s\
        );

    \I__3455\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__22143\,
            I => \N__22140\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__22140\,
            I => \b2v_inst11.mult1_un96_sum_cry_6_s\
        );

    \I__3452\ : InMux
    port map (
            O => \N__22137\,
            I => \b2v_inst11.mult1_un96_sum_cry_5\
        );

    \I__3451\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22131\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__22131\,
            I => \b2v_inst11.mult1_un89_sum_cry_6_s\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__3448\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__22119\,
            I => \b2v_inst11.mult1_un103_sum_axb_8\
        );

    \I__3445\ : InMux
    port map (
            O => \N__22116\,
            I => \b2v_inst11.mult1_un96_sum_cry_6\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__3443\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__22107\,
            I => \b2v_inst11.mult1_un96_sum_axb_8\
        );

    \I__3441\ : InMux
    port map (
            O => \N__22104\,
            I => \b2v_inst11.mult1_un96_sum_cry_7\
        );

    \I__3440\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22097\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__22100\,
            I => \N__22094\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22088\
        );

    \I__3437\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22081\
        );

    \I__3436\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22081\
        );

    \I__3435\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22081\
        );

    \I__3434\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22078\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__22088\,
            I => \N__22073\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__22081\,
            I => \N__22073\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__22078\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__22073\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__3429\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22064\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__22067\,
            I => \N__22060\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__22064\,
            I => \N__22055\
        );

    \I__3426\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22052\
        );

    \I__3425\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22045\
        );

    \I__3424\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22045\
        );

    \I__3423\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22045\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__22055\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__22052\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__22045\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__22038\,
            I => \N__22034\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__22037\,
            I => \N__22030\
        );

    \I__3417\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22023\
        );

    \I__3416\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22023\
        );

    \I__3415\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22023\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__22023\,
            I => \b2v_inst11.mult1_un89_sum_i_0_8\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__3412\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22014\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__22011\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__22011\,
            I => \b2v_inst200.un2_count_1_axb_15\
        );

    \I__3409\ : InMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__22005\,
            I => \b2v_inst200.un2_count_1_axb_8\
        );

    \I__3407\ : InMux
    port map (
            O => \N__22002\,
            I => \b2v_inst11.mult1_un89_sum_cry_4\
        );

    \I__3406\ : InMux
    port map (
            O => \N__21999\,
            I => \b2v_inst11.mult1_un89_sum_cry_5\
        );

    \I__3405\ : InMux
    port map (
            O => \N__21996\,
            I => \b2v_inst11.mult1_un89_sum_cry_6\
        );

    \I__3404\ : InMux
    port map (
            O => \N__21993\,
            I => \b2v_inst11.mult1_un89_sum_cry_7\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__21990\,
            I => \N__21986\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__21989\,
            I => \N__21982\
        );

    \I__3401\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21975\
        );

    \I__3400\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21975\
        );

    \I__3399\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21975\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__21975\,
            I => \b2v_inst11.mult1_un82_sum_i_0_8\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__21972\,
            I => \N__21969\
        );

    \I__3396\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21966\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21963\
        );

    \I__3394\ : Span4Mux_s2_h
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__21960\,
            I => \b2v_inst11.mult1_un96_sum_cry_3_s\
        );

    \I__3392\ : InMux
    port map (
            O => \N__21957\,
            I => \b2v_inst11.mult1_un96_sum_cry_2\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__21954\,
            I => \N__21951\
        );

    \I__3390\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__21948\,
            I => \b2v_inst11.mult1_un89_sum_cry_3_s\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__21945\,
            I => \N__21942\
        );

    \I__3387\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21939\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__21939\,
            I => \N__21936\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__21936\,
            I => \b2v_inst11.mult1_un96_sum_cry_4_s\
        );

    \I__3384\ : InMux
    port map (
            O => \N__21933\,
            I => \b2v_inst11.mult1_un96_sum_cry_3\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__3382\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21924\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__21924\,
            I => \b2v_inst11.mult1_un89_sum_cry_4_s\
        );

    \I__3380\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__21918\,
            I => \N__21915\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__21915\,
            I => \b2v_inst11.mult1_un96_sum_cry_5_s\
        );

    \I__3377\ : InMux
    port map (
            O => \N__21912\,
            I => \b2v_inst11.mult1_un96_sum_cry_4\
        );

    \I__3376\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21906\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__21900\,
            I => \b2v_inst11.mult1_un103_sum_cry_4_s\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__3371\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__21891\,
            I => \b2v_inst11.mult1_un110_sum_cry_5_s\
        );

    \I__3369\ : InMux
    port map (
            O => \N__21888\,
            I => \b2v_inst11.mult1_un110_sum_cry_4\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__21885\,
            I => \N__21881\
        );

    \I__3367\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21876\
        );

    \I__3366\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21876\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21872\
        );

    \I__3364\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21869\
        );

    \I__3363\ : Span4Mux_s3_v
    port map (
            O => \N__21872\,
            I => \N__21862\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21862\
        );

    \I__3361\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21859\
        );

    \I__3360\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21856\
        );

    \I__3359\ : Span4Mux_h
    port map (
            O => \N__21862\,
            I => \N__21853\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__21859\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__21856\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__21853\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__3354\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21840\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__21840\,
            I => \N__21837\
        );

    \I__3352\ : Span4Mux_v
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__21834\,
            I => \b2v_inst11.mult1_un103_sum_cry_5_s\
        );

    \I__3350\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__21828\,
            I => \b2v_inst11.mult1_un110_sum_cry_6_s\
        );

    \I__3348\ : InMux
    port map (
            O => \N__21825\,
            I => \b2v_inst11.mult1_un110_sum_cry_5\
        );

    \I__3347\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21819\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__21819\,
            I => \N__21816\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__21816\,
            I => \N__21813\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__21813\,
            I => \b2v_inst11.mult1_un103_sum_cry_6_s\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__21810\,
            I => \N__21806\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__21809\,
            I => \N__21802\
        );

    \I__3341\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21795\
        );

    \I__3340\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21795\
        );

    \I__3339\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21795\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__21795\,
            I => \b2v_inst11.mult1_un103_sum_i_0_8\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__21792\,
            I => \N__21789\
        );

    \I__3336\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21786\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__21786\,
            I => \b2v_inst11.mult1_un117_sum_axb_8\
        );

    \I__3334\ : InMux
    port map (
            O => \N__21783\,
            I => \b2v_inst11.mult1_un110_sum_cry_6\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__3332\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21774\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__3330\ : Span4Mux_h
    port map (
            O => \N__21771\,
            I => \N__21768\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__21768\,
            I => \b2v_inst11.mult1_un110_sum_axb_8\
        );

    \I__3328\ : InMux
    port map (
            O => \N__21765\,
            I => \b2v_inst11.mult1_un110_sum_cry_7\
        );

    \I__3327\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21758\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__21761\,
            I => \N__21754\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21750\
        );

    \I__3324\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21745\
        );

    \I__3323\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21745\
        );

    \I__3322\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21742\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__21750\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__21745\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__21742\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__21735\,
            I => \b2v_inst11.mult1_un110_sum_s_8_cascade_\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__21732\,
            I => \N__21728\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__21731\,
            I => \N__21724\
        );

    \I__3315\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21717\
        );

    \I__3314\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21717\
        );

    \I__3313\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21717\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__21717\,
            I => \b2v_inst11.mult1_un110_sum_i_0_8\
        );

    \I__3311\ : InMux
    port map (
            O => \N__21714\,
            I => \b2v_inst11.mult1_un89_sum_cry_2\
        );

    \I__3310\ : InMux
    port map (
            O => \N__21711\,
            I => \b2v_inst11.mult1_un89_sum_cry_3\
        );

    \I__3309\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21705\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__21705\,
            I => \b2v_inst11.mult1_un138_sum_i\
        );

    \I__3307\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21699\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__21699\,
            I => \N__21696\
        );

    \I__3305\ : Span4Mux_s1_v
    port map (
            O => \N__21696\,
            I => \N__21693\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__21693\,
            I => \b2v_inst11.mult1_un124_sum_i\
        );

    \I__3303\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21687\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__21687\,
            I => \b2v_inst11.mult1_un110_sum_i\
        );

    \I__3301\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21681\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__21681\,
            I => \b2v_inst11.mult1_un103_sum_i\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__3298\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21672\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__21672\,
            I => \b2v_inst11.mult1_un110_sum_cry_3_s\
        );

    \I__3296\ : InMux
    port map (
            O => \N__21669\,
            I => \b2v_inst11.mult1_un110_sum_cry_2\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__21666\,
            I => \N__21663\
        );

    \I__3294\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21660\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__21660\,
            I => \N__21657\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__21657\,
            I => \N__21654\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__21654\,
            I => \b2v_inst11.mult1_un103_sum_cry_3_s\
        );

    \I__3290\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21648\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__21648\,
            I => \b2v_inst11.mult1_un110_sum_cry_4_s\
        );

    \I__3288\ : InMux
    port map (
            O => \N__21645\,
            I => \b2v_inst11.mult1_un110_sum_cry_3\
        );

    \I__3287\ : InMux
    port map (
            O => \N__21642\,
            I => \bfn_5_12_0_\
        );

    \I__3286\ : InMux
    port map (
            O => \N__21639\,
            I => \b2v_inst20.counter_1_cry_25\
        );

    \I__3285\ : InMux
    port map (
            O => \N__21636\,
            I => \b2v_inst20.counter_1_cry_26\
        );

    \I__3284\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21629\
        );

    \I__3283\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21626\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__21629\,
            I => \N__21623\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__21626\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__3280\ : Odrv12
    port map (
            O => \N__21623\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__3279\ : InMux
    port map (
            O => \N__21618\,
            I => \b2v_inst20.counter_1_cry_27\
        );

    \I__3278\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21611\
        );

    \I__3277\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21608\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__21611\,
            I => \N__21605\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__21608\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__3274\ : Odrv12
    port map (
            O => \N__21605\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__3273\ : InMux
    port map (
            O => \N__21600\,
            I => \b2v_inst20.counter_1_cry_28\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__21597\,
            I => \N__21594\
        );

    \I__3271\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21590\
        );

    \I__3270\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21587\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__21590\,
            I => \N__21584\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__21587\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__3267\ : Odrv12
    port map (
            O => \N__21584\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__3266\ : InMux
    port map (
            O => \N__21579\,
            I => \b2v_inst20.counter_1_cry_29\
        );

    \I__3265\ : InMux
    port map (
            O => \N__21576\,
            I => \b2v_inst20.counter_1_cry_30\
        );

    \I__3264\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21569\
        );

    \I__3263\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21566\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21563\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__21566\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__3260\ : Odrv12
    port map (
            O => \N__21563\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__3259\ : InMux
    port map (
            O => \N__21558\,
            I => \bfn_5_11_0_\
        );

    \I__3258\ : InMux
    port map (
            O => \N__21555\,
            I => \b2v_inst20.counter_1_cry_17\
        );

    \I__3257\ : InMux
    port map (
            O => \N__21552\,
            I => \b2v_inst20.counter_1_cry_18\
        );

    \I__3256\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21545\
        );

    \I__3255\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21542\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__21545\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__21542\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__3252\ : InMux
    port map (
            O => \N__21537\,
            I => \b2v_inst20.counter_1_cry_19\
        );

    \I__3251\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21530\
        );

    \I__3250\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21527\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__21530\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__21527\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__3247\ : InMux
    port map (
            O => \N__21522\,
            I => \b2v_inst20.counter_1_cry_20\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__21519\,
            I => \N__21515\
        );

    \I__3245\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21512\
        );

    \I__3244\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21509\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__21512\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__21509\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__3241\ : InMux
    port map (
            O => \N__21504\,
            I => \b2v_inst20.counter_1_cry_21\
        );

    \I__3240\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21497\
        );

    \I__3239\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21494\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__21497\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__21494\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__3236\ : InMux
    port map (
            O => \N__21489\,
            I => \b2v_inst20.counter_1_cry_22\
        );

    \I__3235\ : InMux
    port map (
            O => \N__21486\,
            I => \b2v_inst20.counter_1_cry_23\
        );

    \I__3234\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21479\
        );

    \I__3233\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21476\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__21479\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__21476\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__3230\ : InMux
    port map (
            O => \N__21471\,
            I => \b2v_inst20.counter_1_cry_7\
        );

    \I__3229\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21464\
        );

    \I__3228\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21461\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__21464\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__21461\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__3225\ : InMux
    port map (
            O => \N__21456\,
            I => \bfn_5_10_0_\
        );

    \I__3224\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21449\
        );

    \I__3223\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21446\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__21449\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__21446\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__3220\ : InMux
    port map (
            O => \N__21441\,
            I => \b2v_inst20.counter_1_cry_9\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__21438\,
            I => \N__21434\
        );

    \I__3218\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21431\
        );

    \I__3217\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21428\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__21431\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__21428\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__3214\ : InMux
    port map (
            O => \N__21423\,
            I => \b2v_inst20.counter_1_cry_10\
        );

    \I__3213\ : InMux
    port map (
            O => \N__21420\,
            I => \b2v_inst20.counter_1_cry_11\
        );

    \I__3212\ : InMux
    port map (
            O => \N__21417\,
            I => \b2v_inst20.counter_1_cry_12\
        );

    \I__3211\ : InMux
    port map (
            O => \N__21414\,
            I => \b2v_inst20.counter_1_cry_13\
        );

    \I__3210\ : InMux
    port map (
            O => \N__21411\,
            I => \b2v_inst20.counter_1_cry_14\
        );

    \I__3209\ : InMux
    port map (
            O => \N__21408\,
            I => \b2v_inst20.counter_1_cry_15\
        );

    \I__3208\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21402\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__21402\,
            I => \b2v_inst200.HDA_SDO_ATP_0\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__21399\,
            I => \N__21396\
        );

    \I__3205\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21391\
        );

    \I__3204\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21386\
        );

    \I__3203\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21386\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__21391\,
            I => \b2v_inst200.N_205\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__21386\,
            I => \b2v_inst200.N_205\
        );

    \I__3200\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21372\
        );

    \I__3199\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21372\
        );

    \I__3198\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21372\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__21372\,
            I => \b2v_inst200.curr_state_i_2\
        );

    \I__3196\ : IoInMux
    port map (
            O => \N__21369\,
            I => \N__21366\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__3194\ : Odrv12
    port map (
            O => \N__21363\,
            I => hda_sdo_atp
        );

    \I__3193\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21351\
        );

    \I__3192\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21351\
        );

    \I__3191\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21351\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21347\
        );

    \I__3189\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21344\
        );

    \I__3188\ : Odrv12
    port map (
            O => \N__21347\,
            I => \b2v_inst200.N_282\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__21344\,
            I => \b2v_inst200.N_282\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__3185\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21332\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__21335\,
            I => \N__21329\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21325\
        );

    \I__3182\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21320\
        );

    \I__3181\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21320\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__21325\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__21320\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__3178\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21309\
        );

    \I__3177\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21309\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21304\
        );

    \I__3175\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21299\
        );

    \I__3174\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21299\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__21304\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__21299\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__3171\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21291\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__21291\,
            I => \N__21288\
        );

    \I__3169\ : Span4Mux_v
    port map (
            O => \N__21288\,
            I => \N__21285\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__21285\,
            I => \b2v_inst200.curr_state_3_1\
        );

    \I__3167\ : InMux
    port map (
            O => \N__21282\,
            I => \b2v_inst20.counter_1_cry_1\
        );

    \I__3166\ : InMux
    port map (
            O => \N__21279\,
            I => \b2v_inst20.counter_1_cry_2\
        );

    \I__3165\ : InMux
    port map (
            O => \N__21276\,
            I => \b2v_inst20.counter_1_cry_3\
        );

    \I__3164\ : InMux
    port map (
            O => \N__21273\,
            I => \b2v_inst20.counter_1_cry_4\
        );

    \I__3163\ : InMux
    port map (
            O => \N__21270\,
            I => \b2v_inst20.counter_1_cry_5\
        );

    \I__3162\ : InMux
    port map (
            O => \N__21267\,
            I => \b2v_inst20.counter_1_cry_6\
        );

    \I__3161\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21258\
        );

    \I__3160\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21258\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__21258\,
            I => \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\
        );

    \I__3158\ : InMux
    port map (
            O => \N__21255\,
            I => \b2v_inst11.un3_count_off_1_cry_13\
        );

    \I__3157\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21248\
        );

    \I__3156\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21245\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__21248\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__21245\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__3153\ : InMux
    port map (
            O => \N__21240\,
            I => \b2v_inst11.un3_count_off_1_cry_14\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__21237\,
            I => \N__21233\
        );

    \I__3151\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21228\
        );

    \I__3150\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21228\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__21228\,
            I => \b2v_inst11.count_offZ0Z_12\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__21225\,
            I => \N__21221\
        );

    \I__3147\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21216\
        );

    \I__3146\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21216\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__21216\,
            I => \b2v_inst11.count_offZ0Z_11\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__21213\,
            I => \N__21209\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__21212\,
            I => \N__21206\
        );

    \I__3142\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21201\
        );

    \I__3141\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21201\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__21201\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__21198\,
            I => \N__21194\
        );

    \I__3138\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21189\
        );

    \I__3137\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21189\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__21189\,
            I => \b2v_inst11.count_offZ0Z_9\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__21186\,
            I => \b2v_inst200.curr_state_i_2_cascade_\
        );

    \I__3134\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__21180\,
            I => \b2v_inst200.i4_mux\
        );

    \I__3132\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21173\
        );

    \I__3131\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21170\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__21173\,
            I => \N__21167\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__21170\,
            I => \b2v_inst200.N_2989_i\
        );

    \I__3128\ : Odrv12
    port map (
            O => \N__21167\,
            I => \b2v_inst200.N_2989_i\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__21162\,
            I => \b2v_inst200.N_205_cascade_\
        );

    \I__3126\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__21156\,
            I => \b2v_inst200.curr_stateZ0Z_2\
        );

    \I__3124\ : InMux
    port map (
            O => \N__21153\,
            I => \b2v_inst11.un3_count_off_1_cry_5\
        );

    \I__3123\ : InMux
    port map (
            O => \N__21150\,
            I => \b2v_inst11.un3_count_off_1_cry_6\
        );

    \I__3122\ : InMux
    port map (
            O => \N__21147\,
            I => \b2v_inst11.un3_count_off_1_cry_7\
        );

    \I__3121\ : InMux
    port map (
            O => \N__21144\,
            I => \bfn_5_7_0_\
        );

    \I__3120\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21137\
        );

    \I__3119\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21134\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__21137\,
            I => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__21134\,
            I => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\
        );

    \I__3116\ : InMux
    port map (
            O => \N__21129\,
            I => \b2v_inst11.un3_count_off_1_cry_9\
        );

    \I__3115\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21120\
        );

    \I__3114\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21120\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__21120\,
            I => \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\
        );

    \I__3112\ : InMux
    port map (
            O => \N__21117\,
            I => \b2v_inst11.un3_count_off_1_cry_10\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__3110\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21105\
        );

    \I__3109\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21105\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__21105\,
            I => \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\
        );

    \I__3107\ : InMux
    port map (
            O => \N__21102\,
            I => \b2v_inst11.un3_count_off_1_cry_11\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__21099\,
            I => \N__21095\
        );

    \I__3105\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21092\
        );

    \I__3104\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21089\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__21092\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__21089\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__3101\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21078\
        );

    \I__3100\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21078\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__21078\,
            I => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\
        );

    \I__3098\ : InMux
    port map (
            O => \N__21075\,
            I => \b2v_inst11.un3_count_off_1_cry_12\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__21072\,
            I => \N__21069\
        );

    \I__3096\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__21066\,
            I => \b2v_inst11.count_offZ0Z_14\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__21063\,
            I => \b2v_inst200.m6_i_0_cascade_\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__21060\,
            I => \b2v_inst200.N_58_cascade_\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__21057\,
            I => \b2v_inst200.curr_stateZ0Z_0_cascade_\
        );

    \I__3091\ : InMux
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21046\
        );

    \I__3089\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21043\
        );

    \I__3088\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21040\
        );

    \I__3087\ : Span4Mux_v
    port map (
            O => \N__21046\,
            I => \N__21037\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__21043\,
            I => \N_411\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N_411\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__21037\,
            I => \N_411\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__21030\,
            I => \N_411_cascade_\
        );

    \I__3082\ : InMux
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__21024\,
            I => \b2v_inst200.m6_i_0\
        );

    \I__3080\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21018\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__21018\,
            I => \b2v_inst200.curr_state_3_0\
        );

    \I__3078\ : InMux
    port map (
            O => \N__21015\,
            I => \b2v_inst11.un3_count_off_1_cry_1\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__21012\,
            I => \N__21008\
        );

    \I__3076\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21003\
        );

    \I__3075\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21003\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__21000\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__21000\,
            I => \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20997\,
            I => \b2v_inst11.un3_count_off_1_cry_2\
        );

    \I__3071\ : InMux
    port map (
            O => \N__20994\,
            I => \b2v_inst11.un3_count_off_1_cry_3\
        );

    \I__3070\ : InMux
    port map (
            O => \N__20991\,
            I => \b2v_inst11.un3_count_off_1_cry_4\
        );

    \I__3069\ : InMux
    port map (
            O => \N__20988\,
            I => \b2v_inst200.un2_count_1_cry_14\
        );

    \I__3068\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20982\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__20982\,
            I => \N__20979\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__20979\,
            I => \b2v_inst200.un2_count_1_axb_16\
        );

    \I__3065\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20967\
        );

    \I__3064\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20967\
        );

    \I__3063\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20967\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__20967\,
            I => \N__20964\
        );

    \I__3061\ : Span4Mux_s0_v
    port map (
            O => \N__20964\,
            I => \N__20961\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__20961\,
            I => \b2v_inst200.count_1_16\
        );

    \I__3059\ : InMux
    port map (
            O => \N__20958\,
            I => \b2v_inst200.un2_count_1_cry_15\
        );

    \I__3058\ : InMux
    port map (
            O => \N__20955\,
            I => \N__20951\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__20954\,
            I => \N__20948\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__20951\,
            I => \N__20945\
        );

    \I__3055\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20942\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__20945\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__20942\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__3052\ : InMux
    port map (
            O => \N__20937\,
            I => \bfn_5_4_0_\
        );

    \I__3051\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20930\
        );

    \I__3050\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20927\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__20930\,
            I => \N__20924\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__20927\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__20924\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__3046\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20916\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20913\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__20913\,
            I => \b2v_inst200.count_0_17\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__20910\,
            I => \b2v_inst200.N_56_cascade_\
        );

    \I__3042\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__20901\,
            I => \N__20898\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__20895\,
            I => gpio_fpga_soc_1
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__20892\,
            I => \b2v_inst200.curr_stateZ0Z_1_cascade_\
        );

    \I__3036\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20885\
        );

    \I__3035\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20882\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__20885\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__20882\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__3032\ : InMux
    port map (
            O => \N__20877\,
            I => \b2v_inst200.un2_count_1_cry_6\
        );

    \I__3031\ : InMux
    port map (
            O => \N__20874\,
            I => \b2v_inst200.un2_count_1_cry_7\
        );

    \I__3030\ : InMux
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__20868\,
            I => \b2v_inst200.un2_count_1_axb_9\
        );

    \I__3028\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20856\
        );

    \I__3027\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20856\
        );

    \I__3026\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20856\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__20856\,
            I => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\
        );

    \I__3024\ : InMux
    port map (
            O => \N__20853\,
            I => \bfn_5_3_0_\
        );

    \I__3023\ : InMux
    port map (
            O => \N__20850\,
            I => \b2v_inst200.un2_count_1_cry_9\
        );

    \I__3022\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__20844\,
            I => \N__20840\
        );

    \I__3020\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20837\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__20840\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__20837\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__3017\ : InMux
    port map (
            O => \N__20832\,
            I => \b2v_inst200.un2_count_1_cry_10\
        );

    \I__3016\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20826\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__20826\,
            I => \b2v_inst200.countZ0Z_12\
        );

    \I__3014\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20817\
        );

    \I__3013\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20817\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__20817\,
            I => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\
        );

    \I__3011\ : InMux
    port map (
            O => \N__20814\,
            I => \b2v_inst200.un2_count_1_cry_11\
        );

    \I__3010\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20808\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__20808\,
            I => \b2v_inst200.un2_count_1_axb_13\
        );

    \I__3008\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20796\
        );

    \I__3007\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20796\
        );

    \I__3006\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20796\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__20796\,
            I => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\
        );

    \I__3004\ : InMux
    port map (
            O => \N__20793\,
            I => \b2v_inst200.un2_count_1_cry_12\
        );

    \I__3003\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20786\
        );

    \I__3002\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20783\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20780\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__20783\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__20780\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__2998\ : InMux
    port map (
            O => \N__20775\,
            I => \b2v_inst200.un2_count_1_cry_13\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__20772\,
            I => \b2v_inst200.count_1_0_cascade_\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__20769\,
            I => \N__20765\
        );

    \I__2995\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20762\
        );

    \I__2994\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20759\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__20762\,
            I => \b2v_inst200.un2_count_1_axb_1\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__20759\,
            I => \b2v_inst200.un2_count_1_axb_1\
        );

    \I__2991\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20750\
        );

    \I__2990\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20747\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__20750\,
            I => \N__20744\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__20747\,
            I => \N__20741\
        );

    \I__2987\ : Odrv12
    port map (
            O => \N__20744\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__20741\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__2985\ : InMux
    port map (
            O => \N__20736\,
            I => \b2v_inst200.un2_count_1_cry_1\
        );

    \I__2984\ : InMux
    port map (
            O => \N__20733\,
            I => \N__20730\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__20730\,
            I => \b2v_inst200.un2_count_1_axb_3\
        );

    \I__2982\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20720\
        );

    \I__2981\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20720\
        );

    \I__2980\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20717\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__20720\,
            I => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__20717\,
            I => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\
        );

    \I__2977\ : InMux
    port map (
            O => \N__20712\,
            I => \b2v_inst200.un2_count_1_cry_2\
        );

    \I__2976\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20705\
        );

    \I__2975\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20697\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__20702\,
            I => \N__20697\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__20697\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__2971\ : InMux
    port map (
            O => \N__20694\,
            I => \b2v_inst200.un2_count_1_cry_3\
        );

    \I__2970\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__20688\,
            I => \b2v_inst200.un2_count_1_axb_5\
        );

    \I__2968\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20680\
        );

    \I__2967\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20675\
        );

    \I__2966\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20675\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__20680\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__20675\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__2963\ : InMux
    port map (
            O => \N__20670\,
            I => \b2v_inst200.un2_count_1_cry_4\
        );

    \I__2962\ : InMux
    port map (
            O => \N__20667\,
            I => \b2v_inst200.un2_count_1_cry_5_cZ0\
        );

    \I__2961\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__20661\,
            I => \b2v_inst11.mult1_un124_sum_cry_5_s\
        );

    \I__2959\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__20655\,
            I => \N__20652\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__20652\,
            I => \b2v_inst11.mult1_un131_sum_cry_6_s\
        );

    \I__2956\ : InMux
    port map (
            O => \N__20649\,
            I => \b2v_inst11.mult1_un131_sum_cry_5\
        );

    \I__2955\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__20643\,
            I => \b2v_inst11.mult1_un124_sum_cry_6_s\
        );

    \I__2953\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__20634\,
            I => \b2v_inst11.mult1_un138_sum_axb_8\
        );

    \I__2950\ : InMux
    port map (
            O => \N__20631\,
            I => \b2v_inst11.mult1_un131_sum_cry_6\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__20628\,
            I => \N__20625\
        );

    \I__2948\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__20622\,
            I => \b2v_inst11.mult1_un131_sum_axb_8\
        );

    \I__2946\ : InMux
    port map (
            O => \N__20619\,
            I => \b2v_inst11.mult1_un131_sum_cry_7\
        );

    \I__2945\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20612\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__20615\,
            I => \N__20609\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20604\
        );

    \I__2942\ : InMux
    port map (
            O => \N__20609\,
            I => \N__20596\
        );

    \I__2941\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20596\
        );

    \I__2940\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20596\
        );

    \I__2939\ : Span4Mux_s3_h
    port map (
            O => \N__20604\,
            I => \N__20593\
        );

    \I__2938\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20590\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__20596\,
            I => \N__20587\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__20593\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__20590\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__2934\ : Odrv12
    port map (
            O => \N__20587\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__2933\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20573\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__20576\,
            I => \N__20569\
        );

    \I__2930\ : Span4Mux_s3_h
    port map (
            O => \N__20573\,
            I => \N__20564\
        );

    \I__2929\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20561\
        );

    \I__2928\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20554\
        );

    \I__2927\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20554\
        );

    \I__2926\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20554\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__20564\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__20561\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__20554\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__20547\,
            I => \N__20543\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__20546\,
            I => \N__20539\
        );

    \I__2920\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20532\
        );

    \I__2919\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20532\
        );

    \I__2918\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20532\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__20532\,
            I => \b2v_inst11.mult1_un124_sum_i_0_8\
        );

    \I__2916\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20526\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__20520\,
            I => \N__20516\
        );

    \I__2912\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20513\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__20516\,
            I => \b2v_inst16.N_208_0\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__20513\,
            I => \b2v_inst16.N_208_0\
        );

    \I__2909\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20505\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20502\
        );

    \I__2907\ : Span12Mux_s8_h
    port map (
            O => \N__20502\,
            I => \N__20499\
        );

    \I__2906\ : Odrv12
    port map (
            O => \N__20499\,
            I => \b2v_inst16.delayed_vddq_pwrgd_en\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__20496\,
            I => \N__20493\
        );

    \I__2904\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20490\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__20490\,
            I => \N__20487\
        );

    \I__2902\ : Span4Mux_s0_v
    port map (
            O => \N__20487\,
            I => \N__20481\
        );

    \I__2901\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20478\
        );

    \I__2900\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20470\
        );

    \I__2899\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20470\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__20481\,
            I => \N__20465\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__20478\,
            I => \N__20465\
        );

    \I__2896\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20462\
        );

    \I__2895\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20457\
        );

    \I__2894\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20457\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20454\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__20465\,
            I => \N__20451\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__20462\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__20457\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__20454\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__20451\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__2887\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__2885\ : Span12Mux_s4_h
    port map (
            O => \N__20436\,
            I => \N__20432\
        );

    \I__2884\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20429\
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__20432\,
            I => \b2v_inst16.delayed_vddq_pwrgdZ0\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__20429\,
            I => \b2v_inst16.delayed_vddq_pwrgdZ0\
        );

    \I__2881\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20420\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__20423\,
            I => \N__20416\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__20420\,
            I => \N__20412\
        );

    \I__2878\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20407\
        );

    \I__2877\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20407\
        );

    \I__2876\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20404\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__20412\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__20407\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__20404\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20394\
        );

    \I__2871\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20391\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__20391\,
            I => \b2v_inst11.mult1_un117_sum_cry_5_s\
        );

    \I__2869\ : InMux
    port map (
            O => \N__20388\,
            I => \b2v_inst11.mult1_un124_sum_cry_5\
        );

    \I__2868\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__20382\,
            I => \b2v_inst11.mult1_un117_sum_cry_6_s\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__20379\,
            I => \N__20375\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__20378\,
            I => \N__20371\
        );

    \I__2864\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20364\
        );

    \I__2863\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20364\
        );

    \I__2862\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20364\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__20364\,
            I => \b2v_inst11.mult1_un117_sum_i_0_8\
        );

    \I__2860\ : InMux
    port map (
            O => \N__20361\,
            I => \b2v_inst11.mult1_un124_sum_cry_6\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__2858\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20352\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__20352\,
            I => \b2v_inst11.mult1_un124_sum_axb_8\
        );

    \I__2856\ : InMux
    port map (
            O => \N__20349\,
            I => \b2v_inst11.mult1_un124_sum_cry_7\
        );

    \I__2855\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__20343\,
            I => \b2v_inst11.mult1_un117_sum_i\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__20340\,
            I => \N__20337\
        );

    \I__2852\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20334\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__20334\,
            I => \N__20331\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__20331\,
            I => \b2v_inst11.mult1_un131_sum_cry_3_s\
        );

    \I__2849\ : InMux
    port map (
            O => \N__20328\,
            I => \b2v_inst11.mult1_un131_sum_cry_2\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20322\
        );

    \I__2847\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20319\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__20319\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \N__20313\
        );

    \I__2844\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__20307\,
            I => \b2v_inst11.mult1_un131_sum_cry_4_s\
        );

    \I__2841\ : InMux
    port map (
            O => \N__20304\,
            I => \b2v_inst11.mult1_un131_sum_cry_3\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__2839\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__20295\,
            I => \b2v_inst11.mult1_un124_sum_cry_4_s\
        );

    \I__2837\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20286\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__20286\,
            I => \b2v_inst11.mult1_un131_sum_cry_5_s\
        );

    \I__2834\ : InMux
    port map (
            O => \N__20283\,
            I => \b2v_inst11.mult1_un131_sum_cry_4\
        );

    \I__2833\ : InMux
    port map (
            O => \N__20280\,
            I => \b2v_inst11.mult1_un117_sum_cry_4\
        );

    \I__2832\ : InMux
    port map (
            O => \N__20277\,
            I => \b2v_inst11.mult1_un117_sum_cry_5\
        );

    \I__2831\ : InMux
    port map (
            O => \N__20274\,
            I => \b2v_inst11.mult1_un117_sum_cry_6\
        );

    \I__2830\ : InMux
    port map (
            O => \N__20271\,
            I => \b2v_inst11.mult1_un117_sum_cry_7\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__20268\,
            I => \b2v_inst11.mult1_un117_sum_s_8_cascade_\
        );

    \I__2828\ : InMux
    port map (
            O => \N__20265\,
            I => \b2v_inst11.mult1_un124_sum_cry_2\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__20262\,
            I => \N__20259\
        );

    \I__2826\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20256\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__20256\,
            I => \b2v_inst11.mult1_un117_sum_cry_3_s\
        );

    \I__2824\ : InMux
    port map (
            O => \N__20253\,
            I => \b2v_inst11.mult1_un124_sum_cry_3\
        );

    \I__2823\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20247\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__20247\,
            I => \b2v_inst11.mult1_un117_sum_cry_4_s\
        );

    \I__2821\ : InMux
    port map (
            O => \N__20244\,
            I => \b2v_inst11.mult1_un124_sum_cry_4\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__2819\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20235\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__20235\,
            I => \b2v_inst11.mult1_un138_sum_cry_4_s\
        );

    \I__2817\ : InMux
    port map (
            O => \N__20232\,
            I => \b2v_inst11.mult1_un138_sum_cry_3\
        );

    \I__2816\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__20226\,
            I => \b2v_inst11.mult1_un138_sum_cry_5_s\
        );

    \I__2814\ : InMux
    port map (
            O => \N__20223\,
            I => \b2v_inst11.mult1_un138_sum_cry_4\
        );

    \I__2813\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20217\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__20217\,
            I => \b2v_inst11.mult1_un138_sum_cry_6_s\
        );

    \I__2811\ : InMux
    port map (
            O => \N__20214\,
            I => \b2v_inst11.mult1_un138_sum_cry_5\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__2809\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20205\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__20205\,
            I => \b2v_inst11.mult1_un145_sum_axb_8\
        );

    \I__2807\ : InMux
    port map (
            O => \N__20202\,
            I => \b2v_inst11.mult1_un138_sum_cry_6\
        );

    \I__2806\ : InMux
    port map (
            O => \N__20199\,
            I => \b2v_inst11.mult1_un138_sum_cry_7\
        );

    \I__2805\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20189\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__20192\,
            I => \N__20185\
        );

    \I__2802\ : Span4Mux_s3_h
    port map (
            O => \N__20189\,
            I => \N__20180\
        );

    \I__2801\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20177\
        );

    \I__2800\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20170\
        );

    \I__2799\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20170\
        );

    \I__2798\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20170\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__20180\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__20177\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__20170\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__20163\,
            I => \N__20159\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__20162\,
            I => \N__20155\
        );

    \I__2792\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20148\
        );

    \I__2791\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20148\
        );

    \I__2790\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20148\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__20148\,
            I => \b2v_inst11.mult1_un131_sum_i_0_8\
        );

    \I__2788\ : InMux
    port map (
            O => \N__20145\,
            I => \b2v_inst11.mult1_un117_sum_cry_2\
        );

    \I__2787\ : InMux
    port map (
            O => \N__20142\,
            I => \b2v_inst11.mult1_un117_sum_cry_3\
        );

    \I__2786\ : InMux
    port map (
            O => \N__20139\,
            I => \b2v_inst11.mult1_un145_sum_cry_2\
        );

    \I__2785\ : InMux
    port map (
            O => \N__20136\,
            I => \b2v_inst11.mult1_un145_sum_cry_3\
        );

    \I__2784\ : InMux
    port map (
            O => \N__20133\,
            I => \b2v_inst11.mult1_un145_sum_cry_4\
        );

    \I__2783\ : InMux
    port map (
            O => \N__20130\,
            I => \b2v_inst11.mult1_un145_sum_cry_5\
        );

    \I__2782\ : InMux
    port map (
            O => \N__20127\,
            I => \b2v_inst11.mult1_un145_sum_cry_6\
        );

    \I__2781\ : InMux
    port map (
            O => \N__20124\,
            I => \b2v_inst11.mult1_un145_sum_cry_7\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__20121\,
            I => \N__20117\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__20120\,
            I => \N__20113\
        );

    \I__2778\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20106\
        );

    \I__2777\ : InMux
    port map (
            O => \N__20116\,
            I => \N__20106\
        );

    \I__2776\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20106\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__20106\,
            I => \b2v_inst11.mult1_un138_sum_i_0_8\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__20103\,
            I => \N__20100\
        );

    \I__2773\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20097\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__20097\,
            I => \b2v_inst11.mult1_un138_sum_cry_3_s\
        );

    \I__2771\ : InMux
    port map (
            O => \N__20094\,
            I => \b2v_inst11.mult1_un138_sum_cry_2\
        );

    \I__2770\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20088\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N__20081\
        );

    \I__2768\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20074\
        );

    \I__2767\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20074\
        );

    \I__2766\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20074\
        );

    \I__2765\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20071\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__20081\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__20074\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__20071\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__2761\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20043\
        );

    \I__2760\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20043\
        );

    \I__2759\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20043\
        );

    \I__2758\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20034\
        );

    \I__2757\ : InMux
    port map (
            O => \N__20060\,
            I => \N__20034\
        );

    \I__2756\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20034\
        );

    \I__2755\ : InMux
    port map (
            O => \N__20058\,
            I => \N__20034\
        );

    \I__2754\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20031\
        );

    \I__2753\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20022\
        );

    \I__2752\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20022\
        );

    \I__2751\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20022\
        );

    \I__2750\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20022\
        );

    \I__2749\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20015\
        );

    \I__2748\ : InMux
    port map (
            O => \N__20051\,
            I => \N__20015\
        );

    \I__2747\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20015\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__20007\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20007\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__20004\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__19999\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__19999\
        );

    \I__2741\ : InMux
    port map (
            O => \N__20014\,
            I => \N__19992\
        );

    \I__2740\ : InMux
    port map (
            O => \N__20013\,
            I => \N__19992\
        );

    \I__2739\ : InMux
    port map (
            O => \N__20012\,
            I => \N__19992\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__20007\,
            I => \N__19987\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__20004\,
            I => \N__19987\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__19999\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__19992\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__19987\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__2733\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__19974\,
            I => \b2v_inst11.count_1_0\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__19971\,
            I => \N__19967\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__19970\,
            I => \N__19963\
        );

    \I__2728\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19956\
        );

    \I__2727\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19956\
        );

    \I__2726\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19956\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__19956\,
            I => \G_2848\
        );

    \I__2724\ : InMux
    port map (
            O => \N__19953\,
            I => \b2v_inst11.mult1_un166_sum_cry_5\
        );

    \I__2723\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19945\
        );

    \I__2722\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19942\
        );

    \I__2721\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19939\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19936\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__19942\,
            I => \N__19933\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19930\
        );

    \I__2717\ : Span4Mux_s3_h
    port map (
            O => \N__19936\,
            I => \N__19925\
        );

    \I__2716\ : Span4Mux_s3_h
    port map (
            O => \N__19933\,
            I => \N__19925\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__19930\,
            I => \b2v_inst11.mult1_un166_sum_s_6\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__19925\,
            I => \b2v_inst11.mult1_un166_sum_s_6\
        );

    \I__2713\ : SRMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__19917\,
            I => \N__19914\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__19914\,
            I => \N__19911\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__19911\,
            I => \b2v_inst11.g0_0_0_rep1_1\
        );

    \I__2709\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19902\
        );

    \I__2708\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19902\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__19902\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__19899\,
            I => \N__19896\
        );

    \I__2705\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19890\
        );

    \I__2704\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19890\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__19890\,
            I => \N__19887\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__19887\,
            I => \b2v_inst11.g0_i_a3_0_1\
        );

    \I__2701\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19881\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__19881\,
            I => \b2v_inst11.N_6\
        );

    \I__2699\ : IoInMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__19875\,
            I => \N__19872\
        );

    \I__2697\ : IoSpan4Mux
    port map (
            O => \N__19872\,
            I => \N__19869\
        );

    \I__2696\ : IoSpan4Mux
    port map (
            O => \N__19869\,
            I => \N__19866\
        );

    \I__2695\ : Span4Mux_s2_h
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__19863\,
            I => pwrbtn_led
        );

    \I__2693\ : IoInMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__2691\ : Odrv12
    port map (
            O => \N__19854\,
            I => \b2v_inst200.count_enZ0\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__19851\,
            I => \b2v_inst16.delayed_vddq_pwrgd_en_cascade_\
        );

    \I__2689\ : IoInMux
    port map (
            O => \N__19848\,
            I => \N__19845\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__2687\ : Span4Mux_s1_h
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__2685\ : Sp12to4
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__2684\ : Odrv12
    port map (
            O => \N__19833\,
            I => vpp_en
        );

    \I__2683\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19826\
        );

    \I__2682\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19823\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__19826\,
            I => \N__19820\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__19823\,
            I => \b2v_inst16.curr_state_RNIBO6I1Z0Z_0\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__19820\,
            I => \b2v_inst16.curr_state_RNIBO6I1Z0Z_0\
        );

    \I__2678\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__19812\,
            I => \b2v_inst16.N_268\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__19809\,
            I => \b2v_inst16.N_268_cascade_\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__19806\,
            I => \N__19799\
        );

    \I__2674\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19786\
        );

    \I__2673\ : InMux
    port map (
            O => \N__19804\,
            I => \N__19786\
        );

    \I__2672\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19786\
        );

    \I__2671\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19786\
        );

    \I__2670\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19786\
        );

    \I__2669\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19783\
        );

    \I__2668\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19759\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19754\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__19783\,
            I => \N__19754\
        );

    \I__2665\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19749\
        );

    \I__2664\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19749\
        );

    \I__2663\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19746\
        );

    \I__2662\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19735\
        );

    \I__2661\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19735\
        );

    \I__2660\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19735\
        );

    \I__2659\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19735\
        );

    \I__2658\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19735\
        );

    \I__2657\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19726\
        );

    \I__2656\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19726\
        );

    \I__2655\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19726\
        );

    \I__2654\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19726\
        );

    \I__2653\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19715\
        );

    \I__2652\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19715\
        );

    \I__2651\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19715\
        );

    \I__2650\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19715\
        );

    \I__2649\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19715\
        );

    \I__2648\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19706\
        );

    \I__2647\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19706\
        );

    \I__2646\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19706\
        );

    \I__2645\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19706\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__19759\,
            I => \N__19701\
        );

    \I__2643\ : Span4Mux_s2_h
    port map (
            O => \N__19754\,
            I => \N__19701\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__19749\,
            I => \N__19698\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__19746\,
            I => \N__19695\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__19735\,
            I => \N__19692\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__19726\,
            I => \N__19689\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19684\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19684\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__19701\,
            I => \N__19681\
        );

    \I__2635\ : Span4Mux_s3_h
    port map (
            O => \N__19698\,
            I => \N__19676\
        );

    \I__2634\ : Span4Mux_s3_h
    port map (
            O => \N__19695\,
            I => \N__19676\
        );

    \I__2633\ : Span4Mux_s3_h
    port map (
            O => \N__19692\,
            I => \N__19671\
        );

    \I__2632\ : Span4Mux_s3_h
    port map (
            O => \N__19689\,
            I => \N__19671\
        );

    \I__2631\ : Span4Mux_s3_h
    port map (
            O => \N__19684\,
            I => \N__19668\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__19681\,
            I => \b2v_inst16.N_26\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__19676\,
            I => \b2v_inst16.N_26\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__19671\,
            I => \b2v_inst16.N_26\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__19668\,
            I => \b2v_inst16.N_26\
        );

    \I__2626\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__19656\,
            I => \b2v_inst11.count_off_0_3\
        );

    \I__2624\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19650\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__19650\,
            I => \N__19647\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__19647\,
            I => \b2v_inst11.count_off_0_14\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__19644\,
            I => \b2v_inst11.count_offZ0Z_14_cascade_\
        );

    \I__2620\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__19638\,
            I => \b2v_inst11.count_off_0_13\
        );

    \I__2618\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19629\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__19629\,
            I => \b2v_inst11.g0_i_o3_0\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__19626\,
            I => \N__19621\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__19625\,
            I => \N__19618\
        );

    \I__2613\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19613\
        );

    \I__2612\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19613\
        );

    \I__2611\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19610\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__19613\,
            I => \N__19605\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19605\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__19605\,
            I => \N__19602\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__19602\,
            I => \N__19599\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__19599\,
            I => \b2v_inst11.un85_clk_100khz1_THRU_CO\
        );

    \I__2605\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19591\
        );

    \I__2604\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19586\
        );

    \I__2603\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19586\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__19591\,
            I => \N__19583\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__19586\,
            I => \N__19580\
        );

    \I__2600\ : Span4Mux_v
    port map (
            O => \N__19583\,
            I => \N__19577\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__19580\,
            I => \N__19574\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__19577\,
            I => \N__19571\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__19574\,
            I => \b2v_inst11.un85_clk_100khz0_THRU_CO\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__19571\,
            I => \b2v_inst11.un85_clk_100khz0_THRU_CO\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__19566\,
            I => \b2v_inst11.N_6_cascade_\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \b2v_inst36.curr_stateZ0Z_0_cascade_\
        );

    \I__2593\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19550\
        );

    \I__2592\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19550\
        );

    \I__2591\ : SRMux
    port map (
            O => \N__19558\,
            I => \N__19550\
        );

    \I__2590\ : SRMux
    port map (
            O => \N__19557\,
            I => \N__19544\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__19550\,
            I => \N__19538\
        );

    \I__2588\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19531\
        );

    \I__2587\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19531\
        );

    \I__2586\ : SRMux
    port map (
            O => \N__19547\,
            I => \N__19531\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19527\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__19543\,
            I => \N__19521\
        );

    \I__2583\ : SRMux
    port map (
            O => \N__19542\,
            I => \N__19518\
        );

    \I__2582\ : SRMux
    port map (
            O => \N__19541\,
            I => \N__19515\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__19538\,
            I => \N__19510\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__19531\,
            I => \N__19510\
        );

    \I__2579\ : SRMux
    port map (
            O => \N__19530\,
            I => \N__19502\
        );

    \I__2578\ : Span4Mux_s1_h
    port map (
            O => \N__19527\,
            I => \N__19499\
        );

    \I__2577\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19492\
        );

    \I__2576\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19492\
        );

    \I__2575\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19492\
        );

    \I__2574\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19489\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__19518\,
            I => \N__19486\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19481\
        );

    \I__2571\ : Span4Mux_s1_v
    port map (
            O => \N__19510\,
            I => \N__19481\
        );

    \I__2570\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19472\
        );

    \I__2569\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19472\
        );

    \I__2568\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19472\
        );

    \I__2567\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19472\
        );

    \I__2566\ : SRMux
    port map (
            O => \N__19505\,
            I => \N__19464\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__19502\,
            I => \N__19453\
        );

    \I__2564\ : IoSpan4Mux
    port map (
            O => \N__19499\,
            I => \N__19446\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__19492\,
            I => \N__19446\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19446\
        );

    \I__2561\ : Span4Mux_v
    port map (
            O => \N__19486\,
            I => \N__19437\
        );

    \I__2560\ : Span4Mux_s1_h
    port map (
            O => \N__19481\,
            I => \N__19437\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__19472\,
            I => \N__19437\
        );

    \I__2558\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19434\
        );

    \I__2557\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19427\
        );

    \I__2556\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19427\
        );

    \I__2555\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19427\
        );

    \I__2554\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19424\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__19464\,
            I => \N__19421\
        );

    \I__2552\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19416\
        );

    \I__2551\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19416\
        );

    \I__2550\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19409\
        );

    \I__2549\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19409\
        );

    \I__2548\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19409\
        );

    \I__2547\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19402\
        );

    \I__2546\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19402\
        );

    \I__2545\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19402\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__19453\,
            I => \N__19397\
        );

    \I__2543\ : Span4Mux_s2_v
    port map (
            O => \N__19446\,
            I => \N__19397\
        );

    \I__2542\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19392\
        );

    \I__2541\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19392\
        );

    \I__2540\ : Sp12to4
    port map (
            O => \N__19437\,
            I => \N__19385\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19385\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__19427\,
            I => \N__19385\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__19424\,
            I => \N__19382\
        );

    \I__2536\ : IoSpan4Mux
    port map (
            O => \N__19421\,
            I => \N__19377\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__19416\,
            I => \N__19377\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19368\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__19402\,
            I => \N__19368\
        );

    \I__2532\ : IoSpan4Mux
    port map (
            O => \N__19397\,
            I => \N__19368\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__19392\,
            I => \N__19368\
        );

    \I__2530\ : Span12Mux_s5_v
    port map (
            O => \N__19385\,
            I => \N__19365\
        );

    \I__2529\ : Span4Mux_s3_h
    port map (
            O => \N__19382\,
            I => \N__19362\
        );

    \I__2528\ : Span4Mux_s3_h
    port map (
            O => \N__19377\,
            I => \N__19357\
        );

    \I__2527\ : Span4Mux_s3_h
    port map (
            O => \N__19368\,
            I => \N__19357\
        );

    \I__2526\ : Odrv12
    port map (
            O => \N__19365\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__19362\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__19357\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__2523\ : InMux
    port map (
            O => \N__19350\,
            I => \N__19347\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__19347\,
            I => \b2v_inst11.count_off_0_11\
        );

    \I__2521\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19341\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__19341\,
            I => \b2v_inst11.count_off_0_10\
        );

    \I__2519\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19335\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__19335\,
            I => \b2v_inst11.count_off_0_12\
        );

    \I__2517\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__19326\,
            I => \N__19322\
        );

    \I__2514\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19319\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__19322\,
            I => \b2v_inst16.count_rst_7\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__19319\,
            I => \b2v_inst16.count_rst_7\
        );

    \I__2511\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19311\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__19311\,
            I => \N__19308\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__19308\,
            I => \b2v_inst16.count_4_2\
        );

    \I__2508\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19301\
        );

    \I__2507\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19298\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19293\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N__19293\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__19293\,
            I => \N__19290\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__19290\,
            I => \b2v_inst16.count_rst_11\
        );

    \I__2502\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19284\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__19281\,
            I => \b2v_inst16.count_4_6\
        );

    \I__2499\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19266\
        );

    \I__2498\ : CEMux
    port map (
            O => \N__19277\,
            I => \N__19266\
        );

    \I__2497\ : CEMux
    port map (
            O => \N__19276\,
            I => \N__19263\
        );

    \I__2496\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19258\
        );

    \I__2495\ : CEMux
    port map (
            O => \N__19274\,
            I => \N__19258\
        );

    \I__2494\ : CEMux
    port map (
            O => \N__19273\,
            I => \N__19253\
        );

    \I__2493\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19248\
        );

    \I__2492\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19248\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__19266\,
            I => \N__19237\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__19263\,
            I => \N__19234\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__19258\,
            I => \N__19231\
        );

    \I__2488\ : CEMux
    port map (
            O => \N__19257\,
            I => \N__19228\
        );

    \I__2487\ : CEMux
    port map (
            O => \N__19256\,
            I => \N__19225\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19218\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19215\
        );

    \I__2484\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19210\
        );

    \I__2483\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19210\
        );

    \I__2482\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19207\
        );

    \I__2481\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19200\
        );

    \I__2480\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19200\
        );

    \I__2479\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19200\
        );

    \I__2478\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19195\
        );

    \I__2477\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19195\
        );

    \I__2476\ : Span4Mux_h
    port map (
            O => \N__19237\,
            I => \N__19190\
        );

    \I__2475\ : Span4Mux_s2_h
    port map (
            O => \N__19234\,
            I => \N__19190\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__19231\,
            I => \N__19185\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__19228\,
            I => \N__19185\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19182\
        );

    \I__2471\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19179\
        );

    \I__2470\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19172\
        );

    \I__2469\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19172\
        );

    \I__2468\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19172\
        );

    \I__2467\ : Span4Mux_s1_h
    port map (
            O => \N__19218\,
            I => \N__19159\
        );

    \I__2466\ : Span4Mux_h
    port map (
            O => \N__19215\,
            I => \N__19159\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__19210\,
            I => \N__19159\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19159\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19159\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__19195\,
            I => \N__19159\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__19190\,
            I => \b2v_inst16.count_en\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__19185\,
            I => \b2v_inst16.count_en\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__19182\,
            I => \b2v_inst16.count_en\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__19179\,
            I => \b2v_inst16.count_en\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__19172\,
            I => \b2v_inst16.count_en\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__19159\,
            I => \b2v_inst16.count_en\
        );

    \I__2455\ : SRMux
    port map (
            O => \N__19146\,
            I => \N__19142\
        );

    \I__2454\ : SRMux
    port map (
            O => \N__19145\,
            I => \N__19138\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19134\
        );

    \I__2452\ : SRMux
    port map (
            O => \N__19141\,
            I => \N__19131\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__19138\,
            I => \N__19127\
        );

    \I__2450\ : SRMux
    port map (
            O => \N__19137\,
            I => \N__19124\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__19134\,
            I => \N__19120\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__19131\,
            I => \N__19117\
        );

    \I__2447\ : SRMux
    port map (
            O => \N__19130\,
            I => \N__19114\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__19127\,
            I => \N__19109\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19109\
        );

    \I__2444\ : SRMux
    port map (
            O => \N__19123\,
            I => \N__19106\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__19120\,
            I => \b2v_inst16.N_3037_i\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__19117\,
            I => \b2v_inst16.N_3037_i\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__19114\,
            I => \b2v_inst16.N_3037_i\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__19109\,
            I => \b2v_inst16.N_3037_i\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__19106\,
            I => \b2v_inst16.N_3037_i\
        );

    \I__2438\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19092\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__19092\,
            I => \b2v_inst36.curr_state_0_1\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__19089\,
            I => \b2v_inst36.curr_state_7_1_cascade_\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__19086\,
            I => \b2v_inst36.curr_stateZ0Z_1_cascade_\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__19083\,
            I => \N__19077\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__19082\,
            I => \N__19074\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__19081\,
            I => \N__19065\
        );

    \I__2431\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19057\
        );

    \I__2430\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19054\
        );

    \I__2429\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19049\
        );

    \I__2428\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19049\
        );

    \I__2427\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19044\
        );

    \I__2426\ : InMux
    port map (
            O => \N__19071\,
            I => \N__19044\
        );

    \I__2425\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19037\
        );

    \I__2424\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19037\
        );

    \I__2423\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19037\
        );

    \I__2422\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19026\
        );

    \I__2421\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19026\
        );

    \I__2420\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19026\
        );

    \I__2419\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19026\
        );

    \I__2418\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19026\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__19060\,
            I => \N__19022\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__19057\,
            I => \N__19014\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__19054\,
            I => \N__19014\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__19049\,
            I => \N__19009\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19009\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19004\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__19026\,
            I => \N__19004\
        );

    \I__2410\ : InMux
    port map (
            O => \N__19025\,
            I => \N__18993\
        );

    \I__2409\ : InMux
    port map (
            O => \N__19022\,
            I => \N__18993\
        );

    \I__2408\ : InMux
    port map (
            O => \N__19021\,
            I => \N__18993\
        );

    \I__2407\ : InMux
    port map (
            O => \N__19020\,
            I => \N__18993\
        );

    \I__2406\ : InMux
    port map (
            O => \N__19019\,
            I => \N__18993\
        );

    \I__2405\ : Span4Mux_s1_v
    port map (
            O => \N__19014\,
            I => \N__18988\
        );

    \I__2404\ : Span4Mux_h
    port map (
            O => \N__19009\,
            I => \N__18988\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__19004\,
            I => \b2v_inst36.N_1_i\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__18993\,
            I => \b2v_inst36.N_1_i\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__18988\,
            I => \b2v_inst36.N_1_i\
        );

    \I__2400\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__18978\,
            I => \b2v_inst36.curr_state_0_0\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__18975\,
            I => \b2v_inst36.curr_state_7_0_cascade_\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__18972\,
            I => \N__18969\
        );

    \I__2396\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18965\
        );

    \I__2395\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18962\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__18965\,
            I => \b2v_inst200.count_3_5\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__18962\,
            I => \b2v_inst200.count_3_5\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__18957\,
            I => \N__18953\
        );

    \I__2391\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18950\
        );

    \I__2390\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18947\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__18950\,
            I => \N__18942\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18942\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__18942\,
            I => \N__18939\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__18939\,
            I => \b2v_inst16.countZ0Z_15\
        );

    \I__2385\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18930\
        );

    \I__2384\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18930\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__18930\,
            I => \N__18927\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__18927\,
            I => \N__18924\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__18924\,
            I => \b2v_inst16.count_rst_4\
        );

    \I__2380\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18918\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__18918\,
            I => \b2v_inst16.count_4_15\
        );

    \I__2378\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18912\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18908\
        );

    \I__2376\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18905\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__18908\,
            I => \N__18900\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__18905\,
            I => \N__18900\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__18900\,
            I => \N__18897\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__18897\,
            I => \b2v_inst16.countZ0Z_13\
        );

    \I__2371\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18888\
        );

    \I__2370\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18888\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__18888\,
            I => \N__18885\
        );

    \I__2368\ : Span4Mux_v
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__2367\ : Sp12to4
    port map (
            O => \N__18882\,
            I => \N__18879\
        );

    \I__2366\ : Odrv12
    port map (
            O => \N__18879\,
            I => \b2v_inst16.count_rst_2\
        );

    \I__2365\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18873\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__18873\,
            I => \b2v_inst16.count_4_13\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__18870\,
            I => \N__18867\
        );

    \I__2362\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18863\
        );

    \I__2361\ : InMux
    port map (
            O => \N__18866\,
            I => \N__18860\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__18863\,
            I => \N__18857\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18854\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__18857\,
            I => \N__18851\
        );

    \I__2357\ : Span4Mux_s3_h
    port map (
            O => \N__18854\,
            I => \N__18848\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__18851\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__18848\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__2354\ : InMux
    port map (
            O => \N__18843\,
            I => \N__18837\
        );

    \I__2353\ : InMux
    port map (
            O => \N__18842\,
            I => \N__18837\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__18837\,
            I => \N__18834\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__18834\,
            I => \N__18831\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__18831\,
            I => \b2v_inst16.count_rst_3\
        );

    \I__2349\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__18825\,
            I => \b2v_inst16.count_4_14\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__2346\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18813\
        );

    \I__2345\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18813\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__18813\,
            I => \b2v_inst200.count_3_3\
        );

    \I__2343\ : InMux
    port map (
            O => \N__18810\,
            I => \N__18807\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__18807\,
            I => \b2v_inst200.un25_clk_100khz_2\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__18804\,
            I => \N__18801\
        );

    \I__2340\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18795\
        );

    \I__2339\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18795\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__18795\,
            I => \b2v_inst200.count_3_13\
        );

    \I__2337\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18789\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__18789\,
            I => \b2v_inst200.un25_clk_100khz_5\
        );

    \I__2335\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__18783\,
            I => \b2v_inst200.count_3_12\
        );

    \I__2333\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18774\
        );

    \I__2332\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18774\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__18774\,
            I => \b2v_inst200.count_3_9\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__18771\,
            I => \b2v_inst200.countZ0Z_12_cascade_\
        );

    \I__2329\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__18765\,
            I => \b2v_inst200.un25_clk_100khz_4\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__18762\,
            I => \b2v_inst200.un25_clk_100khz_1_cascade_\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__18759\,
            I => \b2v_inst200.un2_count_1_axb_1_cascade_\
        );

    \I__2325\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18752\
        );

    \I__2324\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18749\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__18752\,
            I => \b2v_inst200.count_RNIZ0Z_1\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__18749\,
            I => \b2v_inst200.count_RNIZ0Z_1\
        );

    \I__2321\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18738\
        );

    \I__2320\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18738\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__18738\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__2318\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18732\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__18732\,
            I => \b2v_inst200.un25_clk_100khz_0\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__18729\,
            I => \N__18726\
        );

    \I__2315\ : InMux
    port map (
            O => \N__18726\,
            I => \N__18720\
        );

    \I__2314\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18720\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__18720\,
            I => \b2v_inst200.count_3_1\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__18717\,
            I => \b2v_inst200.un25_clk_100khz_3_cascade_\
        );

    \I__2311\ : InMux
    port map (
            O => \N__18714\,
            I => \b2v_inst11.mult1_un103_sum_cry_3\
        );

    \I__2310\ : InMux
    port map (
            O => \N__18711\,
            I => \b2v_inst11.mult1_un103_sum_cry_4\
        );

    \I__2309\ : InMux
    port map (
            O => \N__18708\,
            I => \b2v_inst11.mult1_un103_sum_cry_5\
        );

    \I__2308\ : InMux
    port map (
            O => \N__18705\,
            I => \b2v_inst11.mult1_un103_sum_cry_6\
        );

    \I__2307\ : InMux
    port map (
            O => \N__18702\,
            I => \b2v_inst11.mult1_un103_sum_cry_7\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__18699\,
            I => \N__18695\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__18698\,
            I => \N__18691\
        );

    \I__2304\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18684\
        );

    \I__2303\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18684\
        );

    \I__2302\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18684\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__18684\,
            I => \b2v_inst11.mult1_un96_sum_i_0_8\
        );

    \I__2300\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18677\
        );

    \I__2299\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18674\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__18677\,
            I => \b2v_inst11.N_5862_i\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__18674\,
            I => \b2v_inst11.N_5862_i\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__18669\,
            I => \N__18665\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__18668\,
            I => \N__18662\
        );

    \I__2294\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18659\
        );

    \I__2293\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18656\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__18659\,
            I => \N__18653\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__18656\,
            I => \b2v_inst11.un85_clk_100khz_1_8\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__18653\,
            I => \b2v_inst11.un85_clk_100khz_1_8\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__18648\,
            I => \N__18645\
        );

    \I__2288\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18641\
        );

    \I__2287\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18638\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__18641\,
            I => \b2v_inst11.N_5863_i\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__18638\,
            I => \b2v_inst11.N_5863_i\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__2283\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18626\
        );

    \I__2282\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18623\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__18626\,
            I => \N__18620\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__18623\,
            I => \b2v_inst11.un85_clk_100khz_1_9\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__18620\,
            I => \b2v_inst11.un85_clk_100khz_1_9\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__2277\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18608\
        );

    \I__2276\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18605\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__18608\,
            I => \b2v_inst11.N_5864_i\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__18605\,
            I => \b2v_inst11.N_5864_i\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__18600\,
            I => \N__18596\
        );

    \I__2272\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18593\
        );

    \I__2271\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18590\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__18593\,
            I => \b2v_inst11.un85_clk_100khz_1_10\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__18590\,
            I => \b2v_inst11.un85_clk_100khz_1_10\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__18585\,
            I => \N__18581\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__18584\,
            I => \N__18578\
        );

    \I__2266\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18575\
        );

    \I__2265\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18572\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__18575\,
            I => \b2v_inst11.N_5865_i\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__18572\,
            I => \b2v_inst11.N_5865_i\
        );

    \I__2262\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18563\
        );

    \I__2261\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18560\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18557\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__18560\,
            I => \b2v_inst11.un85_clk_100khz_1_11\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__18557\,
            I => \b2v_inst11.un85_clk_100khz_1_11\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__18552\,
            I => \N__18548\
        );

    \I__2256\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18545\
        );

    \I__2255\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18542\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__18545\,
            I => \b2v_inst11.N_5866_i\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__18542\,
            I => \b2v_inst11.N_5866_i\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__18537\,
            I => \N__18534\
        );

    \I__2251\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18530\
        );

    \I__2250\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18527\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__18530\,
            I => \b2v_inst11.un85_clk_100khz_1_12\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__18527\,
            I => \b2v_inst11.un85_clk_100khz_1_12\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__18522\,
            I => \N__18518\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__18521\,
            I => \N__18515\
        );

    \I__2245\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18512\
        );

    \I__2244\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18509\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__18512\,
            I => \b2v_inst11.N_5867_i\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__18509\,
            I => \b2v_inst11.N_5867_i\
        );

    \I__2241\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18500\
        );

    \I__2240\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18497\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__18500\,
            I => \b2v_inst11.un85_clk_100khz_1_13\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__18497\,
            I => \b2v_inst11.un85_clk_100khz_1_13\
        );

    \I__2237\ : InMux
    port map (
            O => \N__18492\,
            I => \b2v_inst11.un85_clk_100khz1\
        );

    \I__2236\ : InMux
    port map (
            O => \N__18489\,
            I => \b2v_inst11.mult1_un103_sum_cry_2\
        );

    \I__2235\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18482\
        );

    \I__2234\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18479\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__18482\,
            I => \b2v_inst11.N_5855_i\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__18479\,
            I => \b2v_inst11.N_5855_i\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__18474\,
            I => \N__18470\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__18473\,
            I => \N__18467\
        );

    \I__2229\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18464\
        );

    \I__2228\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18461\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__18464\,
            I => \b2v_inst11.un85_clk_100khz_0_1\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__18461\,
            I => \b2v_inst11.un85_clk_100khz_0_1\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__18456\,
            I => \N__18452\
        );

    \I__2224\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18449\
        );

    \I__2223\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18446\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__18449\,
            I => \b2v_inst11.N_5856_i\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__18446\,
            I => \b2v_inst11.N_5856_i\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__18441\,
            I => \N__18438\
        );

    \I__2219\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18434\
        );

    \I__2218\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18431\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__18434\,
            I => \b2v_inst11.un85_clk_100khz_0_2\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__18431\,
            I => \b2v_inst11.un85_clk_100khz_0_2\
        );

    \I__2215\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18422\
        );

    \I__2214\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18419\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__18422\,
            I => \b2v_inst11.N_5857_i\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__18419\,
            I => \b2v_inst11.N_5857_i\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__18414\,
            I => \N__18410\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__18413\,
            I => \N__18407\
        );

    \I__2209\ : InMux
    port map (
            O => \N__18410\,
            I => \N__18404\
        );

    \I__2208\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18401\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18398\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__18401\,
            I => \b2v_inst11.un85_clk_100khz_0_3\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__18398\,
            I => \b2v_inst11.un85_clk_100khz_0_3\
        );

    \I__2204\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18389\
        );

    \I__2203\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18386\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__18389\,
            I => \b2v_inst11.N_5858_i\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__18386\,
            I => \b2v_inst11.N_5858_i\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__18381\,
            I => \N__18377\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__18380\,
            I => \N__18374\
        );

    \I__2198\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__2197\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18368\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__18371\,
            I => \b2v_inst11.un85_clk_100khz_0_4\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__18368\,
            I => \b2v_inst11.un85_clk_100khz_0_4\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__2193\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18356\
        );

    \I__2192\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__18356\,
            I => \b2v_inst11.N_5859_i\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__18353\,
            I => \b2v_inst11.N_5859_i\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__18348\,
            I => \N__18344\
        );

    \I__2188\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18341\
        );

    \I__2187\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18338\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__18341\,
            I => \b2v_inst11.un85_clk_100khz_0_5\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__18338\,
            I => \b2v_inst11.un85_clk_100khz_0_5\
        );

    \I__2184\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18329\
        );

    \I__2183\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18326\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__18329\,
            I => \b2v_inst11.N_5860_i\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__18326\,
            I => \b2v_inst11.N_5860_i\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__18321\,
            I => \N__18317\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__18320\,
            I => \N__18314\
        );

    \I__2178\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18311\
        );

    \I__2177\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18308\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__18311\,
            I => \b2v_inst11.un85_clk_100khz_0_6\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__18308\,
            I => \b2v_inst11.un85_clk_100khz_0_6\
        );

    \I__2174\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18299\
        );

    \I__2173\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18296\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__18299\,
            I => \b2v_inst11.N_5861_i\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__18296\,
            I => \b2v_inst11.N_5861_i\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__18291\,
            I => \N__18287\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__18290\,
            I => \N__18284\
        );

    \I__2168\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18281\
        );

    \I__2167\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18278\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__18281\,
            I => \N__18275\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__18278\,
            I => \b2v_inst11.un85_clk_100khz_0_7\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__18275\,
            I => \b2v_inst11.un85_clk_100khz_0_7\
        );

    \I__2163\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18266\
        );

    \I__2162\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18263\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__18266\,
            I => \N__18259\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__18263\,
            I => \N__18256\
        );

    \I__2159\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18253\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__18259\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__18256\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__18253\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__2155\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18241\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__18245\,
            I => \N__18238\
        );

    \I__2153\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18235\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__18241\,
            I => \N__18232\
        );

    \I__2151\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18229\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__18235\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__18232\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__18229\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__2147\ : InMux
    port map (
            O => \N__18222\,
            I => \N__18217\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__18221\,
            I => \N__18214\
        );

    \I__2145\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18211\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18208\
        );

    \I__2143\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18205\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__18211\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__18208\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__18205\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__2139\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18193\
        );

    \I__2138\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18190\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__18196\,
            I => \N__18187\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__18193\,
            I => \N__18184\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__18190\,
            I => \N__18181\
        );

    \I__2134\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18178\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__18184\,
            I => \N__18175\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__18181\,
            I => \N__18170\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__18178\,
            I => \N__18170\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__18175\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__18170\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__18165\,
            I => \N__18162\
        );

    \I__2127\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18157\
        );

    \I__2126\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18154\
        );

    \I__2125\ : InMux
    port map (
            O => \N__18160\,
            I => \N__18151\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__18157\,
            I => \N__18148\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__18154\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__18151\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__18148\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__18141\,
            I => \b2v_inst11.un79_clk_100khzlt6_cascade_\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__18138\,
            I => \N__18134\
        );

    \I__2118\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18131\
        );

    \I__2117\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18127\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__18131\,
            I => \N__18124\
        );

    \I__2115\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18121\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__18127\,
            I => \N__18118\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__18124\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__18121\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__18118\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__2110\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18107\
        );

    \I__2109\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18103\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__18107\,
            I => \N__18100\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18097\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__18103\,
            I => \N__18094\
        );

    \I__2105\ : Span4Mux_s2_v
    port map (
            O => \N__18100\,
            I => \N__18091\
        );

    \I__2104\ : InMux
    port map (
            O => \N__18097\,
            I => \N__18088\
        );

    \I__2103\ : Odrv12
    port map (
            O => \N__18094\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__18091\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__18088\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__2100\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18078\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__18078\,
            I => \N__18073\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18070\
        );

    \I__2097\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18067\
        );

    \I__2096\ : Span4Mux_s2_v
    port map (
            O => \N__18073\,
            I => \N__18064\
        );

    \I__2095\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18061\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__18067\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__18064\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__18061\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__18054\,
            I => \N__18050\
        );

    \I__2090\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18047\
        );

    \I__2089\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18043\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__18047\,
            I => \N__18040\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__18046\,
            I => \N__18037\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__18032\
        );

    \I__2085\ : Span4Mux_s2_v
    port map (
            O => \N__18040\,
            I => \N__18032\
        );

    \I__2084\ : InMux
    port map (
            O => \N__18037\,
            I => \N__18029\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__18032\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__18029\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__2081\ : InMux
    port map (
            O => \N__18024\,
            I => \N__18019\
        );

    \I__2080\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18016\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__18013\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__18019\,
            I => \N__18008\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__18016\,
            I => \N__18008\
        );

    \I__2076\ : InMux
    port map (
            O => \N__18013\,
            I => \N__18005\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__18008\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__18005\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__2073\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17995\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__17999\,
            I => \N__17992\
        );

    \I__2071\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17989\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__17995\,
            I => \N__17986\
        );

    \I__2069\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17983\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__17989\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__17986\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__17983\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__17976\,
            I => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\
        );

    \I__2064\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17968\
        );

    \I__2063\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17965\
        );

    \I__2062\ : InMux
    port map (
            O => \N__17971\,
            I => \N__17962\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__17968\,
            I => \N__17959\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__17965\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__17962\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__17959\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__2057\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17949\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__17949\,
            I => \b2v_inst11.un79_clk_100khzlto15_3\
        );

    \I__2055\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17942\
        );

    \I__2054\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17938\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__17942\,
            I => \N__17935\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__17941\,
            I => \N__17932\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__17938\,
            I => \N__17927\
        );

    \I__2050\ : Span4Mux_s3_v
    port map (
            O => \N__17935\,
            I => \N__17927\
        );

    \I__2049\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17924\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__17927\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__17924\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__17919\,
            I => \b2v_inst11.un79_clk_100khzlto15_7_cascade_\
        );

    \I__2045\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17912\
        );

    \I__2044\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17908\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17905\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__17911\,
            I => \N__17902\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__17908\,
            I => \N__17899\
        );

    \I__2040\ : Span4Mux_s3_v
    port map (
            O => \N__17905\,
            I => \N__17896\
        );

    \I__2039\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17893\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__17899\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__17896\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__17893\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__17886\,
            I => \N__17881\
        );

    \I__2034\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17871\
        );

    \I__2033\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17871\
        );

    \I__2032\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17871\
        );

    \I__2031\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17871\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__2029\ : Odrv12
    port map (
            O => \N__17868\,
            I => \b2v_inst11.count_RNIZ0Z_8\
        );

    \I__2028\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17861\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__17864\,
            I => \N__17856\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17851\
        );

    \I__2025\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17848\
        );

    \I__2024\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17839\
        );

    \I__2023\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17839\
        );

    \I__2022\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17839\
        );

    \I__2021\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17839\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__17851\,
            I => \N__17836\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__17848\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__17839\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__17836\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__17829\,
            I => \b2v_inst11.count_RNIZ0Z_8_cascade_\
        );

    \I__2015\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17823\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__17823\,
            I => \N__17820\
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__17820\,
            I => \b2v_inst11.curr_state_3_i_m2_0_rep1_1\
        );

    \I__2012\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17813\
        );

    \I__2011\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17810\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__17813\,
            I => \b2v_inst11.N_5853_i\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__17810\,
            I => \b2v_inst11.N_5853_i\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__17805\,
            I => \N__17801\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__17804\,
            I => \N__17798\
        );

    \I__2006\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17795\
        );

    \I__2005\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17792\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__17795\,
            I => \b2v_inst11.un85_clk_100khz_0\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__17792\,
            I => \b2v_inst11.un85_clk_100khz_0\
        );

    \I__2002\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17783\
        );

    \I__2001\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17780\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__17783\,
            I => \b2v_inst11.N_5854_i\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__17780\,
            I => \b2v_inst11.N_5854_i\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__17775\,
            I => \N__17771\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__17774\,
            I => \N__17768\
        );

    \I__1996\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17765\
        );

    \I__1995\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17762\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__17765\,
            I => \N__17759\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__17762\,
            I => \b2v_inst11.un85_clk_100khz_0_0\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__17759\,
            I => \b2v_inst11.un85_clk_100khz_0_0\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__17754\,
            I => \N__17750\
        );

    \I__1990\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17745\
        );

    \I__1989\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17745\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__17745\,
            I => \b2v_inst11.count_1_2\
        );

    \I__1987\ : InMux
    port map (
            O => \N__17742\,
            I => \N__17739\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__17739\,
            I => \b2v_inst11.count_0_2\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__17736\,
            I => \N__17733\
        );

    \I__1984\ : InMux
    port map (
            O => \N__17733\,
            I => \N__17727\
        );

    \I__1983\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17727\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__17727\,
            I => \b2v_inst11.count_1_12\
        );

    \I__1981\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17721\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__17721\,
            I => \b2v_inst11.count_0_12\
        );

    \I__1979\ : InMux
    port map (
            O => \N__17718\,
            I => \N__17712\
        );

    \I__1978\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17712\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__17712\,
            I => \b2v_inst11.count_1_3\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__17709\,
            I => \N__17706\
        );

    \I__1975\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17703\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__17703\,
            I => \b2v_inst11.count_0_3\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__17700\,
            I => \N__17697\
        );

    \I__1972\ : InMux
    port map (
            O => \N__17697\,
            I => \N__17691\
        );

    \I__1971\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17691\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__17691\,
            I => \b2v_inst11.count_1_13\
        );

    \I__1969\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17685\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__17685\,
            I => \b2v_inst11.count_0_13\
        );

    \I__1967\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17676\
        );

    \I__1966\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17676\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__17676\,
            I => \b2v_inst11.count_1_4\
        );

    \I__1964\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17670\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__17670\,
            I => \b2v_inst11.count_0_4\
        );

    \I__1962\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17664\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__17664\,
            I => \N__17658\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__17663\,
            I => \N__17655\
        );

    \I__1959\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17650\
        );

    \I__1958\ : InMux
    port map (
            O => \N__17661\,
            I => \N__17650\
        );

    \I__1957\ : Span4Mux_s3_v
    port map (
            O => \N__17658\,
            I => \N__17647\
        );

    \I__1956\ : InMux
    port map (
            O => \N__17655\,
            I => \N__17644\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__17650\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__17647\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__17644\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__1952\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17634\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__17634\,
            I => \b2v_inst11.count_0_1\
        );

    \I__1950\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17628\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__17628\,
            I => \N__17625\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__17625\,
            I => \b2v_inst11.count_0_8\
        );

    \I__1947\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17618\
        );

    \I__1946\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17615\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__17618\,
            I => \b2v_inst11.count_1_8\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__17615\,
            I => \b2v_inst11.count_1_8\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__17610\,
            I => \N__17607\
        );

    \I__1942\ : InMux
    port map (
            O => \N__17607\,
            I => \N__17601\
        );

    \I__1941\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17601\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__17601\,
            I => \b2v_inst11.count_1_9\
        );

    \I__1939\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17595\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__17595\,
            I => \b2v_inst11.count_0_9\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__17592\,
            I => \N__17589\
        );

    \I__1936\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17583\
        );

    \I__1935\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17583\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__17583\,
            I => \b2v_inst11.count_1_10\
        );

    \I__1933\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17577\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__17577\,
            I => \b2v_inst11.count_0_10\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__17574\,
            I => \N__17571\
        );

    \I__1930\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17565\
        );

    \I__1929\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17565\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__17565\,
            I => \b2v_inst11.count_1_11\
        );

    \I__1927\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17559\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__17559\,
            I => \b2v_inst11.count_0_11\
        );

    \I__1925\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17553\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__17553\,
            I => \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJZ0Z62\
        );

    \I__1923\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17547\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__17547\,
            I => \b2v_inst11.curr_state_4_0\
        );

    \I__1921\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17541\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__17541\,
            I => \b2v_inst11.count_0_0\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__17538\,
            I => \b2v_inst11.countZ0Z_0_cascade_\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__17535\,
            I => \b2v_inst11.count_1_1_cascade_\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__17532\,
            I => \CONSTANT_ONE_NET_cascade_\
        );

    \I__1916\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17526\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__17526\,
            I => \N__17522\
        );

    \I__1914\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17519\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__17522\,
            I => \N__17516\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__17519\,
            I => \b2v_inst11.N_5852_i\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__17516\,
            I => \b2v_inst11.N_5852_i\
        );

    \I__1910\ : InMux
    port map (
            O => \N__17511\,
            I => \N__17505\
        );

    \I__1909\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17505\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__17505\,
            I => \b2v_inst16.un4_count_1_cry_8_THRU_CO\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__17502\,
            I => \b2v_inst16.countZ0Z_9_cascade_\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__17499\,
            I => \N__17495\
        );

    \I__1905\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17480\
        );

    \I__1904\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17480\
        );

    \I__1903\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17480\
        );

    \I__1902\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17464\
        );

    \I__1901\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17464\
        );

    \I__1900\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17464\
        );

    \I__1899\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17464\
        );

    \I__1898\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17464\
        );

    \I__1897\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17459\
        );

    \I__1896\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17459\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__17480\,
            I => \N__17456\
        );

    \I__1894\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17445\
        );

    \I__1893\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17445\
        );

    \I__1892\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17445\
        );

    \I__1891\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17445\
        );

    \I__1890\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17445\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__17464\,
            I => \N__17440\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__17459\,
            I => \N__17440\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__17456\,
            I => \b2v_inst16.N_416\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__17445\,
            I => \b2v_inst16.N_416\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__17440\,
            I => \b2v_inst16.N_416\
        );

    \I__1884\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__17430\,
            I => \b2v_inst16.count_4_9\
        );

    \I__1882\ : InMux
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__17424\,
            I => \b2v_inst16.count_4_10\
        );

    \I__1880\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17415\
        );

    \I__1879\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17415\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__17415\,
            I => \b2v_inst16.count_rst\
        );

    \I__1877\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17409\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__17409\,
            I => \N__17405\
        );

    \I__1875\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17402\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__17405\,
            I => \b2v_inst16.countZ0Z_10\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__17402\,
            I => \b2v_inst16.countZ0Z_10\
        );

    \I__1872\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17393\
        );

    \I__1871\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17390\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__17393\,
            I => \b2v_inst16.count_rst_1\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__17390\,
            I => \b2v_inst16.count_rst_1\
        );

    \I__1868\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17382\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__17382\,
            I => \b2v_inst16.count_4_12\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__17379\,
            I => \b2v_inst11.curr_state_3_0_cascade_\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__17376\,
            I => \b2v_inst11.curr_stateZ0Z_0_cascade_\
        );

    \I__1864\ : InMux
    port map (
            O => \N__17373\,
            I => \b2v_inst16.un4_count_1_cry_10\
        );

    \I__1863\ : InMux
    port map (
            O => \N__17370\,
            I => \b2v_inst16.un4_count_1_cry_11\
        );

    \I__1862\ : InMux
    port map (
            O => \N__17367\,
            I => \b2v_inst16.un4_count_1_cry_12\
        );

    \I__1861\ : InMux
    port map (
            O => \N__17364\,
            I => \b2v_inst16.un4_count_1_cry_13\
        );

    \I__1860\ : InMux
    port map (
            O => \N__17361\,
            I => \b2v_inst16.un4_count_1_cry_14\
        );

    \I__1859\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17354\
        );

    \I__1858\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17351\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__17354\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__17351\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__1855\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17342\
        );

    \I__1854\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17339\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__17342\,
            I => \N__17334\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__17339\,
            I => \N__17334\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__17334\,
            I => \b2v_inst16.un4_count_1_cry_7_THRU_CO\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__1849\ : InMux
    port map (
            O => \N__17328\,
            I => \N__17323\
        );

    \I__1848\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17320\
        );

    \I__1847\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17317\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__17323\,
            I => \N__17314\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__17320\,
            I => \N__17311\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__17317\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__17314\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__17311\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1841\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17301\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__17301\,
            I => \b2v_inst16.count_rst_13\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__17298\,
            I => \b2v_inst16.count_rst_14_cascade_\
        );

    \I__1838\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17291\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__17294\,
            I => \N__17288\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__17291\,
            I => \N__17284\
        );

    \I__1835\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17281\
        );

    \I__1834\ : InMux
    port map (
            O => \N__17287\,
            I => \N__17278\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__17284\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__17281\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__17278\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1830\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17264\
        );

    \I__1829\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17264\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__17269\,
            I => \N__17261\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17258\
        );

    \I__1826\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17255\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__17258\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__17255\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1823\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17246\
        );

    \I__1822\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17243\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__17246\,
            I => \b2v_inst16.un4_count_1_cry_2_THRU_CO\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__17243\,
            I => \b2v_inst16.un4_count_1_cry_2_THRU_CO\
        );

    \I__1819\ : InMux
    port map (
            O => \N__17238\,
            I => \b2v_inst16.un4_count_1_cry_2\
        );

    \I__1818\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17230\
        );

    \I__1817\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17227\
        );

    \I__1816\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17224\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__17230\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__17227\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__17224\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__17217\,
            I => \N__17213\
        );

    \I__1811\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17210\
        );

    \I__1810\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17207\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__17210\,
            I => \b2v_inst16.un4_count_1_cry_3_THRU_CO\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__17207\,
            I => \b2v_inst16.un4_count_1_cry_3_THRU_CO\
        );

    \I__1807\ : InMux
    port map (
            O => \N__17202\,
            I => \b2v_inst16.un4_count_1_cry_3\
        );

    \I__1806\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17196\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__17196\,
            I => \N__17192\
        );

    \I__1804\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17189\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__17192\,
            I => \N__17185\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17182\
        );

    \I__1801\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17179\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__17185\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__17182\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__17179\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__17172\,
            I => \N__17168\
        );

    \I__1796\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17165\
        );

    \I__1795\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17162\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17157\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__17162\,
            I => \N__17157\
        );

    \I__1792\ : Span4Mux_s1_h
    port map (
            O => \N__17157\,
            I => \N__17154\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__17154\,
            I => \b2v_inst16.un4_count_1_cry_4_THRU_CO\
        );

    \I__1790\ : InMux
    port map (
            O => \N__17151\,
            I => \b2v_inst16.un4_count_1_cry_4\
        );

    \I__1789\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17144\
        );

    \I__1788\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17141\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__17144\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__17141\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1785\ : InMux
    port map (
            O => \N__17136\,
            I => \b2v_inst16.un4_count_1_cry_5\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__17133\,
            I => \N__17129\
        );

    \I__1783\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17126\
        );

    \I__1782\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17123\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__17126\,
            I => \N__17119\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17116\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__17122\,
            I => \N__17113\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__17119\,
            I => \N__17110\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__17116\,
            I => \N__17107\
        );

    \I__1776\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17104\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__17110\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__17107\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__17104\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1772\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17091\
        );

    \I__1771\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17091\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__17091\,
            I => \N__17088\
        );

    \I__1769\ : Span4Mux_s1_h
    port map (
            O => \N__17088\,
            I => \N__17085\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__17085\,
            I => \b2v_inst16.un4_count_1_cry_6_THRU_CO\
        );

    \I__1767\ : InMux
    port map (
            O => \N__17082\,
            I => \b2v_inst16.un4_count_1_cry_6\
        );

    \I__1766\ : InMux
    port map (
            O => \N__17079\,
            I => \b2v_inst16.un4_count_1_cry_7\
        );

    \I__1765\ : InMux
    port map (
            O => \N__17076\,
            I => \bfn_2_7_0_\
        );

    \I__1764\ : InMux
    port map (
            O => \N__17073\,
            I => \b2v_inst16.un4_count_1_cry_9\
        );

    \I__1763\ : InMux
    port map (
            O => \N__17070\,
            I => \N__17066\
        );

    \I__1762\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17063\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__17066\,
            I => \N__17059\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__17063\,
            I => \N__17056\
        );

    \I__1759\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17053\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__17059\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__17056\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__17053\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1755\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17040\
        );

    \I__1754\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17040\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__17040\,
            I => \N__17037\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__17037\,
            I => \b2v_inst16.un4_count_1_cry_10_THRU_CO\
        );

    \I__1751\ : InMux
    port map (
            O => \N__17034\,
            I => \N__17031\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__17031\,
            I => \N__17027\
        );

    \I__1749\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17024\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__17027\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__17024\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__1746\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17016\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__17016\,
            I => \b2v_inst36.count_2_14\
        );

    \I__1744\ : CEMux
    port map (
            O => \N__17013\,
            I => \N__17008\
        );

    \I__1743\ : CEMux
    port map (
            O => \N__17012\,
            I => \N__17005\
        );

    \I__1742\ : CEMux
    port map (
            O => \N__17011\,
            I => \N__17002\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__17008\,
            I => \N__16994\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__17005\,
            I => \N__16994\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__17002\,
            I => \N__16994\
        );

    \I__1738\ : CEMux
    port map (
            O => \N__17001\,
            I => \N__16979\
        );

    \I__1737\ : Span4Mux_s2_v
    port map (
            O => \N__16994\,
            I => \N__16976\
        );

    \I__1736\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16973\
        );

    \I__1735\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16968\
        );

    \I__1734\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16968\
        );

    \I__1733\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16959\
        );

    \I__1732\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16959\
        );

    \I__1731\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16959\
        );

    \I__1730\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16959\
        );

    \I__1729\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16948\
        );

    \I__1728\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16948\
        );

    \I__1727\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16948\
        );

    \I__1726\ : InMux
    port map (
            O => \N__16983\,
            I => \N__16948\
        );

    \I__1725\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16948\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__16979\,
            I => \N__16939\
        );

    \I__1723\ : Span4Mux_s1_h
    port map (
            O => \N__16976\,
            I => \N__16924\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__16973\,
            I => \N__16924\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__16968\,
            I => \N__16924\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__16959\,
            I => \N__16924\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__16948\,
            I => \N__16924\
        );

    \I__1718\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16917\
        );

    \I__1717\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16917\
        );

    \I__1716\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16917\
        );

    \I__1715\ : CEMux
    port map (
            O => \N__16944\,
            I => \N__16911\
        );

    \I__1714\ : CEMux
    port map (
            O => \N__16943\,
            I => \N__16908\
        );

    \I__1713\ : CEMux
    port map (
            O => \N__16942\,
            I => \N__16905\
        );

    \I__1712\ : Span4Mux_s2_h
    port map (
            O => \N__16939\,
            I => \N__16902\
        );

    \I__1711\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16893\
        );

    \I__1710\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16893\
        );

    \I__1709\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16893\
        );

    \I__1708\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16893\
        );

    \I__1707\ : Sp12to4
    port map (
            O => \N__16924\,
            I => \N__16888\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16888\
        );

    \I__1705\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16881\
        );

    \I__1704\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16881\
        );

    \I__1703\ : InMux
    port map (
            O => \N__16914\,
            I => \N__16881\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__16911\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__16908\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__16905\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__16902\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__16893\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__16888\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__16881\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0\
        );

    \I__1695\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16860\
        );

    \I__1694\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16860\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__16860\,
            I => \N__16857\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__16857\,
            I => \b2v_inst36.count_rst\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__16854\,
            I => \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_\
        );

    \I__1690\ : InMux
    port map (
            O => \N__16851\,
            I => \N__16848\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__16848\,
            I => \b2v_inst36.count_2_15\
        );

    \I__1688\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16841\
        );

    \I__1687\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16838\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__16841\,
            I => \N__16833\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16833\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__16833\,
            I => \b2v_inst36.countZ0Z_15\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__16830\,
            I => \b2v_inst16.count_en_cascade_\
        );

    \I__1682\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16823\
        );

    \I__1681\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16820\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__16823\,
            I => \b2v_inst16.un4_count_1_axb_1\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__16820\,
            I => \b2v_inst16.un4_count_1_axb_1\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__16815\,
            I => \N__16812\
        );

    \I__1677\ : InMux
    port map (
            O => \N__16812\,
            I => \N__16806\
        );

    \I__1676\ : InMux
    port map (
            O => \N__16811\,
            I => \N__16801\
        );

    \I__1675\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16801\
        );

    \I__1674\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16798\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__16806\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__16801\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__16798\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1670\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16787\
        );

    \I__1669\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16784\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__16787\,
            I => \b2v_inst16.countZ0Z_2\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__16784\,
            I => \b2v_inst16.countZ0Z_2\
        );

    \I__1666\ : InMux
    port map (
            O => \N__16779\,
            I => \b2v_inst16.un4_count_1_cry_1\
        );

    \I__1665\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16773\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__16773\,
            I => \b2v_inst36.count_2_12\
        );

    \I__1663\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16764\
        );

    \I__1662\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16764\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__16764\,
            I => \b2v_inst36.count_rst_2\
        );

    \I__1660\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16758\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__16758\,
            I => \b2v_inst36.countZ0Z_12\
        );

    \I__1658\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16748\
        );

    \I__1657\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16748\
        );

    \I__1656\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16745\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__16748\,
            I => \b2v_inst36.count_rst_5\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__16745\,
            I => \b2v_inst36.count_rst_5\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__16740\,
            I => \b2v_inst36.countZ0Z_12_cascade_\
        );

    \I__1652\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16734\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__16734\,
            I => \N__16730\
        );

    \I__1650\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16727\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__16730\,
            I => \b2v_inst36.count_2_9\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__16727\,
            I => \b2v_inst36.count_2_9\
        );

    \I__1647\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16719\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__16719\,
            I => \b2v_inst36.un12_clk_100khz_6\
        );

    \I__1645\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16713\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__16713\,
            I => \b2v_inst36.countZ0Z_14\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__16710\,
            I => \b2v_inst36.countZ0Z_14_cascade_\
        );

    \I__1642\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16702\
        );

    \I__1641\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16697\
        );

    \I__1640\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16694\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__16702\,
            I => \N__16691\
        );

    \I__1638\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16686\
        );

    \I__1637\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16686\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__16697\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__16694\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__16691\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__16686\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__1632\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16674\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__16674\,
            I => \b2v_inst36.un12_clk_100khz_10\
        );

    \I__1630\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16668\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__16668\,
            I => \b2v_inst36.count_2_13\
        );

    \I__1628\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16659\
        );

    \I__1627\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16659\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__16659\,
            I => \b2v_inst36.count_rst_1\
        );

    \I__1625\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16652\
        );

    \I__1624\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16649\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__16652\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__16649\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__1621\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16641\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__16641\,
            I => \N__16637\
        );

    \I__1619\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16634\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__16637\,
            I => \b2v_inst36.un2_count_1_axb_8\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__16634\,
            I => \b2v_inst36.un2_count_1_axb_8\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__16629\,
            I => \N__16625\
        );

    \I__1615\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16620\
        );

    \I__1614\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16620\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__16620\,
            I => \b2v_inst36.un2_count_1_cry_7_THRU_CO\
        );

    \I__1612\ : InMux
    port map (
            O => \N__16617\,
            I => \b2v_inst36.un2_count_1_cry_7\
        );

    \I__1611\ : InMux
    port map (
            O => \N__16614\,
            I => \bfn_2_3_0_\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__16611\,
            I => \N__16607\
        );

    \I__1609\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16603\
        );

    \I__1608\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16600\
        );

    \I__1607\ : InMux
    port map (
            O => \N__16606\,
            I => \N__16597\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__16603\,
            I => \N__16592\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__16600\,
            I => \N__16592\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__16597\,
            I => \N__16589\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__16592\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__16589\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__1601\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16580\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16577\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__16580\,
            I => \N__16574\
        );

    \I__1598\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16571\
        );

    \I__1597\ : Span4Mux_s2_v
    port map (
            O => \N__16574\,
            I => \N__16566\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16566\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__16566\,
            I => \b2v_inst36.un2_count_1_cry_9_THRU_CO\
        );

    \I__1594\ : InMux
    port map (
            O => \N__16563\,
            I => \b2v_inst36.un2_count_1_cry_9\
        );

    \I__1593\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16556\
        );

    \I__1592\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16552\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__16556\,
            I => \N__16549\
        );

    \I__1590\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16546\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__16552\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__16549\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__16546\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__1586\ : InMux
    port map (
            O => \N__16539\,
            I => \N__16535\
        );

    \I__1585\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16532\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__16535\,
            I => \b2v_inst36.un2_count_1_cry_10_THRU_CO\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__16532\,
            I => \b2v_inst36.un2_count_1_cry_10_THRU_CO\
        );

    \I__1582\ : InMux
    port map (
            O => \N__16527\,
            I => \b2v_inst36.un2_count_1_cry_10\
        );

    \I__1581\ : InMux
    port map (
            O => \N__16524\,
            I => \b2v_inst36.un2_count_1_cry_11\
        );

    \I__1580\ : InMux
    port map (
            O => \N__16521\,
            I => \b2v_inst36.un2_count_1_cry_12\
        );

    \I__1579\ : InMux
    port map (
            O => \N__16518\,
            I => \b2v_inst36.un2_count_1_cry_13\
        );

    \I__1578\ : InMux
    port map (
            O => \N__16515\,
            I => \b2v_inst36.un2_count_1_cry_14\
        );

    \I__1577\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16509\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__16509\,
            I => \b2v_inst36.un2_count_1_axb_9\
        );

    \I__1575\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16503\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__16503\,
            I => \b2v_inst36.count_2_7\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__16500\,
            I => \N__16497\
        );

    \I__1572\ : InMux
    port map (
            O => \N__16497\,
            I => \N__16492\
        );

    \I__1571\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16487\
        );

    \I__1570\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16487\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__16492\,
            I => \N__16484\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__16487\,
            I => \b2v_inst36.un2_count_1_axb_1\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__16484\,
            I => \b2v_inst36.un2_count_1_axb_1\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__16479\,
            I => \N__16475\
        );

    \I__1565\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16469\
        );

    \I__1564\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16469\
        );

    \I__1563\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16466\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__16469\,
            I => \b2v_inst36.un2_count_1_axb_2\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__16466\,
            I => \b2v_inst36.un2_count_1_axb_2\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__16461\,
            I => \N__16458\
        );

    \I__1559\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16452\
        );

    \I__1558\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16452\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__16452\,
            I => \b2v_inst36.un2_count_1_cry_1_THRU_CO\
        );

    \I__1556\ : InMux
    port map (
            O => \N__16449\,
            I => \b2v_inst36.un2_count_1_cry_1\
        );

    \I__1555\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16439\
        );

    \I__1554\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16439\
        );

    \I__1553\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16436\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__16439\,
            I => \b2v_inst36.countZ0Z_3\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__16436\,
            I => \b2v_inst36.countZ0Z_3\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__16431\,
            I => \N__16427\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__16430\,
            I => \N__16424\
        );

    \I__1548\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16419\
        );

    \I__1547\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16419\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__16419\,
            I => \b2v_inst36.un2_count_1_cry_2_THRU_CO\
        );

    \I__1545\ : InMux
    port map (
            O => \N__16416\,
            I => \b2v_inst36.un2_count_1_cry_2\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__16413\,
            I => \N__16410\
        );

    \I__1543\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16407\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__16407\,
            I => \b2v_inst36.un2_count_1_axb_4\
        );

    \I__1541\ : InMux
    port map (
            O => \N__16404\,
            I => \N__16397\
        );

    \I__1540\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16397\
        );

    \I__1539\ : InMux
    port map (
            O => \N__16402\,
            I => \N__16394\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__16397\,
            I => \b2v_inst36.count_rst_10\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__16394\,
            I => \b2v_inst36.count_rst_10\
        );

    \I__1536\ : InMux
    port map (
            O => \N__16389\,
            I => \b2v_inst36.un2_count_1_cry_3\
        );

    \I__1535\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16382\
        );

    \I__1534\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16379\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__16382\,
            I => \b2v_inst36.un2_count_1_axb_5\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__16379\,
            I => \b2v_inst36.un2_count_1_axb_5\
        );

    \I__1531\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16368\
        );

    \I__1530\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16368\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__16368\,
            I => \b2v_inst36.un2_count_1_cry_4_THRU_CO\
        );

    \I__1528\ : InMux
    port map (
            O => \N__16365\,
            I => \b2v_inst36.un2_count_1_cry_4\
        );

    \I__1527\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16359\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__16359\,
            I => \b2v_inst36.un2_count_1_axb_6\
        );

    \I__1525\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16347\
        );

    \I__1524\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16347\
        );

    \I__1523\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16347\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__16347\,
            I => \b2v_inst36.un2_count_1_cry_5_c_RNIE2FZ0Z8\
        );

    \I__1521\ : InMux
    port map (
            O => \N__16344\,
            I => \b2v_inst36.un2_count_1_cry_5\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__16341\,
            I => \N__16338\
        );

    \I__1519\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16333\
        );

    \I__1518\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16329\
        );

    \I__1517\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16326\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__16333\,
            I => \N__16323\
        );

    \I__1515\ : InMux
    port map (
            O => \N__16332\,
            I => \N__16320\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__16329\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__16326\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__16323\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__16320\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__1510\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16307\
        );

    \I__1509\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16304\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__16307\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__16304\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__1506\ : InMux
    port map (
            O => \N__16299\,
            I => \b2v_inst36.un2_count_1_cry_6\
        );

    \I__1505\ : InMux
    port map (
            O => \N__16296\,
            I => \bfn_1_16_0_\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__16293\,
            I => \b2v_inst36.count_rst_12_cascade_\
        );

    \I__1503\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16287\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__16287\,
            I => \b2v_inst36.count_rst_12\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__16284\,
            I => \b2v_inst36.countZ0Z_3_cascade_\
        );

    \I__1500\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16278\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__16278\,
            I => \N__16275\
        );

    \I__1498\ : Span4Mux_s1_h
    port map (
            O => \N__16275\,
            I => \N__16272\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__16272\,
            I => \b2v_inst36.un12_clk_100khz_3\
        );

    \I__1496\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16266\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__16266\,
            I => \b2v_inst36.count_rst_11\
        );

    \I__1494\ : InMux
    port map (
            O => \N__16263\,
            I => \N__16257\
        );

    \I__1493\ : InMux
    port map (
            O => \N__16262\,
            I => \N__16257\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__16257\,
            I => \b2v_inst36.count_2_2\
        );

    \I__1491\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16251\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__16251\,
            I => \b2v_inst36.count_2_3\
        );

    \I__1489\ : InMux
    port map (
            O => \N__16248\,
            I => \N__16242\
        );

    \I__1488\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16242\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__16242\,
            I => \N__16239\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__16239\,
            I => \b2v_inst11.count_1_6\
        );

    \I__1485\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16233\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__16233\,
            I => \b2v_inst11.count_0_6\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__16230\,
            I => \N__16227\
        );

    \I__1482\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16221\
        );

    \I__1481\ : InMux
    port map (
            O => \N__16226\,
            I => \N__16221\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__16221\,
            I => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\
        );

    \I__1479\ : InMux
    port map (
            O => \N__16218\,
            I => \N__16215\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__16215\,
            I => \b2v_inst11.count_0_15\
        );

    \I__1477\ : InMux
    port map (
            O => \N__16212\,
            I => \b2v_inst11.un1_count_cry_11\
        );

    \I__1476\ : InMux
    port map (
            O => \N__16209\,
            I => \b2v_inst11.un1_count_cry_12\
        );

    \I__1475\ : InMux
    port map (
            O => \N__16206\,
            I => \b2v_inst11.un1_count_cry_13\
        );

    \I__1474\ : InMux
    port map (
            O => \N__16203\,
            I => \b2v_inst11.un1_count_cry_14\
        );

    \I__1473\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16194\
        );

    \I__1472\ : InMux
    port map (
            O => \N__16199\,
            I => \N__16194\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16191\
        );

    \I__1470\ : Odrv4
    port map (
            O => \N__16191\,
            I => \b2v_inst11.count_1_5\
        );

    \I__1469\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16185\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__16185\,
            I => \b2v_inst11.count_0_5\
        );

    \I__1467\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16178\
        );

    \I__1466\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16175\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__16178\,
            I => \b2v_inst11.count_1_14\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__16175\,
            I => \b2v_inst11.count_1_14\
        );

    \I__1463\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16167\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__16167\,
            I => \b2v_inst11.count_0_14\
        );

    \I__1461\ : InMux
    port map (
            O => \N__16164\,
            I => \b2v_inst11.un1_count_cry_2_cZ0\
        );

    \I__1460\ : InMux
    port map (
            O => \N__16161\,
            I => \b2v_inst11.un1_count_cry_3\
        );

    \I__1459\ : InMux
    port map (
            O => \N__16158\,
            I => \b2v_inst11.un1_count_cry_4\
        );

    \I__1458\ : InMux
    port map (
            O => \N__16155\,
            I => \b2v_inst11.un1_count_cry_5\
        );

    \I__1457\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16148\
        );

    \I__1456\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16145\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__16148\,
            I => \N__16142\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__16145\,
            I => \b2v_inst11.count_1_7\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__16142\,
            I => \b2v_inst11.count_1_7\
        );

    \I__1452\ : InMux
    port map (
            O => \N__16137\,
            I => \b2v_inst11.un1_count_cry_6\
        );

    \I__1451\ : InMux
    port map (
            O => \N__16134\,
            I => \b2v_inst11.un1_count_cry_7\
        );

    \I__1450\ : InMux
    port map (
            O => \N__16131\,
            I => \bfn_1_12_0_\
        );

    \I__1449\ : InMux
    port map (
            O => \N__16128\,
            I => \b2v_inst11.un1_count_cry_9\
        );

    \I__1448\ : InMux
    port map (
            O => \N__16125\,
            I => \b2v_inst11.un1_count_cry_10\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__16122\,
            I => \b2v_inst16.curr_state_7_0_1_cascade_\
        );

    \I__1446\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16116\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__16116\,
            I => \N__16113\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__16113\,
            I => \N__16110\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__16110\,
            I => \N__16107\
        );

    \I__1442\ : Sp12to4
    port map (
            O => \N__16107\,
            I => \N__16104\
        );

    \I__1441\ : Odrv12
    port map (
            O => \N__16104\,
            I => vddq_ok
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__16101\,
            I => \b2v_inst16.N_208_0_cascade_\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__16098\,
            I => \b2v_inst16.curr_state_RNIBO6I1Z0Z_0_cascade_\
        );

    \I__1438\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16092\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__16092\,
            I => \b2v_inst16.curr_state_2_1\
        );

    \I__1436\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16086\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__16086\,
            I => \b2v_inst16.curr_state_2_0\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__16083\,
            I => \N__16080\
        );

    \I__1433\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16077\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__16077\,
            I => \b2v_inst11.count_0_7\
        );

    \I__1431\ : InMux
    port map (
            O => \N__16074\,
            I => \b2v_inst11.un1_count_cry_1_cZ0\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__16071\,
            I => \b2v_inst16.countZ0Z_7_cascade_\
        );

    \I__1429\ : InMux
    port map (
            O => \N__16068\,
            I => \N__16065\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__16065\,
            I => \b2v_inst16.count_4_7\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__16062\,
            I => \b2v_inst16.count_rst_10_cascade_\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__16059\,
            I => \b2v_inst16.countZ0Z_5_cascade_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16053\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__16053\,
            I => \b2v_inst16.count_4_5\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__16050\,
            I => \b2v_inst16.countZ0Z_8_cascade_\
        );

    \I__1422\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16044\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__16044\,
            I => \b2v_inst16.count_4_8\
        );

    \I__1420\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16038\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__16038\,
            I => \b2v_inst16.count_rst_12\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__16035\,
            I => \b2v_inst16.N_416_cascade_\
        );

    \I__1417\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16029\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__16029\,
            I => \b2v_inst16.count_rst_8\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__16026\,
            I => \b2v_inst16.count_RNIE4RF_2Z0Z_1_cascade_\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__16023\,
            I => \b2v_inst16.count_rst_5_cascade_\
        );

    \I__1413\ : InMux
    port map (
            O => \N__16020\,
            I => \N__16014\
        );

    \I__1412\ : InMux
    port map (
            O => \N__16019\,
            I => \N__16014\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__16014\,
            I => \b2v_inst16.N_414\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__16011\,
            I => \b2v_inst16.countZ0Z_0_cascade_\
        );

    \I__1409\ : InMux
    port map (
            O => \N__16008\,
            I => \N__16005\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__16005\,
            I => \b2v_inst16.count_4_0\
        );

    \I__1407\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15999\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__15999\,
            I => \b2v_inst16.countZ0Z_1\
        );

    \I__1405\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15993\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__15993\,
            I => \b2v_inst16.count_4_i_a3_7_0\
        );

    \I__1403\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15984\
        );

    \I__1402\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15984\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__15984\,
            I => \b2v_inst16.count_RNIE4RF_2Z0Z_1\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__15981\,
            I => \N__15977\
        );

    \I__1399\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15972\
        );

    \I__1398\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15972\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__15972\,
            I => \b2v_inst16.count_4_1\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__15969\,
            I => \b2v_inst16.count_rst_9_cascade_\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__15966\,
            I => \b2v_inst16.countZ0Z_4_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15960\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__15960\,
            I => \b2v_inst16.count_4_4\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__15957\,
            I => \b2v_inst16.countZ0Z_3_cascade_\
        );

    \I__1391\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15951\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__15951\,
            I => \b2v_inst16.count_4_3\
        );

    \I__1389\ : InMux
    port map (
            O => \N__15948\,
            I => \N__15945\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__15945\,
            I => \b2v_inst16.count_4_i_a3_9_0\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__15942\,
            I => \b2v_inst16.count_4_i_a3_8_0_cascade_\
        );

    \I__1386\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15936\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__15936\,
            I => \b2v_inst16.count_4_i_a3_10_0\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__15933\,
            I => \b2v_inst16.N_414_cascade_\
        );

    \I__1383\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15927\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__15927\,
            I => \b2v_inst36.un12_clk_100khz_1\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__15924\,
            I => \b2v_inst36.un12_clk_100khz_0_cascade_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15918\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__15918\,
            I => \N__15915\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__15915\,
            I => \b2v_inst36.un12_clk_100khz_2\
        );

    \I__1377\ : InMux
    port map (
            O => \N__15912\,
            I => \N__15909\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__15909\,
            I => \N__15906\
        );

    \I__1375\ : Odrv12
    port map (
            O => \N__15906\,
            I => \b2v_inst36.un12_clk_100khz_7\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__15903\,
            I => \b2v_inst36.un12_clk_100khz_12_cascade_\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__15900\,
            I => \b2v_inst36.N_1_i_cascade_\
        );

    \I__1372\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15894\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__15894\,
            I => \b2v_inst36.count_2_0\
        );

    \I__1370\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15888\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__15888\,
            I => \b2v_inst36.count_rst_14\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__15885\,
            I => \b2v_inst36.countZ0Z_0_cascade_\
        );

    \I__1367\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15876\
        );

    \I__1366\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15876\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__15876\,
            I => \b2v_inst36.count_2_1\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__15873\,
            I => \b2v_inst16.count_rst_0_cascade_\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__15870\,
            I => \b2v_inst16.countZ0Z_11_cascade_\
        );

    \I__1362\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15864\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__15864\,
            I => \N__15861\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__15861\,
            I => \b2v_inst16.count_4_11\
        );

    \I__1359\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15855\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__15855\,
            I => \b2v_inst36.count_rst_6\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__15852\,
            I => \b2v_inst36.count_rst_6_cascade_\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \b2v_inst36.un2_count_1_axb_8_cascade_\
        );

    \I__1355\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15840\
        );

    \I__1354\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15840\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__15840\,
            I => \b2v_inst36.count_2_8\
        );

    \I__1352\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15834\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__15834\,
            I => \N__15831\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__15831\,
            I => \b2v_inst36.count_rst_4\
        );

    \I__1349\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15825\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__15825\,
            I => \b2v_inst36.count_rst_3\
        );

    \I__1347\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15819\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__15819\,
            I => \b2v_inst36.count_rst_13\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \b2v_inst36.count_rst_13_cascade_\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__15813\,
            I => \b2v_inst36.count_rst_7_cascade_\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__15810\,
            I => \b2v_inst36.countZ0Z_6_cascade_\
        );

    \I__1342\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15801\
        );

    \I__1341\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15801\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__15801\,
            I => \b2v_inst36.count_2_4\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__15798\,
            I => \b2v_inst36.countZ0Z_11_cascade_\
        );

    \I__1338\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15792\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__15792\,
            I => \b2v_inst36.count_2_11\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__15789\,
            I => \N__15785\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__15788\,
            I => \N__15782\
        );

    \I__1334\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15777\
        );

    \I__1333\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15777\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__15777\,
            I => \b2v_inst36.count_2_6\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__15774\,
            I => \b2v_inst36.countZ0Z_10_cascade_\
        );

    \I__1330\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15768\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__15768\,
            I => \b2v_inst36.count_2_10\
        );

    \I__1328\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15762\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__15762\,
            I => \b2v_inst36.count_rst_9\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__15759\,
            I => \b2v_inst36.count_rst_9_cascade_\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__15756\,
            I => \b2v_inst36.un2_count_1_axb_5_cascade_\
        );

    \I__1324\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15747\
        );

    \I__1323\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15747\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__15747\,
            I => \b2v_inst36.count_2_5\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst6.un2_count_1_cry_8\,
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst5.un2_count_1_cry_7\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst36.un2_count_1_cry_8\,
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_8\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_16\,
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => b2v_inst20_un4_counter_7,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_8\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_16\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_24\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst16.un4_count_1_cry_8\,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_0_cry_7\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz0\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un3_count_off_1_cry_8\,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_94_cry_7_s1\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_94_cry_7_s0\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_cry_8\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_1_cry_8\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_12_0_\
        );

    \b2v_inst200.count_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19860\,
            GLOBALBUFFEROUTPUT => \b2v_inst200.count_en_g\
        );

    \N_607_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35828\,
            GLOBALBUFFEROUTPUT => \N_607_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \b2v_inst36.count_RNIJKUH1_0_5_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__15765\,
            in1 => \N__15753\,
            in2 => \N__16341\,
            in3 => \N__16990\,
            lcout => \b2v_inst36.un12_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI4VQN1_10_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16989\,
            in1 => \N__15771\,
            in2 => \_gnd_net_\,
            in3 => \N__15837\,
            lcout => \b2v_inst36.countZ0Z_10\,
            ltout => \b2v_inst36.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_10_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19525\,
            in1 => \N__16584\,
            in2 => \N__15774\,
            in3 => \N__19070\,
            lcout => \b2v_inst36.count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36942\,
            ce => \N__17012\,
            sr => \N__19557\
        );

    \b2v_inst36.un2_count_1_cry_4_c_RNI8RQI_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__19068\,
            in1 => \N__16386\,
            in2 => \N__19543\,
            in3 => \N__16373\,
            lcout => \b2v_inst36.count_rst_9\,
            ltout => \b2v_inst36.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIJKUH1_5_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15752\,
            in2 => \N__15759\,
            in3 => \N__16987\,
            lcout => \b2v_inst36.un2_count_1_axb_5\,
            ltout => \b2v_inst36.un2_count_1_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_5_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19069\,
            in1 => \N__16374\,
            in2 => \N__15756\,
            in3 => \N__19526\,
            lcout => \b2v_inst36.count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36942\,
            ce => \N__17012\,
            sr => \N__19557\
        );

    \b2v_inst36.un2_count_1_cry_6_c_RNIAVSI_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__19524\,
            in1 => \N__16310\,
            in2 => \N__19083\,
            in3 => \N__16337\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNINQ0I1_7_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16988\,
            in1 => \_gnd_net_\,
            in2 => \N__15813\,
            in3 => \N__16506\,
            lcout => \b2v_inst36.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_6_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__16356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19509\,
            lcout => \b2v_inst36.count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36898\,
            ce => \N__17001\,
            sr => \N__19541\
        );

    \b2v_inst36.count_RNIHHTH1_4_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15806\,
            in1 => \N__16982\,
            in2 => \_gnd_net_\,
            in3 => \N__16402\,
            lcout => \b2v_inst36.un2_count_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_4_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16404\,
            lcout => \b2v_inst36.count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36898\,
            ce => \N__17001\,
            sr => \N__19541\
        );

    \b2v_inst36.count_RNILNVH1_6_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__19507\,
            in1 => \N__16985\,
            in2 => \N__15789\,
            in3 => \N__16355\,
            lcout => OPEN,
            ltout => \b2v_inst36.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI69T33_4_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__16986\,
            in1 => \N__16403\,
            in2 => \N__15810\,
            in3 => \N__15807\,
            lcout => \b2v_inst36.un12_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIDPQG1_11_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15795\,
            in1 => \N__16984\,
            in2 => \_gnd_net_\,
            in3 => \N__15828\,
            lcout => \b2v_inst36.countZ0Z_11\,
            ltout => \b2v_inst36.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_11_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__19080\,
            in1 => \N__19508\,
            in2 => \N__15798\,
            in3 => \N__16539\,
            lcout => \b2v_inst36.count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36898\,
            ce => \N__17001\,
            sr => \N__19541\
        );

    \b2v_inst36.count_RNILNVH1_0_6_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__19506\,
            in1 => \N__16983\,
            in2 => \N__15788\,
            in3 => \N__16354\,
            lcout => \b2v_inst36.un2_count_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIPT1I1_0_8_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__15858\,
            in1 => \N__15846\,
            in2 => \N__16611\,
            in3 => \N__16992\,
            lcout => \b2v_inst36.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_c_RNIB1UI_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19456\,
            in1 => \N__16644\,
            in2 => \N__16629\,
            in3 => \N__19020\,
            lcout => \b2v_inst36.count_rst_6\,
            ltout => \b2v_inst36.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIPT1I1_8_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15845\,
            in2 => \N__15852\,
            in3 => \N__16991\,
            lcout => \b2v_inst36.un2_count_1_axb_8\,
            ltout => \b2v_inst36.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_8_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16628\,
            in1 => \N__19445\,
            in2 => \N__15849\,
            in3 => \N__19025\,
            lcout => \b2v_inst36.count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36889\,
            ce => \N__17013\,
            sr => \N__19505\
        );

    \b2v_inst36.un2_count_1_cry_9_c_RNID50J_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19021\,
            in1 => \N__16610\,
            in2 => \N__16583\,
            in3 => \N__19457\,
            lcout => \b2v_inst36.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIRQCA_0_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16705\,
            in1 => \N__19444\,
            in2 => \_gnd_net_\,
            in3 => \N__19019\,
            lcout => \b2v_inst36.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_c_RNILUVB_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__16559\,
            in1 => \N__19458\,
            in2 => \N__19060\,
            in3 => \N__16538\,
            lcout => \b2v_inst36.count_rst_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI2GG91_1_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15881\,
            in1 => \N__16915\,
            in2 => \_gnd_net_\,
            in3 => \N__15822\,
            lcout => \b2v_inst36.un2_count_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIRQCA_1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__16495\,
            in1 => \N__16700\,
            in2 => \_gnd_net_\,
            in3 => \N__19467\,
            lcout => \b2v_inst36.count_rst_13\,
            ltout => \b2v_inst36.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI2GG91_0_1_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__15882\,
            in1 => \N__16916\,
            in2 => \N__15816\,
            in3 => \N__16560\,
            lcout => OPEN,
            ltout => \b2v_inst36.un12_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIRDCV5_1_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16281\,
            in1 => \N__15930\,
            in2 => \N__15924\,
            in3 => \N__15921\,
            lcout => OPEN,
            ltout => \b2v_inst36.un12_clk_100khz_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNISNCLA_4_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15912\,
            in1 => \N__16722\,
            in2 => \N__15903\,
            in3 => \N__16677\,
            lcout => \b2v_inst36.N_1_i\,
            ltout => \b2v_inst36.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_0_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16701\,
            in2 => \N__15900\,
            in3 => \N__19559\,
            lcout => \b2v_inst36.count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37101\,
            ce => \N__16944\,
            sr => \N__19558\
        );

    \b2v_inst36.count_RNI1FG91_0_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15897\,
            in1 => \N__16914\,
            in2 => \_gnd_net_\,
            in3 => \N__15891\,
            lcout => \b2v_inst36.countZ0Z_0\,
            ltout => \b2v_inst36.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__16496\,
            in1 => \_gnd_net_\,
            in2 => \N__15885\,
            in3 => \N__19560\,
            lcout => \b2v_inst36.count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37101\,
            ce => \N__16944\,
            sr => \N__19558\
        );

    \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__17062\,
            in1 => \N__17045\,
            in2 => \N__19806\,
            in3 => \N__17476\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIV7UA_11_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19222\,
            in1 => \_gnd_net_\,
            in2 => \N__15873\,
            in3 => \N__15867\,
            lcout => \b2v_inst16.countZ0Z_11\,
            ltout => \b2v_inst16.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_11_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__19803\,
            in1 => \N__17046\,
            in2 => \N__15870\,
            in3 => \N__17479\,
            lcout => \b2v_inst16.count_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37108\,
            ce => \N__19256\,
            sr => \N__19141\
        );

    \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17475\,
            in1 => \N__19802\,
            in2 => \N__17217\,
            in3 => \N__17233\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNITRJU_4_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15963\,
            in1 => \_gnd_net_\,
            in2 => \N__15969\,
            in3 => \N__19221\,
            lcout => \b2v_inst16.countZ0Z_4\,
            ltout => \b2v_inst16.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_4_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17478\,
            in1 => \N__19805\,
            in2 => \N__15966\,
            in3 => \N__17216\,
            lcout => \b2v_inst16.count_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37108\,
            ce => \N__19256\,
            sr => \N__19141\
        );

    \b2v_inst16.count_RNIROIU_3_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15954\,
            in1 => \N__16032\,
            in2 => \_gnd_net_\,
            in3 => \N__19223\,
            lcout => \b2v_inst16.countZ0Z_3\,
            ltout => \b2v_inst16.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_3_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17477\,
            in1 => \N__19804\,
            in2 => \N__15957\,
            in3 => \N__17249\,
            lcout => \b2v_inst16.count_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37108\,
            ce => \N__19256\,
            sr => \N__19141\
        );

    \b2v_inst16.count_RNI_10_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__17412\,
            in1 => \N__18915\,
            in2 => \N__18870\,
            in3 => \N__17327\,
            lcout => \b2v_inst16.count_4_i_a3_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_15_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17358\,
            in1 => \N__16791\,
            in2 => \N__18957\,
            in3 => \N__17148\,
            lcout => \b2v_inst16.count_4_i_a3_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17270\,
            in1 => \N__17195\,
            in2 => \N__17133\,
            in3 => \N__17234\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_4_i_a3_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIE4RF_3_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15996\,
            in1 => \N__15948\,
            in2 => \N__15942\,
            in3 => \N__15939\,
            lcout => \b2v_inst16.N_414\,
            ltout => \b2v_inst16.N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15933\,
            in3 => \N__16809\,
            lcout => \b2v_inst16.N_416\,
            ltout => \b2v_inst16.N_416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__19780\,
            in1 => \N__17271\,
            in2 => \N__16035\,
            in3 => \N__17250\,
            lcout => \b2v_inst16.count_rst_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIE4RF_2_1_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16810\,
            in2 => \_gnd_net_\,
            in3 => \N__16827\,
            lcout => \b2v_inst16.count_RNIE4RF_2Z0Z_1\,
            ltout => \b2v_inst16.count_RNIE4RF_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIE4RF_1_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19779\,
            in1 => \N__15980\,
            in2 => \N__16026\,
            in3 => \N__19275\,
            lcout => \b2v_inst16.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_0_0_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__16019\,
            in1 => \N__19775\,
            in2 => \_gnd_net_\,
            in3 => \N__16811\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNID3RF_0_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19241\,
            in1 => \_gnd_net_\,
            in2 => \N__16023\,
            in3 => \N__16008\,
            lcout => \b2v_inst16.countZ0Z_0\,
            ltout => \b2v_inst16.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_0_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__16020\,
            in1 => \_gnd_net_\,
            in2 => \N__16011\,
            in3 => \N__19778\,
            lcout => \b2v_inst16.count_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37109\,
            ce => \N__19274\,
            sr => \N__19130\
        );

    \b2v_inst16.count_RNIE4RF_1_1_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17295\,
            in1 => \N__16002\,
            in2 => \_gnd_net_\,
            in3 => \N__17069\,
            lcout => \b2v_inst16.count_4_i_a3_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIE4RF_0_1_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15989\,
            in1 => \N__19776\,
            in2 => \N__15981\,
            in3 => \N__19240\,
            lcout => \b2v_inst16.un4_count_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_1_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__19777\,
            in1 => \N__15990\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37109\,
            ce => \N__19274\,
            sr => \N__19130\
        );

    \b2v_inst16.count_RNI35NU_7_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19242\,
            in1 => \N__16068\,
            in2 => \_gnd_net_\,
            in3 => \N__16041\,
            lcout => \b2v_inst16.countZ0Z_7\,
            ltout => \b2v_inst16.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_7_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__19768\,
            in1 => \N__17493\,
            in2 => \N__16071\,
            in3 => \N__17097\,
            lcout => \b2v_inst16.count_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37139\,
            ce => \N__19273\,
            sr => \N__19137\
        );

    \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__17490\,
            in1 => \N__17188\,
            in2 => \N__17172\,
            in3 => \N__19767\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIVUKU_5_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16056\,
            in2 => \N__16062\,
            in3 => \N__19243\,
            lcout => \b2v_inst16.countZ0Z_5\,
            ltout => \b2v_inst16.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_5_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__17491\,
            in1 => \N__17171\,
            in2 => \N__16059\,
            in3 => \N__19770\,
            lcout => \b2v_inst16.count_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37139\,
            ce => \N__19273\,
            sr => \N__19137\
        );

    \b2v_inst16.count_RNI58OU_8_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16047\,
            in1 => \N__17304\,
            in2 => \_gnd_net_\,
            in3 => \N__19244\,
            lcout => \b2v_inst16.countZ0Z_8\,
            ltout => \b2v_inst16.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_8_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17492\,
            in1 => \N__19769\,
            in2 => \N__16050\,
            in3 => \N__17346\,
            lcout => \b2v_inst16.count_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37139\,
            ce => \N__19273\,
            sr => \N__19137\
        );

    \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__19766\,
            in1 => \N__17489\,
            in2 => \N__17122\,
            in3 => \N__17096\,
            lcout => \b2v_inst16.count_rst_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIBO6I1_1_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20477\,
            in1 => \N__19829\,
            in2 => \_gnd_net_\,
            in3 => \N__17487\,
            lcout => OPEN,
            ltout => \b2v_inst16.curr_state_7_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI4KJ02_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__28397\,
            in1 => \_gnd_net_\,
            in2 => \N__16122\,
            in3 => \N__16095\,
            lcout => \b2v_inst16.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__38529\,
            in1 => \N__16119\,
            in2 => \_gnd_net_\,
            in3 => \N__34833\,
            lcout => \b2v_inst16.N_208_0\,
            ltout => \b2v_inst16.N_208_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIBO6I1_0_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111111"
        )
    port map (
            in0 => \N__28395\,
            in1 => \_gnd_net_\,
            in2 => \N__16101\,
            in3 => \N__16089\,
            lcout => \b2v_inst16.curr_state_RNIBO6I1Z0Z_0\,
            ltout => \b2v_inst16.curr_state_RNIBO6I1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_1_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20475\,
            in2 => \N__16098\,
            in3 => \N__17488\,
            lcout => \b2v_inst16.curr_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37125\,
            ce => \N__27542\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIU6GN_7_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__28396\,
            in1 => \_gnd_net_\,
            in2 => \N__16083\,
            in3 => \N__16152\,
            lcout => \b2v_inst11.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_0_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__20476\,
            in1 => \N__20519\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37125\,
            ce => \N__27542\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_8_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17622\,
            lcout => \b2v_inst11.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37141\,
            ce => \N__27540\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_7_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16151\,
            lcout => \b2v_inst11.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37141\,
            ce => \N__27540\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20084\,
            in2 => \N__17663\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \b2v_inst11.un1_count_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20058\,
            in1 => \N__18262\,
            in2 => \_gnd_net_\,
            in3 => \N__16074\,
            lcout => \b2v_inst11.count_1_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_1_cZ0\,
            carryout => \b2v_inst11.un1_count_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20050\,
            in1 => \_gnd_net_\,
            in2 => \N__18245\,
            in3 => \N__16164\,
            lcout => \b2v_inst11.count_1_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_2_cZ0\,
            carryout => \b2v_inst11.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20059\,
            in1 => \_gnd_net_\,
            in2 => \N__18221\,
            in3 => \N__16161\,
            lcout => \b2v_inst11.count_1_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_3\,
            carryout => \b2v_inst11.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20051\,
            in1 => \_gnd_net_\,
            in2 => \N__18138\,
            in3 => \N__16158\,
            lcout => \b2v_inst11.count_1_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_4\,
            carryout => \b2v_inst11.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20060\,
            in1 => \_gnd_net_\,
            in2 => \N__18165\,
            in3 => \N__16155\,
            lcout => \b2v_inst11.count_1_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_5\,
            carryout => \b2v_inst11.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20052\,
            in1 => \_gnd_net_\,
            in2 => \N__18196\,
            in3 => \N__16137\,
            lcout => \b2v_inst11.count_1_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_6\,
            carryout => \b2v_inst11.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20061\,
            in1 => \_gnd_net_\,
            in2 => \N__17941\,
            in3 => \N__16134\,
            lcout => \b2v_inst11.count_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_7\,
            carryout => \b2v_inst11.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20053\,
            in1 => \_gnd_net_\,
            in2 => \N__17911\,
            in3 => \N__16131\,
            lcout => \b2v_inst11.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \b2v_inst11.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20062\,
            in1 => \_gnd_net_\,
            in2 => \N__18106\,
            in3 => \N__16128\,
            lcout => \b2v_inst11.count_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_9\,
            carryout => \b2v_inst11.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20054\,
            in1 => \_gnd_net_\,
            in2 => \N__18046\,
            in3 => \N__16125\,
            lcout => \b2v_inst11.count_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_10\,
            carryout => \b2v_inst11.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20063\,
            in1 => \_gnd_net_\,
            in2 => \N__18077\,
            in3 => \N__16212\,
            lcout => \b2v_inst11.count_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_11\,
            carryout => \b2v_inst11.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20055\,
            in1 => \_gnd_net_\,
            in2 => \N__18022\,
            in3 => \N__16209\,
            lcout => \b2v_inst11.count_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_12\,
            carryout => \b2v_inst11.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20064\,
            in1 => \_gnd_net_\,
            in2 => \N__17999\,
            in3 => \N__16206\,
            lcout => \b2v_inst11.count_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_13\,
            carryout => \b2v_inst11.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20056\,
            in1 => \N__17972\,
            in2 => \_gnd_net_\,
            in3 => \N__16203\,
            lcout => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQF4M_14_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16170\,
            in1 => \N__28409\,
            in2 => \_gnd_net_\,
            in3 => \N__16181\,
            lcout => \b2v_inst11.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQ0EN_5_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28406\,
            in1 => \N__16188\,
            in2 => \_gnd_net_\,
            in3 => \N__16199\,
            lcout => \b2v_inst11.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_5_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37148\,
            ce => \N__27533\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_14_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16182\,
            lcout => \b2v_inst11.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37148\,
            ce => \N__27533\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIS3FN_6_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28407\,
            in1 => \N__16236\,
            in2 => \_gnd_net_\,
            in3 => \N__16247\,
            lcout => \b2v_inst11.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_6_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16248\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37148\,
            ce => \N__27533\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNISI5M_15_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28408\,
            in1 => \N__16218\,
            in2 => \_gnd_net_\,
            in3 => \N__16226\,
            lcout => \b2v_inst11.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_15_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16230\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37148\,
            ce => \N__27533\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_0_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17529\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_1_c_inv_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17816\,
            in2 => \N__17804\,
            in3 => \N__17667\,
            lcout => \b2v_inst11.N_5853_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_0\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_2_c_inv_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17786\,
            in2 => \N__17775\,
            in3 => \N__18269\,
            lcout => \b2v_inst11.N_5854_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_1\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_3_c_inv_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18485\,
            in2 => \N__18473\,
            in3 => \N__18246\,
            lcout => \b2v_inst11.N_5855_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_2\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_4_c_inv_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18437\,
            in2 => \N__18456\,
            in3 => \N__18222\,
            lcout => \b2v_inst11.N_5856_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_3\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_5_c_inv_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18130\,
            in1 => \N__18425\,
            in2 => \N__18414\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5857_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_4\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_6_c_inv_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18392\,
            in2 => \N__18380\,
            in3 => \N__18160\,
            lcout => \b2v_inst11.N_5858_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_5\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_7_c_inv_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18359\,
            in2 => \N__18348\,
            in3 => \N__18197\,
            lcout => \b2v_inst11.N_5859_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_6\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_8_c_inv_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18332\,
            in2 => \N__18320\,
            in3 => \N__17946\,
            lcout => \b2v_inst11.N_5860_i\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_9_c_inv_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18302\,
            in2 => \N__18291\,
            in3 => \N__17916\,
            lcout => \b2v_inst11.N_5861_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_8\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_10_c_inv_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18680\,
            in2 => \N__18669\,
            in3 => \N__18111\,
            lcout => \b2v_inst11.N_5862_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_9\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_11_c_inv_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18644\,
            in2 => \N__18633\,
            in3 => \N__18053\,
            lcout => \b2v_inst11.N_5863_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_10\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_12_c_inv_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18611\,
            in2 => \N__18600\,
            in3 => \N__18081\,
            lcout => \b2v_inst11.N_5864_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_11\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_13_c_inv_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18567\,
            in2 => \N__18584\,
            in3 => \N__18023\,
            lcout => \b2v_inst11.N_5865_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_12\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_14_c_inv_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18533\,
            in2 => \N__18552\,
            in3 => \N__18000\,
            lcout => \b2v_inst11.N_5866_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_13\,
            carryout => \b2v_inst11.un85_clk_100khz_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_15_c_inv_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18503\,
            in2 => \N__18521\,
            in3 => \N__17973\,
            lcout => \b2v_inst11.N_5867_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_0_cry_14\,
            carryout => \b2v_inst11.un85_clk_100khz0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz0_THRU_LUT4_0_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16296\,
            lcout => \b2v_inst11.un85_clk_100khz0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_c_RNI5LNI_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19468\,
            in1 => \N__16457\,
            in2 => \N__16479\,
            in3 => \N__19061\,
            lcout => \b2v_inst36.count_rst_12\,
            ltout => \b2v_inst36.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIDBRH1_2_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16262\,
            in2 => \N__16293\,
            in3 => \N__16945\,
            lcout => \b2v_inst36.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIFESH1_3_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16946\,
            in1 => \N__16254\,
            in2 => \_gnd_net_\,
            in3 => \N__16269\,
            lcout => \b2v_inst36.countZ0Z_3\,
            ltout => \b2v_inst36.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIDBRH1_0_2_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__16290\,
            in1 => \N__16263\,
            in2 => \N__16284\,
            in3 => \N__16947\,
            lcout => \b2v_inst36.un12_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_c_RNI6NOI_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__19469\,
            in1 => \N__19062\,
            in2 => \N__16430\,
            in3 => \N__16446\,
            lcout => \b2v_inst36.count_rst_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_2_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19063\,
            in1 => \N__16478\,
            in2 => \N__16461\,
            in3 => \N__19549\,
            lcout => \b2v_inst36.count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36801\,
            ce => \N__17011\,
            sr => \N__19547\
        );

    \b2v_inst36.count_3_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__19470\,
            in1 => \N__19064\,
            in2 => \N__16431\,
            in3 => \N__16445\,
            lcout => \b2v_inst36.count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36801\,
            ce => \N__17011\,
            sr => \N__19547\
        );

    \b2v_inst36.count_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__16311\,
            in1 => \N__16336\,
            in2 => \N__19081\,
            in3 => \N__19548\,
            lcout => \b2v_inst36.count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36801\,
            ce => \N__17011\,
            sr => \N__19547\
        );

    \b2v_inst36.un2_count_1_cry_1_c_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16707\,
            in2 => \N__16500\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16474\,
            in2 => \_gnd_net_\,
            in3 => \N__16449\,
            lcout => \b2v_inst36.un2_count_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_1\,
            carryout => \b2v_inst36.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16444\,
            in2 => \_gnd_net_\,
            in3 => \N__16416\,
            lcout => \b2v_inst36.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_2\,
            carryout => \b2v_inst36.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_3_c_RNI7PPI_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19471\,
            in1 => \_gnd_net_\,
            in2 => \N__16413\,
            in3 => \N__16389\,
            lcout => \b2v_inst36.count_rst_10\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_3\,
            carryout => \b2v_inst36.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16385\,
            in2 => \_gnd_net_\,
            in3 => \N__16365\,
            lcout => \b2v_inst36.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_4\,
            carryout => \b2v_inst36.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16362\,
            in2 => \_gnd_net_\,
            in3 => \N__16344\,
            lcout => \b2v_inst36.un2_count_1_cry_5_c_RNIE2FZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_5\,
            carryout => \b2v_inst36.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16332\,
            in2 => \_gnd_net_\,
            in3 => \N__16299\,
            lcout => \b2v_inst36.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_6\,
            carryout => \b2v_inst36.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16640\,
            in2 => \_gnd_net_\,
            in3 => \N__16617\,
            lcout => \b2v_inst36.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_7\,
            carryout => \b2v_inst36.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_8_c_RNIC3VI_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19459\,
            in1 => \N__16512\,
            in2 => \_gnd_net_\,
            in3 => \N__16614\,
            lcout => \b2v_inst36.count_rst_5\,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16606\,
            in2 => \_gnd_net_\,
            in3 => \N__16563\,
            lcout => \b2v_inst36.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_9\,
            carryout => \b2v_inst36.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16555\,
            in2 => \_gnd_net_\,
            in3 => \N__16527\,
            lcout => \b2v_inst36.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_10\,
            carryout => \b2v_inst36.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_11_c_RNIM01C_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19462\,
            in1 => \N__16761\,
            in2 => \_gnd_net_\,
            in3 => \N__16524\,
            lcout => \b2v_inst36.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_11\,
            carryout => \b2v_inst36.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_12_c_RNIN22C_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19460\,
            in1 => \N__16655\,
            in2 => \_gnd_net_\,
            in3 => \N__16521\,
            lcout => \b2v_inst36.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_12\,
            carryout => \b2v_inst36.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_13_c_RNIO43C_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19463\,
            in1 => \N__16716\,
            in2 => \_gnd_net_\,
            in3 => \N__16518\,
            lcout => \b2v_inst36.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_13\,
            carryout => \b2v_inst36.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_14_c_RNIP64C_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19461\,
            in1 => \N__16845\,
            in2 => \_gnd_net_\,
            in3 => \N__16515\,
            lcout => \b2v_inst36.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIR03I1_9_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16733\,
            in1 => \N__16993\,
            in2 => \_gnd_net_\,
            in3 => \N__16753\,
            lcout => \b2v_inst36.un2_count_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_12_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16770\,
            lcout => \b2v_inst36.count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37027\,
            ce => \N__16943\,
            sr => \N__19530\
        );

    \b2v_inst36.count_9_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16755\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37027\,
            ce => \N__16943\,
            sr => \N__19530\
        );

    \b2v_inst36.count_RNIFSRG1_12_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16776\,
            in1 => \N__16935\,
            in2 => \_gnd_net_\,
            in3 => \N__16769\,
            lcout => \b2v_inst36.countZ0Z_12\,
            ltout => \b2v_inst36.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIR03I1_0_9_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__16938\,
            in1 => \N__16754\,
            in2 => \N__16740\,
            in3 => \N__16737\,
            lcout => \b2v_inst36.un12_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_13_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16665\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37027\,
            ce => \N__16943\,
            sr => \N__19530\
        );

    \b2v_inst36.count_RNIJ2UG1_14_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16937\,
            in1 => \N__17019\,
            in2 => \_gnd_net_\,
            in3 => \N__17030\,
            lcout => \b2v_inst36.countZ0Z_14\,
            ltout => \b2v_inst36.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_15_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16656\,
            in1 => \N__16844\,
            in2 => \N__16710\,
            in3 => \N__16706\,
            lcout => \b2v_inst36.un12_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIHVSG1_13_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16936\,
            in1 => \N__16671\,
            in2 => \_gnd_net_\,
            in3 => \N__16664\,
            lcout => \b2v_inst36.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_15_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16865\,
            lcout => \b2v_inst36.count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36966\,
            ce => \N__16942\,
            sr => \N__19542\
        );

    \b2v_inst36.count_14_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17034\,
            lcout => \b2v_inst36.count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36966\,
            ce => \N__16942\,
            sr => \N__19542\
        );

    \b2v_inst36.curr_state_RNINSDS_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__23090\,
            in1 => \N__23036\,
            in2 => \N__23148\,
            in3 => \N__27562\,
            lcout => \b2v_inst36.curr_state_RNINSDSZ0Z_0\,
            ltout => \b2v_inst36.curr_state_RNINSDSZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIL5VG1_15_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16866\,
            in1 => \_gnd_net_\,
            in2 => \N__16854\,
            in3 => \N__16851\,
            lcout => \b2v_inst36.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIPLHU_2_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19314\,
            in1 => \N__19325\,
            in2 => \_gnd_net_\,
            in3 => \N__19224\,
            lcout => \b2v_inst16.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIKEBL_1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__27563\,
            in1 => \N__19798\,
            in2 => \_gnd_net_\,
            in3 => \N__20486\,
            lcout => \b2v_inst16.count_en\,
            ltout => \b2v_inst16.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI12MU_6_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19287\,
            in2 => \N__16830\,
            in3 => \N__19305\,
            lcout => \b2v_inst16.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16826\,
            in2 => \N__16815\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__19781\,
            in1 => \N__16790\,
            in2 => \_gnd_net_\,
            in3 => \N__16779\,
            lcout => \b2v_inst16.count_rst_7\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_1\,
            carryout => \b2v_inst16.un4_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17269\,
            in3 => \N__17238\,
            lcout => \b2v_inst16.un4_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_2\,
            carryout => \b2v_inst16.un4_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17235\,
            in2 => \_gnd_net_\,
            in3 => \N__17202\,
            lcout => \b2v_inst16.un4_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_3\,
            carryout => \b2v_inst16.un4_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17199\,
            in2 => \_gnd_net_\,
            in3 => \N__17151\,
            lcout => \b2v_inst16.un4_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_4\,
            carryout => \b2v_inst16.un4_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__19782\,
            in1 => \N__17147\,
            in2 => \_gnd_net_\,
            in3 => \N__17136\,
            lcout => \b2v_inst16.count_rst_11\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_5\,
            carryout => \b2v_inst16.un4_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17132\,
            in2 => \_gnd_net_\,
            in3 => \N__17082\,
            lcout => \b2v_inst16.un4_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_6\,
            carryout => \b2v_inst16.un4_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17331\,
            in3 => \N__17079\,
            lcout => \b2v_inst16.un4_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_7\,
            carryout => \b2v_inst16.un4_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17287\,
            in2 => \_gnd_net_\,
            in3 => \N__17076\,
            lcout => \b2v_inst16.un4_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__19773\,
            in1 => \N__17408\,
            in2 => \_gnd_net_\,
            in3 => \N__17073\,
            lcout => \b2v_inst16.count_rst\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_9\,
            carryout => \b2v_inst16.un4_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17070\,
            in2 => \_gnd_net_\,
            in3 => \N__17373\,
            lcout => \b2v_inst16.un4_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_10\,
            carryout => \b2v_inst16.un4_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__19774\,
            in1 => \N__17357\,
            in2 => \_gnd_net_\,
            in3 => \N__17370\,
            lcout => \b2v_inst16.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_11\,
            carryout => \b2v_inst16.un4_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__19797\,
            in1 => \N__18911\,
            in2 => \_gnd_net_\,
            in3 => \N__17367\,
            lcout => \b2v_inst16.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_12\,
            carryout => \b2v_inst16.un4_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__19772\,
            in1 => \N__18866\,
            in2 => \_gnd_net_\,
            in3 => \N__17364\,
            lcout => \b2v_inst16.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_13\,
            carryout => \b2v_inst16.un4_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__18956\,
            in1 => \N__19771\,
            in2 => \_gnd_net_\,
            in3 => \N__17361\,
            lcout => \b2v_inst16.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIR4KE_12_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17385\,
            in1 => \N__17397\,
            in2 => \_gnd_net_\,
            in3 => \N__19245\,
            lcout => \b2v_inst16.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__19763\,
            in1 => \N__17345\,
            in2 => \N__17499\,
            in3 => \N__17326\,
            lcout => \b2v_inst16.count_rst_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__17511\,
            in1 => \N__19762\,
            in2 => \N__17294\,
            in3 => \N__17498\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI7BPU_9_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17433\,
            in2 => \N__17298\,
            in3 => \N__19247\,
            lcout => \b2v_inst16.countZ0Z_9\,
            ltout => \b2v_inst16.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_9_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__17510\,
            in1 => \N__19765\,
            in2 => \N__17502\,
            in3 => \N__17494\,
            lcout => \b2v_inst16.count_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37095\,
            ce => \N__19276\,
            sr => \N__19123\
        );

    \b2v_inst16.curr_state_RNI_0_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.N_3037_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_10_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17420\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37095\,
            ce => \N__19276\,
            sr => \N__19123\
        );

    \b2v_inst16.count_RNIG7TP_10_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17427\,
            in1 => \N__17421\,
            in2 => \_gnd_net_\,
            in3 => \N__19246\,
            lcout => \b2v_inst16.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_12_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17396\,
            lcout => \b2v_inst16.count_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37095\,
            ce => \N__19276\,
            sr => \N__19123\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_0_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__17859\,
            in1 => \N__17885\,
            in2 => \_gnd_net_\,
            in3 => \N__17556\,
            lcout => OPEN,
            ltout => \b2v_inst11.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNI82MVJ62_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17550\,
            in2 => \N__17379\,
            in3 => \N__28390\,
            lcout => \b2v_inst11.curr_stateZ0Z_0\,
            ltout => \b2v_inst11.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__28391\,
            in1 => \_gnd_net_\,
            in2 => \N__17376\,
            in3 => \N__17884\,
            lcout => \b2v_inst11.count_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNO_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17855\,
            in2 => \N__17886\,
            in3 => \N__28392\,
            lcout => \b2v_inst11.g0_0_0_rep1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJ62_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19595\,
            in1 => \N__19624\,
            in2 => \_gnd_net_\,
            in3 => \N__19949\,
            lcout => \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNILDIRJZ0Z62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__17860\,
            in1 => \N__17826\,
            in2 => \N__19626\,
            in3 => \N__19594\,
            lcout => \b2v_inst11.curr_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37062\,
            ce => \N__27541\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_0_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__28393\,
            in1 => \_gnd_net_\,
            in2 => \N__17864\,
            in3 => \N__17880\,
            lcout => \b2v_inst11.g0_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIKEBL_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27567\,
            in2 => \_gnd_net_\,
            in3 => \N__17854\,
            lcout => \b2v_inst11.g0_i_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__20086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20013\,
            lcout => \b2v_inst11.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37140\,
            ce => \N__27538\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI03G9_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17544\,
            in1 => \N__28351\,
            in2 => \_gnd_net_\,
            in3 => \N__19980\,
            lcout => \b2v_inst11.countZ0Z_0\,
            ltout => \b2v_inst11.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_1_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17662\,
            in2 => \N__17538\,
            in3 => \N__20012\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI14G9_1_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__28394\,
            in1 => \N__17637\,
            in2 => \N__17535\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => \CONSTANT_ONE_NET_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_0_cry_0_c_inv_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__17525\,
            in1 => \_gnd_net_\,
            in2 => \N__17532\,
            in3 => \N__20085\,
            lcout => \b2v_inst11.N_5852_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__20087\,
            in1 => \N__17661\,
            in2 => \_gnd_net_\,
            in3 => \N__20014\,
            lcout => \b2v_inst11.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37140\,
            ce => \N__27538\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI0AHN_8_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17631\,
            in1 => \N__28352\,
            in2 => \_gnd_net_\,
            in3 => \N__17621\,
            lcout => \b2v_inst11.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI2DIN_9_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17598\,
            in1 => \N__28399\,
            in2 => \_gnd_net_\,
            in3 => \N__17606\,
            lcout => \b2v_inst11.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_9_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17610\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37135\,
            ce => \N__27535\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIB49T_10_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17580\,
            in1 => \N__28400\,
            in2 => \_gnd_net_\,
            in3 => \N__17588\,
            lcout => \b2v_inst11.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_10_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17592\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37135\,
            ce => \N__27535\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIK61M_11_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17562\,
            in1 => \N__28401\,
            in2 => \_gnd_net_\,
            in3 => \N__17570\,
            lcout => \b2v_inst11.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_11_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17574\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37135\,
            ce => \N__27535\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIKNAN_2_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17742\,
            in2 => \N__17754\,
            in3 => \N__28398\,
            lcout => \b2v_inst11.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_2_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17753\,
            lcout => \b2v_inst11.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37135\,
            ce => \N__27535\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIM92M_12_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28404\,
            in1 => \N__17724\,
            in2 => \_gnd_net_\,
            in3 => \N__17732\,
            lcout => \b2v_inst11.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_12_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17736\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37134\,
            ce => \N__27534\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIMQBN_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28402\,
            in2 => \N__17709\,
            in3 => \N__17717\,
            lcout => \b2v_inst11.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37134\,
            ce => \N__27534\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOC3M_13_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28405\,
            in1 => \N__17688\,
            in2 => \_gnd_net_\,
            in3 => \N__17696\,
            lcout => \b2v_inst11.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_13_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17700\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37134\,
            ce => \N__27534\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOTCN_4_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28403\,
            in1 => \N__17673\,
            in2 => \_gnd_net_\,
            in3 => \N__17681\,
            lcout => \b2v_inst11.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_4_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37134\,
            ce => \N__27534\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_2_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18270\,
            in1 => \N__18244\,
            in2 => \_gnd_net_\,
            in3 => \N__18220\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_5_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__18198\,
            in1 => \N__18161\,
            in2 => \N__18141\,
            in3 => \N__18137\,
            lcout => \b2v_inst11.un79_clk_100khzlto15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_10_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18110\,
            in1 => \N__18076\,
            in2 => \N__18054\,
            in3 => \N__18024\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_15_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17998\,
            in2 => \N__17976\,
            in3 => \N__17971\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_8_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17952\,
            in1 => \N__17945\,
            in2 => \N__17919\,
            in3 => \N__17915\,
            lcout => \b2v_inst11.count_RNIZ0Z_8\,
            ltout => \b2v_inst11.count_RNIZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNO_0_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17865\,
            in2 => \N__17829\,
            in3 => \N__19950\,
            lcout => \b2v_inst11.curr_state_3_i_m2_0_rep1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_1_c_inv_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17817\,
            in2 => \N__17805\,
            in3 => \N__23886\,
            lcout => \b2v_inst11.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_2_c_inv_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17787\,
            in2 => \N__17774\,
            in3 => \N__24027\,
            lcout => \b2v_inst11.un85_clk_100khz_0_0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_1\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_3_c_inv_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18486\,
            in2 => \N__18474\,
            in3 => \N__23766\,
            lcout => \b2v_inst11.un85_clk_100khz_0_1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_2\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_4_c_inv_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18455\,
            in2 => \N__18441\,
            in3 => \N__20196\,
            lcout => \b2v_inst11.un85_clk_100khz_0_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_3\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_5_c_inv_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18426\,
            in2 => \N__18413\,
            in3 => \N__20616\,
            lcout => \b2v_inst11.un85_clk_100khz_0_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_4\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_6_c_inv_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18393\,
            in2 => \N__18381\,
            in3 => \N__20580\,
            lcout => \b2v_inst11.un85_clk_100khz_0_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_5\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_7_c_inv_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18347\,
            in2 => \N__18363\,
            in3 => \N__20424\,
            lcout => \b2v_inst11.un85_clk_100khz_0_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_6\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_8_c_inv_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18333\,
            in2 => \N__18321\,
            in3 => \N__21762\,
            lcout => \b2v_inst11.un85_clk_100khz_0_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_7\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_9_c_inv_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18303\,
            in2 => \N__18290\,
            in3 => \N__21868\,
            lcout => \b2v_inst11.un85_clk_100khz_0_7\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_10_c_inv_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18681\,
            in2 => \N__18668\,
            in3 => \N__22101\,
            lcout => \b2v_inst11.un85_clk_100khz_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_9\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_11_c_inv_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22068\,
            in1 => \N__18629\,
            in2 => \N__18648\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_1_9\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_10\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_12_c_inv_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18599\,
            in2 => \N__18615\,
            in3 => \N__24102\,
            lcout => \b2v_inst11.un85_clk_100khz_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_11\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_13_c_inv_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18566\,
            in2 => \N__18585\,
            in3 => \N__24198\,
            lcout => \b2v_inst11.un85_clk_100khz_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_12\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_14_c_inv_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18551\,
            in2 => \N__18537\,
            in3 => \N__25362\,
            lcout => \b2v_inst11.un85_clk_100khz_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_13\,
            carryout => \b2v_inst11.un85_clk_100khz_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_15_c_inv_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \N__18522\,
            in3 => \N__25326\,
            lcout => \b2v_inst11.un85_clk_100khz_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_1_cry_14\,
            carryout => \b2v_inst11.un85_clk_100khz1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz1_THRU_LUT4_0_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18492\,
            lcout => \b2v_inst11.un85_clk_100khz1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27069\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23964\,
            in2 => \N__18698\,
            in3 => \N__18489\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18694\,
            in2 => \N__21972\,
            in3 => \N__18714\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22093\,
            in2 => \N__21945\,
            in3 => \N__18711\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21921\,
            in2 => \N__22100\,
            in3 => \N__18708\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21867\,
            in1 => \N__22146\,
            in2 => \N__18699\,
            in3 => \N__18705\,
            lcout => \b2v_inst11.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22128\,
            in3 => \N__18702\,
            lcout => \b2v_inst11.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22092\,
            lcout => \b2v_inst11.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9S71_16_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18743\,
            in1 => \N__20974\,
            in2 => \_gnd_net_\,
            in3 => \N__22612\,
            lcout => \b2v_inst200.un2_count_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_16_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36800\,
            ce => \N__22541\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNID13N_0_1_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000111"
        )
    port map (
            in0 => \N__18756\,
            in1 => \N__22614\,
            in2 => \N__18729\,
            in3 => \N__20754\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIOAVU1_1_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20847\,
            in1 => \N__18735\,
            in2 => \N__18762\,
            in3 => \N__22283\,
            lcout => \b2v_inst200.un25_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNID13N_1_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18725\,
            in1 => \N__18755\,
            in2 => \_gnd_net_\,
            in3 => \N__22611\,
            lcout => \b2v_inst200.un2_count_1_axb_1\,
            ltout => \b2v_inst200.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_1_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18759\,
            in3 => \N__22282\,
            lcout => \b2v_inst200.count_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9S71_0_16_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__18744\,
            in1 => \N__20975\,
            in2 => \N__20954\,
            in3 => \N__22613\,
            lcout => \b2v_inst200.un25_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_1_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20768\,
            in2 => \_gnd_net_\,
            in3 => \N__22284\,
            lcout => \b2v_inst200.count_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36800\,
            ce => \N__22541\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3T051_3_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18818\,
            in1 => \N__20725\,
            in2 => \_gnd_net_\,
            in3 => \N__22617\,
            lcout => \b2v_inst200.un2_count_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_3_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20727\,
            lcout => \b2v_inst200.count_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36755\,
            ce => \N__22539\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73351_0_5_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000101"
        )
    port map (
            in0 => \N__20889\,
            in1 => \N__22621\,
            in2 => \N__18972\,
            in3 => \N__20685\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIUF4N4_3_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18810\,
            in1 => \N__18768\,
            in2 => \N__18717\,
            in3 => \N__18792\,
            lcout => \b2v_inst200.un25_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3T051_0_3_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000111"
        )
    port map (
            in0 => \N__20726\,
            in1 => \N__22619\,
            in2 => \N__18822\,
            in3 => \N__20709\,
            lcout => \b2v_inst200.un25_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_13_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20805\,
            lcout => \b2v_inst200.count_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36755\,
            ce => \N__22539\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50P71_13_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20803\,
            in1 => \N__18800\,
            in2 => \_gnd_net_\,
            in3 => \N__22618\,
            lcout => \b2v_inst200.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50P71_0_13_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100111"
        )
    port map (
            in0 => \N__22620\,
            in1 => \N__20804\,
            in2 => \N__18804\,
            in3 => \N__20789\,
            lcout => \b2v_inst200.un25_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_12_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36719\,
            ce => \N__22538\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_9_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36719\,
            ce => \N__22538\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIFF751_9_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22623\,
            in1 => \N__18779\,
            in2 => \_gnd_net_\,
            in3 => \N__20863\,
            lcout => \b2v_inst200.un2_count_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3TN71_12_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18786\,
            in1 => \N__20822\,
            in2 => \_gnd_net_\,
            in3 => \N__22625\,
            lcout => \b2v_inst200.countZ0Z_12\,
            ltout => \b2v_inst200.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIFF751_0_9_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__22626\,
            in1 => \N__18780\,
            in2 => \N__18771\,
            in3 => \N__20864\,
            lcout => \b2v_inst200.un25_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73351_5_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18968\,
            in1 => \N__22622\,
            in2 => \_gnd_net_\,
            in3 => \N__20683\,
            lcout => \b2v_inst200.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_5_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20684\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36719\,
            ce => \N__22538\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QM71_11_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22239\,
            in1 => \N__22250\,
            in2 => \_gnd_net_\,
            in3 => \N__22624\,
            lcout => \b2v_inst200.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI1ENE_15_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19278\,
            in1 => \N__18921\,
            in2 => \_gnd_net_\,
            in3 => \N__18935\,
            lcout => \b2v_inst16.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_15_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36872\,
            ce => \N__19277\,
            sr => \N__19146\
        );

    \b2v_inst16.count_RNIT7LE_13_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18894\,
            in1 => \N__18876\,
            in2 => \_gnd_net_\,
            in3 => \N__19271\,
            lcout => \b2v_inst16.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_13_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18893\,
            lcout => \b2v_inst16.count_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36872\,
            ce => \N__19277\,
            sr => \N__19146\
        );

    \b2v_inst16.count_RNIVAME_14_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18843\,
            in1 => \N__18828\,
            in2 => \_gnd_net_\,
            in3 => \N__19272\,
            lcout => \b2v_inst16.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_14_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18842\,
            lcout => \b2v_inst16.count_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36872\,
            ce => \N__19277\,
            sr => \N__19146\
        );

    \b2v_inst200.count_RNI1QV41_2_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22206\,
            in1 => \N__22191\,
            in2 => \_gnd_net_\,
            in3 => \N__22615\,
            lcout => \b2v_inst200.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50251_4_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22616\,
            in1 => \N__22164\,
            in2 => \_gnd_net_\,
            in3 => \N__22179\,
            lcout => \b2v_inst200.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_2_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19332\,
            lcout => \b2v_inst16.count_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36965\,
            ce => \N__19257\,
            sr => \N__19145\
        );

    \b2v_inst16.count_6_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19304\,
            lcout => \b2v_inst16.count_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36965\,
            ce => \N__19257\,
            sr => \N__19145\
        );

    \b2v_inst36.curr_state_0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__23150\,
            in1 => \N__23021\,
            in2 => \N__19082\,
            in3 => \N__23072\,
            lcout => \b2v_inst36.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36873\,
            ce => \N__27543\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100010000"
        )
    port map (
            in0 => \N__23020\,
            in1 => \N__19073\,
            in2 => \N__23082\,
            in3 => \N__23151\,
            lcout => \b2v_inst36.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36873\,
            ce => \N__27543\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m6_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110010"
        )
    port map (
            in0 => \N__23153\,
            in1 => \N__23016\,
            in2 => \N__23086\,
            in3 => \N__19072\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIU72Q_1_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19095\,
            in2 => \N__19089\,
            in3 => \N__28330\,
            lcout => \b2v_inst36.curr_stateZ0Z_1\,
            ltout => \b2v_inst36.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m4_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000001000"
        )
    port map (
            in0 => \N__23152\,
            in1 => \N__23022\,
            in2 => \N__19086\,
            in3 => \N__19071\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIT62Q_0_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18981\,
            in2 => \N__18975\,
            in3 => \N__28329\,
            lcout => \b2v_inst36.curr_stateZ0Z_0\,
            ltout => \b2v_inst36.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIRQCA_0_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__23154\,
            in1 => \N__28343\,
            in2 => \N__19563\,
            in3 => \N__23067\,
            lcout => \b2v_inst36.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__23068\,
            in1 => \_gnd_net_\,
            in2 => \N__23029\,
            in3 => \N__23149\,
            lcout => \b2v_inst36.DSW_PWROK_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36873\,
            ce => \N__27543\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI5MK6V3_11_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19350\,
            in1 => \N__28545\,
            in2 => \N__26556\,
            in3 => \N__21125\,
            lcout => \b2v_inst11.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_11_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26552\,
            lcout => \b2v_inst11.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37071\,
            ce => \N__28532\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_10_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26547\,
            in2 => \_gnd_net_\,
            in3 => \N__21141\,
            lcout => \b2v_inst11.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37071\,
            ce => \N__28532\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIS7D3V3_10_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28544\,
            in1 => \N__19344\,
            in2 => \N__26554\,
            in3 => \N__21140\,
            lcout => \b2v_inst11.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI7PL6V3_12_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28546\,
            in1 => \N__19338\,
            in2 => \N__26555\,
            in3 => \N__21110\,
            lcout => \b2v_inst11.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_12_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21114\,
            in3 => \N__26548\,
            lcout => \b2v_inst11.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37071\,
            ce => \N__28532\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIJMQ2V3_9_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28543\,
            in1 => \N__24795\,
            in2 => \N__26553\,
            in3 => \N__24806\,
            lcout => \b2v_inst11.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI74K2V3_3_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19659\,
            in1 => \N__28533\,
            in2 => \N__21012\,
            in3 => \N__26523\,
            lcout => \b2v_inst11.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_3_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21011\,
            lcout => \b2v_inst11.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37007\,
            ce => \N__28547\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_13_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26528\,
            lcout => \b2v_inst11.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37007\,
            ce => \N__28547\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNID2P6V3_15_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__26526\,
            in1 => \N__22938\,
            in2 => \N__28551\,
            in3 => \N__22949\,
            lcout => \b2v_inst11.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_14_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26529\,
            lcout => \b2v_inst11.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37007\,
            ce => \N__28547\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIBVN6V3_14_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__26525\,
            in1 => \N__19653\,
            in2 => \N__28550\,
            in3 => \N__21263\,
            lcout => \b2v_inst11.count_offZ0Z_14\,
            ltout => \b2v_inst11.count_offZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_15_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21098\,
            in1 => \N__22905\,
            in2 => \N__19644\,
            in3 => \N__21251\,
            lcout => \b2v_inst11.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI9SM6V3_13_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__26524\,
            in1 => \N__19641\,
            in2 => \N__28549\,
            in3 => \N__21083\,
            lcout => \b2v_inst11.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_1_cry_15_c_RNI9STGK62_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__19635\,
            in1 => \N__19948\,
            in2 => \N__19625\,
            in3 => \N__19596\,
            lcout => \b2v_inst11.N_6\,
            ltout => \b2v_inst11.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__19907\,
            in1 => \N__35808\,
            in2 => \N__19566\,
            in3 => \N__19895\,
            lcout => \b2v_inst11.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37001\,
            ce => 'H',
            sr => \N__19920\
        );

    \b2v_inst11.pwm_out_RNINR3DL62_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__27566\,
            in1 => \N__19908\,
            in2 => \N__19899\,
            in3 => \N__19884\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_en_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27564\,
            in2 => \_gnd_net_\,
            in3 => \N__21054\,
            lcout => \b2v_inst200.count_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIV6I72_0_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19815\,
            lcout => \b2v_inst16.delayed_vddq_pwrgd_en\,
            ltout => \b2v_inst16.delayed_vddq_pwrgd_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_RNIPAU73_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011111111"
        )
    port map (
            in0 => \N__20485\,
            in1 => \N__20442\,
            in2 => \N__19851\,
            in3 => \N__26784\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIBO6I1_0_0_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19830\,
            in2 => \_gnd_net_\,
            in3 => \N__20484\,
            lcout => \b2v_inst16.N_268\,
            ltout => \b2v_inst16.N_268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI35HL1_0_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19809\,
            in3 => \N__28389\,
            lcout => \b2v_inst16.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_RNO_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21452\,
            in1 => \N__21467\,
            in2 => \N__21438\,
            in3 => \N__21482\,
            lcout => \b2v_inst20.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_RNO_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21548\,
            in1 => \N__21533\,
            in2 => \N__21519\,
            in3 => \N__21500\,
            lcout => \b2v_inst20.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_0_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__20091\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \b2v_inst11.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31582\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23850\,
            in2 => \N__19970\,
            in3 => \N__23877\,
            lcout => \G_2848\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_0\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19966\,
            in2 => \N__23586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23878\,
            in2 => \N__23571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23556\,
            in2 => \N__23885\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23544\,
            in2 => \N__19971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_s_6_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23532\,
            in2 => \_gnd_net_\,
            in3 => \N__19953\,
            lcout => \b2v_inst11.mult1_un166_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27255\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21708\,
            in2 => \N__20120\,
            in3 => \N__20139\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20116\,
            in2 => \N__20103\,
            in3 => \N__20136\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20184\,
            in2 => \N__20241\,
            in3 => \N__20133\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20229\,
            in2 => \N__20192\,
            in3 => \N__20130\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23749\,
            in1 => \N__20220\,
            in2 => \N__20121\,
            in3 => \N__20127\,
            lcout => \b2v_inst11.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20211\,
            in3 => \N__20124\,
            lcout => \b2v_inst11.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20183\,
            lcout => \b2v_inst11.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27222\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25092\,
            in2 => \N__20162\,
            in3 => \N__20094\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20158\,
            in2 => \N__20340\,
            in3 => \N__20232\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20608\,
            in2 => \N__20316\,
            in3 => \N__20223\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20292\,
            in2 => \N__20615\,
            in3 => \N__20214\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20188\,
            in1 => \N__20658\,
            in2 => \N__20163\,
            in3 => \N__20202\,
            lcout => \b2v_inst11.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20640\,
            in2 => \_gnd_net_\,
            in3 => \N__20199\,
            lcout => \b2v_inst11.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20607\,
            lcout => \b2v_inst11.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27110\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21690\,
            in2 => \N__21731\,
            in3 => \N__20145\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21727\,
            in2 => \N__21678\,
            in3 => \N__20142\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21651\,
            in2 => \N__21761\,
            in3 => \N__20280\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21757\,
            in2 => \N__21897\,
            in3 => \N__20277\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20415\,
            in1 => \N__21831\,
            in2 => \N__21732\,
            in3 => \N__20274\,
            lcout => \b2v_inst11.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21792\,
            in3 => \N__20271\,
            lcout => \b2v_inst11.mult1_un117_sum_s_8\,
            ltout => \b2v_inst11.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20268\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27146\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20346\,
            in2 => \N__20378\,
            in3 => \N__20265\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20374\,
            in2 => \N__20262\,
            in3 => \N__20253\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20250\,
            in2 => \N__20423\,
            in3 => \N__20244\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20419\,
            in2 => \N__20397\,
            in3 => \N__20388\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20572\,
            in1 => \N__20385\,
            in2 => \N__20379\,
            in3 => \N__20361\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20358\,
            in3 => \N__20349\,
            lcout => \b2v_inst11.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27186\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21702\,
            in2 => \N__20546\,
            in3 => \N__20328\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20542\,
            in2 => \N__20325\,
            in3 => \N__20304\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20568\,
            in2 => \N__20301\,
            in3 => \N__20283\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20664\,
            in2 => \N__20576\,
            in3 => \N__20649\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20603\,
            in1 => \N__20646\,
            in2 => \N__20547\,
            in3 => \N__20631\,
            lcout => \b2v_inst11.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20628\,
            in3 => \N__20619\,
            lcout => \b2v_inst11.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20567\,
            lcout => \b2v_inst11.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111000100"
        )
    port map (
            in0 => \N__20529\,
            in1 => \N__20508\,
            in2 => \N__20496\,
            in3 => \N__20435\,
            lcout => \b2v_inst16.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73Q71_14_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22609\,
            in1 => \N__22227\,
            in2 => \_gnd_net_\,
            in3 => \N__22212\,
            lcout => \b2v_inst200.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI96451_6_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22685\,
            in1 => \N__22674\,
            in2 => \_gnd_net_\,
            in3 => \N__22606\,
            lcout => \b2v_inst200.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9551_7_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22607\,
            in1 => \N__22656\,
            in2 => \_gnd_net_\,
            in3 => \N__22667\,
            lcout => \b2v_inst200.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDCT71_17_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20919\,
            in1 => \N__20934\,
            in2 => \_gnd_net_\,
            in3 => \N__22610\,
            lcout => \b2v_inst200.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_0_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__22287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22314\,
            lcout => OPEN,
            ltout => \b2v_inst200.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_0_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22257\,
            in2 => \N__20772\,
            in3 => \N__22605\,
            lcout => \b2v_inst200.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIOMPC1_10_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__22608\,
            in1 => \_gnd_net_\,
            in2 => \N__22635\,
            in3 => \N__22650\,
            lcout => \b2v_inst200.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_1_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22285\,
            in2 => \N__20769\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20753\,
            in2 => \_gnd_net_\,
            in3 => \N__20736\,
            lcout => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_1\,
            carryout => \b2v_inst200.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20733\,
            in2 => \_gnd_net_\,
            in3 => \N__20712\,
            lcout => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_2\,
            carryout => \b2v_inst200.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20708\,
            in2 => \_gnd_net_\,
            in3 => \N__20694\,
            lcout => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_3\,
            carryout => \b2v_inst200.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20691\,
            in2 => \_gnd_net_\,
            in3 => \N__20670\,
            lcout => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_4\,
            carryout => \b2v_inst200.un2_count_1_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22339\,
            in1 => \N__22457\,
            in2 => \_gnd_net_\,
            in3 => \N__20667\,
            lcout => \b2v_inst200.count_1_6\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_5_cZ0\,
            carryout => \b2v_inst200.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20888\,
            in2 => \_gnd_net_\,
            in3 => \N__20877\,
            lcout => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_6\,
            carryout => \b2v_inst200.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22340\,
            in1 => \N__22008\,
            in2 => \_gnd_net_\,
            in3 => \N__20874\,
            lcout => \b2v_inst200.count_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_7\,
            carryout => \b2v_inst200.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20871\,
            in2 => \_gnd_net_\,
            in3 => \N__20853\,
            lcout => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22341\,
            in1 => \N__22403\,
            in2 => \_gnd_net_\,
            in3 => \N__20850\,
            lcout => \b2v_inst200.count_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_9\,
            carryout => \b2v_inst200.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22355\,
            in1 => \N__20843\,
            in2 => \_gnd_net_\,
            in3 => \N__20832\,
            lcout => \b2v_inst200.count_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_10\,
            carryout => \b2v_inst200.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20829\,
            in2 => \_gnd_net_\,
            in3 => \N__20814\,
            lcout => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_11\,
            carryout => \b2v_inst200.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20811\,
            in2 => \_gnd_net_\,
            in3 => \N__20793\,
            lcout => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_12\,
            carryout => \b2v_inst200.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20790\,
            in2 => \_gnd_net_\,
            in3 => \N__20775\,
            lcout => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_13\,
            carryout => \b2v_inst200.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_14_c_RNI96R71_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22020\,
            in3 => \N__20988\,
            lcout => \b2v_inst200.un2_count_1_cry_14_c_RNI96RZ0Z71\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_14\,
            carryout => \b2v_inst200.un2_count_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22342\,
            in1 => \N__20985\,
            in2 => \_gnd_net_\,
            in3 => \N__20958\,
            lcout => \b2v_inst200.count_1_16\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_15\,
            carryout => \b2v_inst200.un2_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__20955\,
            in1 => \N__22344\,
            in2 => \_gnd_net_\,
            in3 => \N__20937\,
            lcout => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_17_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20933\,
            lcout => \b2v_inst200.count_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36810\,
            ce => \N__22542\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21049\,
            in2 => \_gnd_net_\,
            in3 => \N__22343\,
            lcout => \b2v_inst200.N_282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI_1_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21328\,
            lcout => \b2v_inst200.N_2989_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m8_i_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111100"
        )
    port map (
            in0 => \N__21307\,
            in1 => \N__21350\,
            in2 => \N__21335\,
            in3 => \N__27762\,
            lcout => OPEN,
            ltout => \b2v_inst200.N_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI26MQ4_1_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__28320\,
            in1 => \_gnd_net_\,
            in2 => \N__20910\,
            in3 => \N__21294\,
            lcout => \b2v_inst200.curr_stateZ0Z_1\,
            ltout => \b2v_inst200.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110101"
        )
    port map (
            in0 => \N__21308\,
            in1 => \N__20907\,
            in2 => \N__20892\,
            in3 => \N__27761\,
            lcout => \b2v_inst200.m6_i_0\,
            ltout => \b2v_inst200.m6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__21050\,
            in1 => \_gnd_net_\,
            in2 => \N__21063\,
            in3 => \N__22354\,
            lcout => OPEN,
            ltout => \b2v_inst200.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI19645_0_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21021\,
            in2 => \N__21060\,
            in3 => \N__28319\,
            lcout => \b2v_inst200.curr_stateZ0Z_0\,
            ltout => \b2v_inst200.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21057\,
            in3 => \N__21176\,
            lcout => \N_411\,
            ltout => \N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_0_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22356\,
            in2 => \N__21030\,
            in3 => \N__21027\,
            lcout => \b2v_inst200.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36823\,
            ce => \N__27544\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22856\,
            in2 => \N__22901\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22842\,
            in3 => \N__21015\,
            lcout => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_1\,
            carryout => \b2v_inst11.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23201\,
            in3 => \N__20997\,
            lcout => \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_2\,
            carryout => \b2v_inst11.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22992\,
            in3 => \N__20994\,
            lcout => \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_3\,
            carryout => \b2v_inst11.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23361\,
            in3 => \N__20991\,
            lcout => \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_4\,
            carryout => \b2v_inst11.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23310\,
            in3 => \N__21153\,
            lcout => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_5\,
            carryout => \b2v_inst11.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24609\,
            in3 => \N__21150\,
            lcout => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_6\,
            carryout => \b2v_inst11.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24525\,
            in2 => \_gnd_net_\,
            in3 => \N__21147\,
            lcout => \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_7\,
            carryout => \b2v_inst11.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21198\,
            in3 => \N__21144\,
            lcout => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21212\,
            in3 => \N__21129\,
            lcout => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_9\,
            carryout => \b2v_inst11.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21225\,
            in3 => \N__21117\,
            lcout => \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_10\,
            carryout => \b2v_inst11.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21237\,
            in3 => \N__21102\,
            lcout => \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_11\,
            carryout => \b2v_inst11.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21099\,
            in3 => \N__21075\,
            lcout => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_12\,
            carryout => \b2v_inst11.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21072\,
            in3 => \N__21255\,
            lcout => \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_13\,
            carryout => \b2v_inst11.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21252\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21240\,
            lcout => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_9_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21236\,
            in1 => \N__21224\,
            in2 => \N__21213\,
            in3 => \N__21197\,
            lcout => \b2v_inst11.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI37MQ4_2_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__21159\,
            in1 => \N__21183\,
            in2 => \_gnd_net_\,
            in3 => \N__28257\,
            lcout => \b2v_inst200.curr_state_i_2\,
            ltout => \b2v_inst200.curr_state_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_ATP_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__21395\,
            in1 => \_gnd_net_\,
            in2 => \N__21186\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.HDA_SDO_ATP_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36996\,
            ce => \N__27536\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101010"
        )
    port map (
            in0 => \N__21358\,
            in1 => \N__21394\,
            in2 => \N__27782\,
            in3 => \N__21381\,
            lcout => \b2v_inst200.i4_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI_0_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21314\,
            in2 => \_gnd_net_\,
            in3 => \N__21177\,
            lcout => \b2v_inst200.N_205\,
            ltout => \b2v_inst200.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_2_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100010001"
        )
    port map (
            in0 => \N__21359\,
            in1 => \N__21379\,
            in2 => \N__21162\,
            in3 => \N__27778\,
            lcout => \b2v_inst200.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36996\,
            ce => \N__27536\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_RNO_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21573\,
            in1 => \N__21615\,
            in2 => \N__21597\,
            in3 => \N__21633\,
            lcout => \b2v_inst20.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_ATP_RNILDHE_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__28259\,
            in1 => \N__21405\,
            in2 => \N__21399\,
            in3 => \N__21380\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_1_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011111100"
        )
    port map (
            in0 => \N__27777\,
            in1 => \N__21360\,
            in2 => \N__21339\,
            in3 => \N__21315\,
            lcout => \b2v_inst200.curr_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36996\,
            ce => \N__27536\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25013\,
            in2 => \N__23178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \b2v_inst20.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24969\,
            in2 => \_gnd_net_\,
            in3 => \N__21282\,
            lcout => \b2v_inst20.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_1\,
            carryout => \b2v_inst20.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24939\,
            in2 => \_gnd_net_\,
            in3 => \N__21279\,
            lcout => \b2v_inst20.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_2\,
            carryout => \b2v_inst20.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24909\,
            in2 => \_gnd_net_\,
            in3 => \N__21276\,
            lcout => \b2v_inst20.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_3\,
            carryout => \b2v_inst20.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23256\,
            in3 => \N__21273\,
            lcout => \b2v_inst20.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_4\,
            carryout => \b2v_inst20.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23226\,
            in2 => \_gnd_net_\,
            in3 => \N__21270\,
            lcout => \b2v_inst20.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_5\,
            carryout => \b2v_inst20.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_7_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22826\,
            in2 => \_gnd_net_\,
            in3 => \N__21267\,
            lcout => \b2v_inst20.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_6\,
            carryout => \b2v_inst20.counter_1_cry_7\,
            clk => \N__37072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_8_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21483\,
            in2 => \_gnd_net_\,
            in3 => \N__21471\,
            lcout => \b2v_inst20.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_7\,
            carryout => \b2v_inst20.counter_1_cry_8\,
            clk => \N__37072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_9_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21468\,
            in2 => \_gnd_net_\,
            in3 => \N__21456\,
            lcout => \b2v_inst20.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \b2v_inst20.counter_1_cry_9\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_10_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21453\,
            in2 => \_gnd_net_\,
            in3 => \N__21441\,
            lcout => \b2v_inst20.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_9\,
            carryout => \b2v_inst20.counter_1_cry_10\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_11_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21437\,
            in2 => \_gnd_net_\,
            in3 => \N__21423\,
            lcout => \b2v_inst20.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_10\,
            carryout => \b2v_inst20.counter_1_cry_11\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_12_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23400\,
            in2 => \_gnd_net_\,
            in3 => \N__21420\,
            lcout => \b2v_inst20.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_11\,
            carryout => \b2v_inst20.counter_1_cry_12\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_13_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23427\,
            in2 => \_gnd_net_\,
            in3 => \N__21417\,
            lcout => \b2v_inst20.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_12\,
            carryout => \b2v_inst20.counter_1_cry_13\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_14_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23414\,
            in2 => \_gnd_net_\,
            in3 => \N__21414\,
            lcout => \b2v_inst20.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_13\,
            carryout => \b2v_inst20.counter_1_cry_14\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_15_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23439\,
            in2 => \_gnd_net_\,
            in3 => \N__21411\,
            lcout => \b2v_inst20.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_14\,
            carryout => \b2v_inst20.counter_1_cry_15\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_16_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23496\,
            in2 => \_gnd_net_\,
            in3 => \N__21408\,
            lcout => \b2v_inst20.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_15\,
            carryout => \b2v_inst20.counter_1_cry_16\,
            clk => \N__36997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_17_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23484\,
            in2 => \_gnd_net_\,
            in3 => \N__21558\,
            lcout => \b2v_inst20.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \b2v_inst20.counter_1_cry_17\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_18_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23471\,
            in2 => \_gnd_net_\,
            in3 => \N__21555\,
            lcout => \b2v_inst20.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_17\,
            carryout => \b2v_inst20.counter_1_cry_18\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_19_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23457\,
            in2 => \_gnd_net_\,
            in3 => \N__21552\,
            lcout => \b2v_inst20.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_18\,
            carryout => \b2v_inst20.counter_1_cry_19\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_20_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21549\,
            in2 => \_gnd_net_\,
            in3 => \N__21537\,
            lcout => \b2v_inst20.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_19\,
            carryout => \b2v_inst20.counter_1_cry_20\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_21_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21534\,
            in2 => \_gnd_net_\,
            in3 => \N__21522\,
            lcout => \b2v_inst20.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_20\,
            carryout => \b2v_inst20.counter_1_cry_21\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_22_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21518\,
            in2 => \_gnd_net_\,
            in3 => \N__21504\,
            lcout => \b2v_inst20.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_21\,
            carryout => \b2v_inst20.counter_1_cry_22\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_23_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21501\,
            in2 => \_gnd_net_\,
            in3 => \N__21489\,
            lcout => \b2v_inst20.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_22\,
            carryout => \b2v_inst20.counter_1_cry_23\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_24_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23652\,
            in2 => \_gnd_net_\,
            in3 => \N__21486\,
            lcout => \b2v_inst20.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_23\,
            carryout => \b2v_inst20.counter_1_cry_24\,
            clk => \N__37002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_25_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23621\,
            in2 => \_gnd_net_\,
            in3 => \N__21642\,
            lcout => \b2v_inst20.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \b2v_inst20.counter_1_cry_25\,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_26_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23639\,
            in2 => \_gnd_net_\,
            in3 => \N__21639\,
            lcout => \b2v_inst20.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_25\,
            carryout => \b2v_inst20.counter_1_cry_26\,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_27_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23606\,
            in2 => \_gnd_net_\,
            in3 => \N__21636\,
            lcout => \b2v_inst20.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_26\,
            carryout => \b2v_inst20.counter_1_cry_27\,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_28_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21632\,
            in2 => \_gnd_net_\,
            in3 => \N__21618\,
            lcout => \b2v_inst20.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_27\,
            carryout => \b2v_inst20.counter_1_cry_28\,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_29_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21614\,
            in2 => \_gnd_net_\,
            in3 => \N__21600\,
            lcout => \b2v_inst20.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_28\,
            carryout => \b2v_inst20.counter_1_cry_29\,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_30_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21593\,
            in2 => \_gnd_net_\,
            in3 => \N__21579\,
            lcout => \b2v_inst20.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_29\,
            carryout => \b2v_inst20.counter_1_cry_30\,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_31_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21572\,
            in2 => \_gnd_net_\,
            in3 => \N__21576\,
            lcout => \b2v_inst20.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_4_l_fx_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23819\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23748\,
            lcout => \b2v_inst11.mult1_un152_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23746\,
            lcout => \b2v_inst11.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27221\,
            lcout => \b2v_inst11.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_7_l_fx_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23747\,
            lcout => \b2v_inst11.mult1_un152_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31987\,
            lcout => \b2v_inst11.N_2943_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27147\,
            lcout => \b2v_inst11.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21875\,
            lcout => \b2v_inst11.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27090\,
            lcout => \b2v_inst11.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27068\,
            lcout => \b2v_inst11.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27086\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21684\,
            in2 => \N__21809\,
            in3 => \N__21669\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21805\,
            in2 => \N__21666\,
            in3 => \N__21645\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21909\,
            in2 => \N__21885\,
            in3 => \N__21888\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21884\,
            in2 => \N__21846\,
            in3 => \N__21825\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21753\,
            in1 => \N__21822\,
            in2 => \N__21810\,
            in3 => \N__21783\,
            lcout => \b2v_inst11.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21780\,
            in3 => \N__21765\,
            lcout => \b2v_inst11.mult1_un110_sum_s_8\,
            ltout => \b2v_inst11.mult1_un110_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21735\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23973\,
            in2 => \N__21989\,
            in3 => \N__21714\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21985\,
            in2 => \N__23898\,
            in3 => \N__21711\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24090\,
            in2 => \N__24147\,
            in3 => \N__22002\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24135\,
            in2 => \N__24098\,
            in3 => \N__21999\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22063\,
            in1 => \N__24126\,
            in2 => \N__21990\,
            in3 => \N__21996\,
            lcout => \b2v_inst11.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24117\,
            in3 => \N__21993\,
            lcout => \b2v_inst11.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24089\,
            lcout => \b2v_inst11.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27038\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27375\,
            in2 => \N__22037\,
            in3 => \N__21957\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22033\,
            in2 => \N__21954\,
            in3 => \N__21933\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22059\,
            in2 => \N__21930\,
            in3 => \N__21912\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22152\,
            in2 => \N__22067\,
            in3 => \N__22137\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22091\,
            in1 => \N__22134\,
            in2 => \N__22038\,
            in3 => \N__22116\,
            lcout => \b2v_inst11.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22113\,
            in3 => \N__22104\,
            lcout => \b2v_inst11.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22058\,
            lcout => \b2v_inst11.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI2KKU_15_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22603\,
            in1 => \N__22472\,
            in2 => \_gnd_net_\,
            in3 => \N__22444\,
            lcout => \b2v_inst200.un2_count_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_15_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => \N__22537\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_8_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => \N__22537\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDC651_8_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22416\,
            in1 => \N__22429\,
            in2 => \_gnd_net_\,
            in3 => \N__22602\,
            lcout => \b2v_inst200.un2_count_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI2KKU_0_15_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__22604\,
            in1 => \N__22473\,
            in2 => \N__22464\,
            in3 => \N__22445\,
            lcout => \b2v_inst200.un25_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDC651_0_8_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__22431\,
            in1 => \N__22415\,
            in2 => \N__22404\,
            in3 => \N__22601\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI5RUP8_8_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22386\,
            in1 => \N__22374\,
            in2 => \N__22368\,
            in3 => \N__22365\,
            lcout => \b2v_inst200.count_RNI5RUP8Z0Z_8\,
            ltout => \b2v_inst200.count_RNI5RUP8Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_0_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22290\,
            in3 => \N__22286\,
            lcout => \b2v_inst200.count_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36436\,
            ce => \N__22537\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_11_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22251\,
            lcout => \b2v_inst200.count_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_14_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22226\,
            lcout => \b2v_inst200.count_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_2_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22205\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_4_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22178\,
            lcout => \b2v_inst200.count_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_6_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22686\,
            lcout => \b2v_inst200.count_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_7_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22668\,
            lcout => \b2v_inst200.count_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_10_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22649\,
            lcout => \b2v_inst200.count_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36775\,
            ce => \N__22540\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_0_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24348\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_0_c_RNILCP9_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24275\,
            in2 => \_gnd_net_\,
            in3 => \N__22488\,
            lcout => \b2v_inst5.un2_count_1_cry_0_c_RNILCPZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_0\,
            carryout => \b2v_inst5.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_1_c_RNIMEQ9_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25656\,
            in2 => \_gnd_net_\,
            in3 => \N__22485\,
            lcout => \b2v_inst5.un2_count_1_cry_1_c_RNIMEQZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_1\,
            carryout => \b2v_inst5.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24288\,
            in2 => \_gnd_net_\,
            in3 => \N__22482\,
            lcout => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_2\,
            carryout => \b2v_inst5.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22739\,
            in2 => \_gnd_net_\,
            in3 => \N__22479\,
            lcout => \b2v_inst5.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_3\,
            carryout => \b2v_inst5.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_4_c_RNIPKT9_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25595\,
            in2 => \_gnd_net_\,
            in3 => \N__22476\,
            lcout => \b2v_inst5.un2_count_1_cry_4_c_RNIPKTZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_4\,
            carryout => \b2v_inst5.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_5_c_RNIQMU9_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25571\,
            in2 => \_gnd_net_\,
            in3 => \N__22713\,
            lcout => \b2v_inst5.un2_count_1_cry_5_c_RNIQMUZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_5\,
            carryout => \b2v_inst5.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_6_c_RNIROV9_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25449\,
            in2 => \_gnd_net_\,
            in3 => \N__22710\,
            lcout => \b2v_inst5.un2_count_1_cry_6_c_RNIROVZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_6\,
            carryout => \b2v_inst5.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22796\,
            in3 => \N__22707\,
            lcout => \b2v_inst5.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26028\,
            in2 => \_gnd_net_\,
            in3 => \N__22704\,
            lcout => \b2v_inst5.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_8\,
            carryout => \b2v_inst5.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25560\,
            in2 => \_gnd_net_\,
            in3 => \N__22701\,
            lcout => \b2v_inst5.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_9\,
            carryout => \b2v_inst5.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_10_c_RNI5KTC1_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25882\,
            in1 => \N__25482\,
            in2 => \_gnd_net_\,
            in3 => \N__22698\,
            lcout => \b2v_inst5.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_10\,
            carryout => \b2v_inst5.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_11_c_RNI76O2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24362\,
            in2 => \_gnd_net_\,
            in3 => \N__22695\,
            lcout => \b2v_inst5.un2_count_1_cry_11_c_RNI76OZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_11\,
            carryout => \b2v_inst5.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26163\,
            in3 => \N__22692\,
            lcout => \b2v_inst5.un2_count_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_12\,
            carryout => \b2v_inst5.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_13_c_RNI9AQ2_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24372\,
            in2 => \_gnd_net_\,
            in3 => \N__22689\,
            lcout => \b2v_inst5.un2_count_1_cry_13_c_RNI9AQZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_13\,
            carryout => \b2v_inst5.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_14_c_RNI9S1D1_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24438\,
            in1 => \N__25883\,
            in2 => \_gnd_net_\,
            in3 => \N__22812\,
            lcout => \b2v_inst5.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIH08H3_4_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22719\,
            in1 => \N__26250\,
            in2 => \_gnd_net_\,
            in3 => \N__22758\,
            lcout => \b2v_inst5.countZ0Z_4\,
            ltout => \b2v_inst5.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIU15T1_0_8_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__26252\,
            in1 => \N__22767\,
            in2 => \N__22809\,
            in3 => \N__22806\,
            lcout => \b2v_inst5.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_c_RNIPCCH3_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26104\,
            in1 => \N__22778\,
            in2 => \N__22797\,
            in3 => \N__25855\,
            lcout => \b2v_inst5.count_rst_6\,
            ltout => \b2v_inst5.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIU15T1_8_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26251\,
            in1 => \_gnd_net_\,
            in2 => \N__22800\,
            in3 => \N__22766\,
            lcout => \b2v_inst5.un2_count_1_axb_8\,
            ltout => \b2v_inst5.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_8_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26108\,
            in1 => \N__22779\,
            in2 => \N__22770\,
            in3 => \N__25857\,
            lcout => \b2v_inst5.count_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36822\,
            ce => \N__26294\,
            sr => \N__25991\
        );

    \b2v_inst5.un2_count_1_cry_3_c_RNIN23K1_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__25854\,
            in1 => \N__22751\,
            in2 => \N__22740\,
            in3 => \N__26103\,
            lcout => \b2v_inst5.count_rst_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_4_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__22752\,
            in1 => \N__22735\,
            in2 => \N__26109\,
            in3 => \N__25856\,
            lcout => \b2v_inst5.count_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36822\,
            ce => \N__26294\,
            sr => \N__25991\
        );

    \b2v_inst5.count_RNIL9B73_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__25853\,
            in1 => \N__24484\,
            in2 => \_gnd_net_\,
            in3 => \N__26102\,
            lcout => \b2v_inst5.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22872\,
            in2 => \_gnd_net_\,
            in3 => \N__26473\,
            lcout => \b2v_inst11.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36639\,
            ce => \N__28531\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_2_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22923\,
            lcout => \b2v_inst11.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36639\,
            ce => \N__28531\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_0_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26472\,
            lcout => \b2v_inst11.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36639\,
            ce => \N__28531\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI51J2V3_2_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22929\,
            in1 => \N__28502\,
            in2 => \N__26522\,
            in3 => \N__22922\,
            lcout => \b2v_inst11.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI5TD0V3_0_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__22899\,
            in1 => \N__28500\,
            in2 => \N__22914\,
            in3 => \N__26466\,
            lcout => \b2v_inst11.count_offZ0Z_0\,
            ltout => \b2v_inst11.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_1_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22875\,
            in3 => \N__22857\,
            lcout => \b2v_inst11.count_off_RNIZ0Z_1\,
            ltout => \b2v_inst11.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI6UD0V3_1_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22866\,
            in1 => \N__28501\,
            in2 => \N__22860\,
            in3 => \N__26467\,
            lcout => \b2v_inst11.count_offZ0Z_1\,
            ltout => \b2v_inst11.count_offZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_0_1_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23306\,
            in1 => \N__23360\,
            in2 => \N__22845\,
            in3 => \N__22841\,
            lcout => \b2v_inst11.un34_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_RNO_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__23167\,
            in1 => \N__23248\,
            in2 => \N__23225\,
            in3 => \N__22827\,
            lcout => \b2v_inst20.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_5_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000110"
        )
    port map (
            in0 => \N__23249\,
            in1 => \N__23265\,
            in2 => \N__26697\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst20.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_6_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__23221\,
            in1 => \N__26691\,
            in2 => \_gnd_net_\,
            in3 => \N__23235\,
            lcout => \b2v_inst20.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24605\,
            in1 => \N__22988\,
            in2 => \N__23205\,
            in3 => \N__24521\,
            lcout => \b2v_inst11.un34_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28258\,
            lcout => \SYNTHESIZED_WIRE_1keep_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__23168\,
            in1 => \N__25017\,
            in2 => \_gnd_net_\,
            in3 => \N__26692\,
            lcout => \b2v_inst20.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI3E27_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__23147\,
            in1 => \N__23091\,
            in2 => \_gnd_net_\,
            in3 => \N__23040\,
            lcout => \b2v_inst36.curr_state_RNI3E27Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI97L2V3_4_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22956\,
            in1 => \N__28526\,
            in2 => \N__22974\,
            in3 => \N__26531\,
            lcout => \b2v_inst11.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_4_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22970\,
            lcout => \b2v_inst11.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36891\,
            ce => \N__28548\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_15_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22950\,
            in2 => \_gnd_net_\,
            in3 => \N__26537\,
            lcout => \b2v_inst11.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36891\,
            ce => \N__28548\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_5_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23372\,
            lcout => \b2v_inst11.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36891\,
            ce => \N__28548\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIBAM2V3_5_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23382\,
            in1 => \N__28527\,
            in2 => \N__23376\,
            in3 => \N__26532\,
            lcout => \b2v_inst11.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_6_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__26535\,
            in1 => \_gnd_net_\,
            in2 => \N__23333\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36891\,
            ce => \N__28548\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIDDN2V3_6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23343\,
            in1 => \N__28525\,
            in2 => \N__23337\,
            in3 => \N__26530\,
            lcout => \b2v_inst11.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_7_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24632\,
            lcout => \b2v_inst11.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36891\,
            ce => \N__28548\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24984\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \b2v_inst20.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23286\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_0\,
            carryout => \b2v_inst20.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23277\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_1\,
            carryout => \b2v_inst20.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23388\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_2\,
            carryout => \b2v_inst20.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23445\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_3\,
            carryout => \b2v_inst20.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23517\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_4\,
            carryout => \b2v_inst20.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23592\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_5\,
            carryout => \b2v_inst20.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23505\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_6\,
            carryout => b2v_inst20_un4_counter_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23499\,
            lcout => \b2v_inst20_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_RNO_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23495\,
            in1 => \N__23483\,
            in2 => \N__23472\,
            in3 => \N__23456\,
            lcout => \b2v_inst20.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.G_149_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34240\,
            in2 => \_gnd_net_\,
            in3 => \N__26654\,
            lcout => \G_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_RNO_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23438\,
            in1 => \N__23426\,
            in2 => \N__23415\,
            in3 => \N__23399\,
            lcout => \b2v_inst20.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_rep1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__34241\,
            in1 => \_gnd_net_\,
            in2 => \N__26672\,
            in3 => \_gnd_net_\,
            lcout => \SYNTHESIZED_WIRE_1keep_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_RNO_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23651\,
            in1 => \N__23640\,
            in2 => \N__23625\,
            in3 => \N__23607\,
            lcout => \b2v_inst20.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31460\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25026\,
            in2 => \N__23990\,
            in3 => \N__23574\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23986\,
            in2 => \N__23832\,
            in3 => \N__23559\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23796\,
            in2 => \N__24020\,
            in3 => \N__23547\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24016\,
            in2 => \N__23778\,
            in3 => \N__23535\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23873\,
            in1 => \N__23709\,
            in2 => \N__23991\,
            in3 => \N__23523\,
            lcout => \b2v_inst11.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23676\,
            in3 => \N__23520\,
            lcout => \b2v_inst11.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_2_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31302\,
            in3 => \N__26813\,
            lcout => \b2v_inst11.N_366\,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25101\,
            in2 => \N__23841\,
            in3 => \N__23823\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23820\,
            in2 => \N__23805\,
            in3 => \N__23790\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23787\,
            in2 => \N__23765\,
            in3 => \N__23769\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23761\,
            in2 => \N__23721\,
            in3 => \N__23703\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__24012\,
            in1 => \N__23700\,
            in2 => \N__23685\,
            in3 => \N__23667\,
            lcout => \b2v_inst11.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23664\,
            in3 => \N__24030\,
            lcout => \b2v_inst11.mult1_un152_sum_s_8\,
            ltout => \b2v_inst11.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23994\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27315\,
            lcout => \b2v_inst11.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27339\,
            lcout => \b2v_inst11.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27360\,
            lcout => \b2v_inst11.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27039\,
            lcout => \b2v_inst11.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27786\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_6_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33879\,
            lcout => \b2v_inst11.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37063\,
            ce => \N__33837\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27359\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23907\,
            in2 => \N__24068\,
            in3 => \N__23889\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24064\,
            in2 => \N__24042\,
            in3 => \N__24138\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24186\,
            in2 => \N__24243\,
            in3 => \N__24129\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24231\,
            in2 => \N__24194\,
            in3 => \N__24120\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__24094\,
            in1 => \N__24222\,
            in2 => \N__24069\,
            in3 => \N__24108\,
            lcout => \b2v_inst11.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24213\,
            in3 => \N__24105\,
            lcout => \b2v_inst11.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24185\,
            lcout => \b2v_inst11.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27335\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24051\,
            in2 => \N__24164\,
            in3 => \N__24033\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24160\,
            in2 => \N__25176\,
            in3 => \N__24234\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25347\,
            in2 => \N__25437\,
            in3 => \N__24225\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25416\,
            in2 => \N__25355\,
            in3 => \N__24216\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__24190\,
            in1 => \N__25401\,
            in2 => \N__24165\,
            in3 => \N__24204\,
            lcout => \b2v_inst11.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25386\,
            in3 => \N__24201\,
            lcout => \b2v_inst11.mult1_un75_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25346\,
            lcout => \b2v_inst11.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_15_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24456\,
            lcout => \b2v_inst5.count_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36427\,
            ce => \N__26310\,
            sr => \N__25990\
        );

    \b2v_inst5.count_RNIL6AH3_6_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26266\,
            in1 => \N__24317\,
            in2 => \N__24306\,
            in3 => \N__25966\,
            lcout => \b2v_inst5.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_5_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__24336\,
            in1 => \_gnd_net_\,
            in2 => \N__25989\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36774\,
            ce => \N__26270\,
            sr => \N__25988\
        );

    \b2v_inst5.count_RNIJ39H3_5_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26265\,
            in1 => \N__24335\,
            in2 => \N__24327\,
            in3 => \N__25965\,
            lcout => \b2v_inst5.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_6_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25970\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24318\,
            lcout => \b2v_inst5.count_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36774\,
            ce => \N__26270\,
            sr => \N__25988\
        );

    \b2v_inst5.count_RNIH6CN3_13_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26118\,
            in1 => \_gnd_net_\,
            in2 => \N__26278\,
            in3 => \N__24294\,
            lcout => \b2v_inst5.countZ0Z_13\,
            ltout => \b2v_inst5.countZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_13_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__26136\,
            in1 => \N__25976\,
            in2 => \N__24297\,
            in3 => \N__26090\,
            lcout => \b2v_inst5.count_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36774\,
            ce => \N__26270\,
            sr => \N__25988\
        );

    \b2v_inst5.count_RNIFT6H3_3_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26264\,
            in1 => \N__25631\,
            in2 => \N__25614\,
            in3 => \N__25964\,
            lcout => \b2v_inst5.countZ0Z_3\,
            ltout => \b2v_inst5.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI_1_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25655\,
            in1 => \N__24279\,
            in2 => \N__24282\,
            in3 => \N__26155\,
            lcout => \b2v_inst5.un12_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIBN4H3_1_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__24263\,
            in1 => \N__26223\,
            in2 => \N__24252\,
            in3 => \N__25897\,
            lcout => \b2v_inst5.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_1_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25978\,
            in2 => \_gnd_net_\,
            in3 => \N__24264\,
            lcout => \b2v_inst5.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36512\,
            ce => \N__26287\,
            sr => \N__25977\
        );

    \b2v_inst5.count_12_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__24405\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25902\,
            lcout => \b2v_inst5.count_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36512\,
            ce => \N__26287\,
            sr => \N__25977\
        );

    \b2v_inst5.count_RNIF3BN3_12_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__25898\,
            in1 => \N__24404\,
            in2 => \N__24396\,
            in3 => \N__26256\,
            lcout => \b2v_inst5.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_14_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__24381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25903\,
            lcout => \b2v_inst5.count_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36512\,
            ce => \N__26287\,
            sr => \N__25977\
        );

    \b2v_inst5.count_RNIJ9DN3_14_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__24387\,
            in1 => \N__24380\,
            in2 => \N__25958\,
            in3 => \N__26257\,
            lcout => \b2v_inst5.countZ0Z_14\,
            ltout => \b2v_inst5.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIMP4T1_0_0_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__24434\,
            in1 => \N__24485\,
            in2 => \N__24366\,
            in3 => \N__24363\,
            lcout => \b2v_inst5.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24486\,
            in1 => \N__25979\,
            in2 => \_gnd_net_\,
            in3 => \N__26089\,
            lcout => \b2v_inst5.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36512\,
            ce => \N__26287\,
            sr => \N__25977\
        );

    \b2v_inst5.curr_state_1_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24420\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36744\,
            ce => \N__27539\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIRH7S1_0_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__24679\,
            in1 => \N__35827\,
            in2 => \N__27735\,
            in3 => \N__24666\,
            lcout => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0\,
            ltout => \b2v_inst5.curr_state_RNIRH7S1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_0_c_RNO_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24507\,
            in2 => \N__24351\,
            in3 => \N__24494\,
            lcout => \b2v_inst5.un2_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIKEUB2_1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24342\,
            in2 => \N__28325\,
            in3 => \N__24419\,
            lcout => \b2v_inst5.curr_stateZ0Z_1\,
            ltout => \b2v_inst5.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24510\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.curr_state_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIMP4T1_0_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__24506\,
            in1 => \_gnd_net_\,
            in2 => \N__24498\,
            in3 => \N__26221\,
            lcout => \b2v_inst5.count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24471\,
            in2 => \_gnd_net_\,
            in3 => \N__26081\,
            lcout => \N_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNILCEN3_15_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24465\,
            in1 => \N__26222\,
            in2 => \_gnd_net_\,
            in3 => \N__24449\,
            lcout => \b2v_inst5.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI65HI_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24705\,
            in2 => \N__28324\,
            in3 => \N__24411\,
            lcout => \b2v_inst5.curr_stateZ0Z_0\,
            ltout => \b2v_inst5.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m6_i_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__24664\,
            in1 => \N__27732\,
            in2 => \N__24423\,
            in3 => \N__24716\,
            lcout => \b2v_inst5.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__27731\,
            in1 => \_gnd_net_\,
            in2 => \N__24699\,
            in3 => \N__24663\,
            lcout => \RSMRSTn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36611\,
            ce => \N__27537\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__28790\,
            in1 => \N__24681\,
            in2 => \_gnd_net_\,
            in3 => \N__24715\,
            lcout => \b2v_inst5.m4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNID8DP1_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__27733\,
            in1 => \_gnd_net_\,
            in2 => \N__24698\,
            in3 => \N__24662\,
            lcout => \curr_state_RNID8DP1_0_0\,
            ltout => \curr_state_RNID8DP1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_0_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24680\,
            in2 => \N__24720\,
            in3 => \N__24717\,
            lcout => \b2v_inst5.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36611\,
            ce => \N__27537\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI65HI_0_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.N_2856_i\,
            ltout => \b2v_inst5.N_2856_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIVF6A1_0_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24665\,
            in1 => \N__27734\,
            in2 => \N__24645\,
            in3 => \N__28260\,
            lcout => \b2v_inst5.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIFGO2V3_7_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24642\,
            in1 => \N__28499\,
            in2 => \N__24633\,
            in3 => \N__26457\,
            lcout => \b2v_inst11.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_8_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24545\,
            lcout => \b2v_inst11.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36745\,
            ce => \N__28524\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_1_1_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24591\,
            in1 => \N__24579\,
            in2 => \N__24573\,
            in3 => \N__24558\,
            lcout => \b2v_inst11.count_off_RNI_1Z0Z_1\,
            ltout => \b2v_inst11.count_off_RNI_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI794G3_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__24822\,
            in1 => \N__32305\,
            in2 => \N__24552\,
            in3 => \N__28003\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNICMPB4_0_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28718\,
            in2 => \N__24549\,
            in3 => \N__30761\,
            lcout => \b2v_inst11.func_state_RNICMPB4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIHJP2V3_8_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24546\,
            in1 => \N__26460\,
            in2 => \N__24534\,
            in3 => \N__28498\,
            lcout => \b2v_inst11.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_9_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24813\,
            lcout => \b2v_inst11.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36745\,
            ce => \N__28524\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI6IFF4_0_1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__26628\,
            in1 => \N__37346\,
            in2 => \N__28719\,
            in3 => \N__24768\,
            lcout => \b2v_inst11.func_state_RNI6IFF4_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI05F44_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011111"
        )
    port map (
            in0 => \N__38982\,
            in1 => \N__26583\,
            in2 => \N__37357\,
            in3 => \N__33940\,
            lcout => \b2v_inst11.N_76\,
            ltout => \b2v_inst11.N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNII89R8_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24759\,
            in2 => \N__24783\,
            in3 => \N__24780\,
            lcout => \b2v_inst11.func_state_1_m2_1\,
            ltout => \b2v_inst11.func_state_1_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNICD8EB_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__24878\,
            in1 => \N__26773\,
            in2 => \N__24774\,
            in3 => \N__26732\,
            lcout => \b2v_inst11.func_state\,
            ltout => \b2v_inst11.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNITPVU_1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__38562\,
            in1 => \N__38725\,
            in2 => \N__24771\,
            in3 => \N__28240\,
            lcout => \b2v_inst11.N_339\,
            ltout => \b2v_inst11.N_339_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI6IFF4_1_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__37350\,
            in1 => \N__26627\,
            in2 => \N__24762\,
            in3 => \N__28714\,
            lcout => \b2v_inst11.func_state_RNI6IFF4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_RNIPUMD_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24753\,
            in1 => \N__24741\,
            in2 => \_gnd_net_\,
            in3 => \N__28241\,
            lcout => dsw_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__24879\,
            in1 => \N__26774\,
            in2 => \N__24888\,
            in3 => \N__26733\,
            lcout => \b2v_inst11.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI3NQD_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__28893\,
            in1 => \N__38983\,
            in2 => \N__38565\,
            in3 => \N__32266\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_51_and_i_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNILBJP_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__34261\,
            in1 => \N__28800\,
            in2 => \N__24870\,
            in3 => \N__28107\,
            lcout => \b2v_inst11.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.VCCST_EN_i_0_o3_0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111011111"
        )
    port map (
            in0 => \N__38554\,
            in1 => \N__34259\,
            in2 => \N__28115\,
            in3 => \N__28795\,
            lcout => \VCCST_EN_i_0_o3_0\,
            ltout => \VCCST_EN_i_0_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un1_vddq_en_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__24867\,
            in1 => \_gnd_net_\,
            in2 => \N__24849\,
            in3 => \_gnd_net_\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_en_0_x1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011001100"
        )
    port map (
            in0 => \N__38555\,
            in1 => \N__34258\,
            in2 => \N__38675\,
            in3 => \N__28794\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clk_en_0_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_en_0_ns_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24825\,
            in3 => \N__26673\,
            lcout => \b2v_inst11.count_clk_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38556\,
            in1 => \N__34260\,
            in2 => \N__38676\,
            in3 => \N__28796\,
            lcout => \b2v_inst11.N_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVT4P1_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__30767\,
            in1 => \N__37356\,
            in2 => \N__39060\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__34265\,
            in1 => \N__28116\,
            in2 => \N__38674\,
            in3 => \N__28809\,
            lcout => v5s_enn,
            ltout => \v5s_enn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIKAJP_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001110"
        )
    port map (
            in0 => \N__39001\,
            in1 => \N__32304\,
            in2 => \N__25020\,
            in3 => \N__31295\,
            lcout => \b2v_inst11.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__26669\,
            in1 => \_gnd_net_\,
            in2 => \N__25012\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst20.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__38528\,
            in1 => \N__38645\,
            in2 => \N__39085\,
            in3 => \N__34800\,
            lcout => \b2v_inst11.func_state_RNIDQ4A1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_RNO_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25002\,
            in1 => \N__24961\,
            in2 => \N__24938\,
            in3 => \N__24904\,
            lcout => \b2v_inst20.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__24978\,
            in1 => \_gnd_net_\,
            in2 => \N__24968\,
            in3 => \N__26670\,
            lcout => \b2v_inst20.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_3_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__24934\,
            in1 => \_gnd_net_\,
            in2 => \N__26680\,
            in3 => \N__24948\,
            lcout => \b2v_inst20.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_4_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__24905\,
            in1 => \N__24918\,
            in2 => \_gnd_net_\,
            in3 => \N__26671\,
            lcout => \b2v_inst20.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI498D2_5_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001101"
        )
    port map (
            in0 => \N__25041\,
            in1 => \N__39296\,
            in2 => \N__29087\,
            in3 => \N__29151\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_52_and_i_o3_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIB79JE_3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011101"
        )
    port map (
            in0 => \N__37345\,
            in1 => \N__30824\,
            in2 => \N__24891\,
            in3 => \N__25071\,
            lcout => \b2v_inst11.dutycycle_eena_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVK_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31179\,
            in1 => \N__35946\,
            in2 => \_gnd_net_\,
            in3 => \N__30534\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIRCVKZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNIKJFD2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__39057\,
            in1 => \N__38641\,
            in2 => \N__25044\,
            in3 => \N__25032\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_5_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__32303\,
            in1 => \N__39059\,
            in2 => \_gnd_net_\,
            in3 => \N__35947\,
            lcout => \b2v_inst11.N_236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI34G9_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32301\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINGLA1_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__38404\,
            in1 => \N__34251\,
            in2 => \N__25035\,
            in3 => \N__39056\,
            lcout => \b2v_inst11.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_9_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39058\,
            in1 => \N__38159\,
            in2 => \_gnd_net_\,
            in3 => \N__32302\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31296\,
            lcout => \b2v_inst11.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_14_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__26832\,
            in1 => \N__28860\,
            in2 => \N__34194\,
            in3 => \N__34036\,
            lcout => \b2v_inst11.dutycycle_RNI_14Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_13_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__28859\,
            in1 => \N__25050\,
            in2 => \N__34049\,
            in3 => \N__34189\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_3055_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIK9J85_5_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101100"
        )
    port map (
            in0 => \N__25059\,
            in1 => \N__26883\,
            in2 => \N__25083\,
            in3 => \N__36019\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_172_m3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIRO179_3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__26898\,
            in1 => \N__25080\,
            in2 => \N__25074\,
            in3 => \N__26952\,
            lcout => \b2v_inst11.un1_dutycycle_172_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_6_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38850\,
            in2 => \_gnd_net_\,
            in3 => \N__34032\,
            lcout => \b2v_inst11.N_19_i\,
            ltout => \b2v_inst11.N_19_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNII7Q52_5_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011110010"
        )
    port map (
            in0 => \N__38484\,
            in1 => \N__38615\,
            in2 => \N__25065\,
            in3 => \N__26877\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_172_m0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_5_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101100"
        )
    port map (
            in0 => \N__34823\,
            in1 => \N__28858\,
            in2 => \N__25062\,
            in3 => \N__36020\,
            lcout => \b2v_inst11.un1_dutycycle_172_m0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__38346\,
            in1 => \N__29276\,
            in2 => \_gnd_net_\,
            in3 => \N__28956\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_0_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__31454\,
            in1 => \N__31577\,
            in2 => \N__25053\,
            in3 => \N__37749\,
            lcout => \b2v_inst11.N_293_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_0_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__34024\,
            in1 => \N__25113\,
            in2 => \N__31583\,
            in3 => \N__31453\,
            lcout => \b2v_inst11.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_12_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29278\,
            in1 => \N__37747\,
            in2 => \N__28964\,
            in3 => \N__38347\,
            lcout => \b2v_inst11.g0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_12_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__37748\,
            in1 => \N__29279\,
            in2 => \N__38352\,
            in3 => \N__28960\,
            lcout => \b2v_inst11.g0_3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_13_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__34591\,
            in1 => \N__35084\,
            in2 => \N__37935\,
            in3 => \N__35193\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_a2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_15_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29331\,
            in1 => \N__38168\,
            in2 => \N__25107\,
            in3 => \N__37594\,
            lcout => \b2v_inst11.N_363\,
            ltout => \b2v_inst11.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_12_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__29277\,
            in1 => \_gnd_net_\,
            in2 => \N__25104\,
            in3 => \N__37746\,
            lcout => \b2v_inst11.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27248\,
            lcout => \b2v_inst11.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27185\,
            lcout => \b2v_inst11.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_8_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39055\,
            in1 => \N__37930\,
            in2 => \_gnd_net_\,
            in3 => \N__32310\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27288\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_3_sf_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29446\,
            lcout => \b2v_inst11.mult1_un54_sum_s_3_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27284\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25155\,
            in3 => \N__25146\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29394\,
            in3 => \N__25143\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30946\,
            in2 => \N__29460\,
            in3 => \N__25140\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30947\,
            in2 => \N__29493\,
            in3 => \N__25137\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27408\,
            in2 => \_gnd_net_\,
            in3 => \N__25134\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25131\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25261\,
            lcout => \b2v_inst11.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27438\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25262\,
            in2 => \N__25128\,
            in3 => \N__25116\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25272\,
            in2 => \N__25266\,
            in3 => \N__25248\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25198\,
            in2 => \N__25245\,
            in3 => \N__25236\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25233\,
            in2 => \N__25205\,
            in3 => \N__25227\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25321\,
            in1 => \N__25224\,
            in2 => \N__25185\,
            in3 => \N__25218\,
            lcout => \b2v_inst11.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25215\,
            in1 => \N__27407\,
            in2 => \N__25206\,
            in3 => \N__25209\,
            lcout => \b2v_inst11.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25197\,
            lcout => \b2v_inst11.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27311\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27423\,
            in2 => \N__25295\,
            in3 => \N__25167\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25291\,
            in2 => \N__25164\,
            in3 => \N__25428\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25317\,
            in2 => \N__25425\,
            in3 => \N__25410\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25407\,
            in2 => \N__25325\,
            in3 => \N__25395\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25351\,
            in1 => \N__25392\,
            in2 => \N__25296\,
            in3 => \N__25377\,
            lcout => \b2v_inst11.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25374\,
            in3 => \N__25365\,
            lcout => \b2v_inst11.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25316\,
            lcout => \b2v_inst11.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_c_RNI440L1_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__33137\,
            in1 => \N__29717\,
            in2 => \N__29738\,
            in3 => \N__29780\,
            lcout => \b2v_inst6.count_rst_11\,
            ltout => \b2v_inst6.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNINOEF5_3_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25508\,
            in2 => \N__25278\,
            in3 => \N__33450\,
            lcout => \b2v_inst6.un2_count_1_axb_3\,
            ltout => \b2v_inst6.un2_count_1_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__33140\,
            in1 => \N__29718\,
            in2 => \N__25275\,
            in3 => \N__29783\,
            lcout => \b2v_inst6.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36437\,
            ce => \N__33456\,
            sr => \N__33236\
        );

    \b2v_inst6.un2_count_1_cry_3_c_RNI561L1_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__29781\,
            in1 => \N__29672\,
            in2 => \N__29699\,
            in3 => \N__33138\,
            lcout => \b2v_inst6.count_rst_10\,
            ltout => \b2v_inst6.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIPRFF5_4_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33451\,
            in1 => \_gnd_net_\,
            in2 => \N__25518\,
            in3 => \N__25490\,
            lcout => \b2v_inst6.un2_count_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNINOEF5_0_3_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25515\,
            in1 => \N__25509\,
            in2 => \_gnd_net_\,
            in3 => \N__33453\,
            lcout => OPEN,
            ltout => \b2v_inst6.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIGKUUA_4_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__33452\,
            in1 => \N__25500\,
            in2 => \N__25494\,
            in3 => \N__25491\,
            lcout => \b2v_inst6.count_1_i_a3_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_4_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__29782\,
            in1 => \N__33139\,
            in2 => \N__29698\,
            in3 => \N__29673\,
            lcout => \b2v_inst6.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36437\,
            ce => \N__33456\,
            sr => \N__33236\
        );

    \b2v_inst5.count_7_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__25464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25963\,
            lcout => \b2v_inst5.count_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36834\,
            ce => \N__26276\,
            sr => \N__25998\
        );

    \b2v_inst5.count_RNID0AN3_11_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26262\,
            in1 => \N__25694\,
            in2 => \_gnd_net_\,
            in3 => \N__25711\,
            lcout => \b2v_inst5.un2_count_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_11_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36834\,
            ce => \N__26276\,
            sr => \N__25998\
        );

    \b2v_inst5.count_RNIN9BH3_7_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__25960\,
            in1 => \N__25470\,
            in2 => \N__26277\,
            in3 => \N__25463\,
            lcout => \b2v_inst5.countZ0Z_7\,
            ltout => \b2v_inst5.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNID0AN3_0_11_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__25712\,
            in1 => \N__25695\,
            in2 => \N__25683\,
            in3 => \N__26263\,
            lcout => \b2v_inst5.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_2_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25680\,
            lcout => \b2v_inst5.count_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36834\,
            ce => \N__26276\,
            sr => \N__25998\
        );

    \b2v_inst5.count_RNIDQ5H3_2_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__25679\,
            in1 => \N__26258\,
            in2 => \N__25665\,
            in3 => \N__25959\,
            lcout => \b2v_inst5.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_3_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25962\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25635\,
            lcout => \b2v_inst5.count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36834\,
            ce => \N__26276\,
            sr => \N__25998\
        );

    \b2v_inst5.count_RNI7BCA2_10_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26253\,
            in1 => \N__25524\,
            in2 => \_gnd_net_\,
            in3 => \N__26352\,
            lcout => \b2v_inst5.un2_count_1_axb_10\,
            ltout => \b2v_inst5.un2_count_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_10_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__25541\,
            in1 => \N__25975\,
            in2 => \N__25605\,
            in3 => \N__26086\,
            lcout => \b2v_inst5.count_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37014\,
            ce => \N__26306\,
            sr => \N__25980\
        );

    \b2v_inst5.count_RNI3QEK5_11_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25602\,
            in1 => \N__25596\,
            in2 => \N__25584\,
            in3 => \N__25575\,
            lcout => \b2v_inst5.un12_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_9_c_RNI4QLU3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__25556\,
            in1 => \N__25974\,
            in2 => \N__25542\,
            in3 => \N__26085\,
            lcout => \b2v_inst5.count_rst_4\,
            ltout => \b2v_inst5.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI7BCA2_0_10_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__26254\,
            in1 => \N__26351\,
            in2 => \N__26343\,
            in3 => \N__26016\,
            lcout => OPEN,
            ltout => \b2v_inst5.un12_clk_100khz_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI870S9_8_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26340\,
            in1 => \N__26328\,
            in2 => \N__26322\,
            in3 => \N__26319\,
            lcout => \b2v_inst5.N_1_i\,
            ltout => \b2v_inst5.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_9_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__26046\,
            in1 => \N__25981\,
            in2 => \N__26313\,
            in3 => \N__26017\,
            lcout => \b2v_inst5.count_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37014\,
            ce => \N__26306\,
            sr => \N__25980\
        );

    \b2v_inst5.count_RNIRFDH3_9_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26255\,
            in2 => \N__26172\,
            in3 => \N__25794\,
            lcout => \b2v_inst5.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_12_c_RNI7OVC1_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__26162\,
            in1 => \N__26135\,
            in2 => \N__25896\,
            in3 => \N__26087\,
            lcout => \b2v_inst5.count_rst_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_c_RNISC8K1_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__26088\,
            in1 => \N__26045\,
            in2 => \N__26027\,
            in3 => \N__25849\,
            lcout => \b2v_inst5.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un8_rsmrst_pwrgd_4_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25788\,
            in1 => \N__25773\,
            in2 => \N__25761\,
            in3 => \N__25740\,
            lcout => \SYNTHESIZED_WIRE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI_1_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27466\,
            lcout => \b2v_inst6.N_3011_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__25728\,
            in1 => \N__38730\,
            in2 => \N__26394\,
            in3 => \N__34817\,
            lcout => \b2v_inst6.N_192\,
            ltout => \b2v_inst6.N_192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__27645\,
            in1 => \_gnd_net_\,
            in2 => \N__26373\,
            in3 => \N__27861\,
            lcout => \b2v_inst6.N_241\,
            ltout => \b2v_inst6.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_1_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001111"
        )
    port map (
            in0 => \N__27467\,
            in1 => \_gnd_net_\,
            in2 => \N__26370\,
            in3 => \N__29820\,
            lcout => \b2v_inst6.curr_state_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36836\,
            ce => \N__27545\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIG8KAH_7_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__30153\,
            in1 => \N__29977\,
            in2 => \_gnd_net_\,
            in3 => \N__26361\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clk_RNIG8KAHZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNITV5AU_7_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27948\,
            in1 => \N__30440\,
            in2 => \N__26367\,
            in3 => \N__32296\,
            lcout => \b2v_inst11.count_clk_RNITV5AUZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI7SOFB_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__30479\,
            in1 => \N__27958\,
            in2 => \N__32946\,
            in3 => \N__29978\,
            lcout => \b2v_inst11.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIB2RFB_1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__27960\,
            in1 => \N__30151\,
            in2 => \_gnd_net_\,
            in3 => \N__30480\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIG510T_5_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32945\,
            in1 => \N__27947\,
            in2 => \N__26364\,
            in3 => \N__29979\,
            lcout => \b2v_inst11.count_clk_RNIG510TZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI7SOFB_0_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__27959\,
            in1 => \N__32944\,
            in2 => \_gnd_net_\,
            in3 => \N__30478\,
            lcout => \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1\,
            ltout => \b2v_inst11.count_clk_RNI7SOFB_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIG510T_0_7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__30152\,
            in1 => \N__27946\,
            in2 => \N__26355\,
            in3 => \N__29976\,
            lcout => \b2v_inst11.N_428\,
            ltout => \b2v_inst11.N_428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__39094\,
            in1 => \N__30441\,
            in2 => \N__26565\,
            in3 => \N__32297\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_332_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.N_224_i_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__39284\,
            in1 => \N__34771\,
            in2 => \N__38417\,
            in3 => \N__28328\,
            lcout => \b2v_inst11.N_224_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNILG61T1_5_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__28579\,
            in1 => \N__27990\,
            in2 => \N__26601\,
            in3 => \N__26562\,
            lcout => \b2v_inst11.count_clk_RNILG61T1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__39285\,
            in1 => \N__34769\,
            in2 => \N__38418\,
            in3 => \N__28326\,
            lcout => \b2v_inst11.N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_4_i_a2_sx_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__38722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39286\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_4_i_a2_sxZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_4_i_a2_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__28770\,
            in1 => \N__28142\,
            in2 => \N__26412\,
            in3 => \N__28085\,
            lcout => \b2v_inst11.N_417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28078\,
            in2 => \N__28146\,
            in3 => \N__28769\,
            lcout => rsmrstn,
            ltout => \rsmrstn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110011111"
        )
    port map (
            in0 => \N__38563\,
            in1 => \N__38718\,
            in2 => \N__26409\,
            in3 => \N__28327\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNI1EKN3_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010111"
        )
    port map (
            in0 => \N__34770\,
            in1 => \N__38564\,
            in2 => \N__38729\,
            in3 => \N__26406\,
            lcout => \b2v_inst11.N_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30749\,
            in1 => \N__28158\,
            in2 => \_gnd_net_\,
            in3 => \N__34059\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_331_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_fast_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26681\,
            lcout => \SYNTHESIZED_WIRE_1keep_3_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_2_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39053\,
            lcout => \b2v_inst11.func_state_RNI_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI5DLR_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000010001"
        )
    port map (
            in0 => \N__32276\,
            in1 => \N__38981\,
            in2 => \N__28734\,
            in3 => \N__30748\,
            lcout => \b2v_inst11.func_state_1_ss0_i_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__38724\,
            in1 => \N__39288\,
            in2 => \N__30377\,
            in3 => \N__32277\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__26777\,
            in1 => \N__26619\,
            in2 => \N__26613\,
            in3 => \N__26610\,
            lcout => \b2v_inst11.un1_func_state25_6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_0_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26597\,
            in1 => \N__28733\,
            in2 => \N__34818\,
            in3 => \N__32274\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_0_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110001"
        )
    port map (
            in0 => \N__32275\,
            in1 => \N__38980\,
            in2 => \N__26586\,
            in3 => \N__28892\,
            lcout => \b2v_inst11.func_state_1_m2s2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNITU8B9_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28017\,
            in1 => \N__26577\,
            in2 => \_gnd_net_\,
            in3 => \N__26571\,
            lcout => \b2v_inst11.func_state_1_m2_0\,
            ltout => \b2v_inst11.func_state_1_m2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIM28UB_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__26775\,
            in1 => \N__26747\,
            in2 => \N__26796\,
            in3 => \N__26734\,
            lcout => \b2v_inst11.func_stateZ0Z_0\,
            ltout => \b2v_inst11.func_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111001100"
        )
    port map (
            in0 => \N__39294\,
            in1 => \N__38560\,
            in2 => \N__26793\,
            in3 => \N__38693\,
            lcout => \b2v_inst11.g3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__38967\,
            in1 => \N__31395\,
            in2 => \_gnd_net_\,
            in3 => \N__32249\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26748\,
            in1 => \N__26790\,
            in2 => \N__26739\,
            in3 => \N__26776\,
            lcout => \b2v_inst11.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36980\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_1_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29224\,
            lcout => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI6M5R2_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010101"
        )
    port map (
            in0 => \N__26735\,
            in1 => \_gnd_net_\,
            in2 => \N__26715\,
            in3 => \N__37402\,
            lcout => \b2v_inst11.func_state_RNI6M5R2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_clk_100khz_52_and_i_a3_1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__38561\,
            in1 => \_gnd_net_\,
            in2 => \N__38717\,
            in3 => \N__34801\,
            lcout => \b2v_inst11.un1_clk_100khz_25_and_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111110000"
        )
    port map (
            in0 => \N__31297\,
            in1 => \N__26712\,
            in2 => \N__26706\,
            in3 => \N__31423\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_4_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26854\,
            in2 => \_gnd_net_\,
            in3 => \N__35002\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_3_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34362\,
            in2 => \_gnd_net_\,
            in3 => \N__38310\,
            lcout => \b2v_inst11.d_N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQH45K_5_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__34455\,
            in1 => \N__35789\,
            in2 => \N__33924\,
            in3 => \N__34466\,
            lcout => \b2v_inst11.dutycycleZ1Z_5\,
            ltout => \b2v_inst11.dutycycleZ1Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26838\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_5\,
            ltout => \b2v_inst11.dutycycle_RNI_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__38311\,
            in1 => \N__31463\,
            in2 => \N__26835\,
            in3 => \N__31532\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__31533\,
            in1 => \N__31424\,
            in2 => \N__26823\,
            in3 => \N__38312\,
            lcout => \b2v_inst11.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31425\,
            in1 => \N__31534\,
            in2 => \N__38343\,
            in3 => \N__26819\,
            lcout => \b2v_inst11.dutycycle_RNI_9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_2_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28902\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28666\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__28629\,
            in1 => \N__30637\,
            in2 => \N__32307\,
            in3 => \N__28901\,
            lcout => \b2v_inst11.N_159\,
            ltout => \b2v_inst11.N_159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26799\,
            in3 => \N__28670\,
            lcout => \b2v_inst11.N_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_1_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__28630\,
            in1 => \N__30438\,
            in2 => \N__28678\,
            in3 => \N__34183\,
            lcout => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__26855\,
            in1 => \N__38847\,
            in2 => \_gnd_net_\,
            in3 => \N__26892\,
            lcout => \b2v_inst11.dutycycle_RNI_11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_14_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__32284\,
            in1 => \_gnd_net_\,
            in2 => \N__39093\,
            in3 => \N__35211\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_10_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__35472\,
            in1 => \N__39012\,
            in2 => \_gnd_net_\,
            in3 => \N__32282\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_13_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__32283\,
            in1 => \_gnd_net_\,
            in2 => \N__39092\,
            in3 => \N__34605\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_0_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__32292\,
            in1 => \N__26946\,
            in2 => \N__31290\,
            in3 => \N__36175\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_172_m3_d_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111100001"
        )
    port map (
            in0 => \N__26931\,
            in1 => \N__26915\,
            in2 => \N__26886\,
            in3 => \N__30429\,
            lcout => \b2v_inst11.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_5_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__32294\,
            in1 => \N__26862\,
            in2 => \_gnd_net_\,
            in3 => \N__36177\,
            lcout => \b2v_inst11.dutycycle_RNIDQ4A1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__36176\,
            in1 => \N__27015\,
            in2 => \N__31291\,
            in3 => \N__32293\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_172_m4_rn_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQK9K2_0_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__32295\,
            in1 => \N__36178\,
            in2 => \N__26871\,
            in3 => \N__26868\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_172_m4_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI7FEU3_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__26861\,
            in1 => \N__27014\,
            in2 => \N__26955\,
            in3 => \N__30428\,
            lcout => \b2v_inst11.un1_dutycycle_172_m4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_16_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__26916\,
            in1 => \N__26939\,
            in2 => \N__34193\,
            in3 => \N__28861\,
            lcout => \b2v_inst11.N_3057_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_17_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__26940\,
            in1 => \N__28862\,
            in2 => \_gnd_net_\,
            in3 => \N__34187\,
            lcout => \b2v_inst11.N_3055_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_3_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__34388\,
            in1 => \_gnd_net_\,
            in2 => \N__38859\,
            in3 => \N__34986\,
            lcout => \b2v_inst11.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_2_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29241\,
            in2 => \_gnd_net_\,
            in3 => \N__38851\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5AV24_4_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__34976\,
            in1 => \N__37508\,
            in2 => \N__26925\,
            in3 => \N__37408\,
            lcout => \b2v_inst11.dutycycle_RNI5AV24Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31554\,
            in1 => \N__26922\,
            in2 => \N__34047\,
            in3 => \N__31449\,
            lcout => \b2v_inst11.g1_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111101"
        )
    port map (
            in0 => \N__26907\,
            in1 => \N__31552\,
            in2 => \N__31462\,
            in3 => \N__34188\,
            lcout => OPEN,
            ltout => \b2v_inst11.g2_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__29178\,
            in1 => \N__34978\,
            in2 => \N__26901\,
            in3 => \N__34387\,
            lcout => \b2v_inst11.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31448\,
            in1 => \N__31553\,
            in2 => \N__38858\,
            in3 => \N__29327\,
            lcout => \b2v_inst11.dutycycle_RNI_10Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__31555\,
            in1 => \N__34977\,
            in2 => \_gnd_net_\,
            in3 => \N__31444\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIPKS23_4_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__35799\,
            in1 => \N__36173\,
            in2 => \N__26997\,
            in3 => \N__27003\,
            lcout => \b2v_inst11.dutycycle_RNIPKS23Z0Z_4\,
            ltout => \b2v_inst11.dutycycle_RNIPKS23Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_4_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__26982\,
            in1 => \N__37361\,
            in2 => \N__27006\,
            in3 => \N__26996\,
            lcout => \b2v_inst11.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37069\,
            ce => 'H',
            sr => \N__36341\
        );

    \b2v_inst11.dutycycle_RNI_1_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__31443\,
            in1 => \N__31299\,
            in2 => \N__35009\,
            in3 => \N__36011\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08U_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31128\,
            in1 => \N__30969\,
            in2 => \_gnd_net_\,
            in3 => \N__36010\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIV08UZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIM7549_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__26995\,
            in1 => \N__26981\,
            in2 => \N__37362\,
            in3 => \N__26973\,
            lcout => \b2v_inst11.dutycycleZ0Z_6\,
            ltout => \b2v_inst11.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__38345\,
            in1 => \N__31442\,
            in2 => \N__26967\,
            in3 => \N__34381\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__29529\,
            in1 => \N__26961\,
            in2 => \N__26964\,
            in3 => \N__36012\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__38344\,
            in1 => \N__31441\,
            in2 => \_gnd_net_\,
            in3 => \N__34380\,
            lcout => \b2v_inst11.d_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34389\,
            in2 => \N__31581\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_0\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31570\,
            in2 => \N__27234\,
            in3 => \N__27195\,
            lcout => \b2v_inst11.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27192\,
            in2 => \N__31301\,
            in3 => \N__27165\,
            lcout => \b2v_inst11.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_1\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31289\,
            in2 => \N__27162\,
            in3 => \N__27126\,
            lcout => \b2v_inst11.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_2\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29525\,
            in2 => \N__27123\,
            in3 => \N__27093\,
            lcout => \b2v_inst11.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_3\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29514\,
            in2 => \N__36060\,
            in3 => \N__27072\,
            lcout => \b2v_inst11.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_4\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31746\,
            in2 => \N__36061\,
            in3 => \N__27042\,
            lcout => \b2v_inst11.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_5\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35468\,
            in2 => \N__32028\,
            in3 => \N__27018\,
            lcout => \b2v_inst11.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_6\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31969\,
            in2 => \N__31872\,
            in3 => \N__27363\,
            lcout => \b2v_inst11.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37766\,
            in2 => \N__37653\,
            in3 => \N__27342\,
            lcout => \b2v_inst11.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_8\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34600\,
            in2 => \N__27417\,
            in3 => \N__27318\,
            lcout => \b2v_inst11.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_9\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29592\,
            in2 => \N__35210\,
            in3 => \N__27294\,
            lcout => \b2v_inst11.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_10\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29379\,
            in2 => \N__37595\,
            in3 => \N__27291\,
            lcout => \b2v_inst11.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_11\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31794\,
            in2 => \N__34608\,
            in3 => \N__27267\,
            lcout => \b2v_inst11.mult1_un47_sum_1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_12\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35203\,
            in2 => \N__31758\,
            in3 => \N__27264\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3BZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_13\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37588\,
            in2 => \N__29586\,
            in3 => \N__27261\,
            lcout => \b2v_inst11.mult1_un40_sum_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_14\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37589\,
            in2 => \N__29577\,
            in3 => \N__27258\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \b2v_inst11.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.CO2_THRU_LUT4_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27441\,
            lcout => \b2v_inst11.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27437\,
            lcout => \b2v_inst11.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_13_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29538\,
            in3 => \N__34604\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_m_0_6_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__29414\,
            in1 => \N__29507\,
            in2 => \N__29448\,
            in3 => \N__29476\,
            lcout => \b2v_inst11.mult1_un47_sum_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27389\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_9_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__29894\,
            in1 => \N__29796\,
            in2 => \N__33209\,
            in3 => \N__29877\,
            lcout => \b2v_inst6.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36709\,
            ce => \N__33463\,
            sr => \N__33237\
        );

    \b2v_inst6.count_RNI18KF5_8_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__27605\,
            in2 => \_gnd_net_\,
            in3 => \N__33460\,
            lcout => \b2v_inst6.un2_count_1_axb_8\,
            ltout => \b2v_inst6.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_7_c_RNI9E5L1_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__33141\,
            in1 => \N__29793\,
            in2 => \N__27366\,
            in3 => \N__29912\,
            lcout => \b2v_inst6.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI3BLF5_9_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27584\,
            in1 => \N__27596\,
            in2 => \_gnd_net_\,
            in3 => \N__33461\,
            lcout => \b2v_inst6.un2_count_1_axb_9\,
            ltout => \b2v_inst6.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_c_RNIAG6L1_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__33142\,
            in1 => \N__29794\,
            in2 => \N__27609\,
            in3 => \N__29876\,
            lcout => \b2v_inst6.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI18KF5_0_8_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27576\,
            in1 => \N__27606\,
            in2 => \_gnd_net_\,
            in3 => \N__33464\,
            lcout => OPEN,
            ltout => \b2v_inst6.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI4J9VA_9_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__27597\,
            in1 => \N__33462\,
            in2 => \N__27588\,
            in3 => \N__27585\,
            lcout => \b2v_inst6.count_1_i_a3_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_8_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__29795\,
            in1 => \N__33143\,
            in2 => \N__29916\,
            in3 => \N__29930\,
            lcout => \b2v_inst6.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36709\,
            ce => \N__33463\,
            sr => \N__33237\
        );

    \b2v_inst6.curr_state_0_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__29813\,
            in1 => \N__27875\,
            in2 => \N__27468\,
            in3 => \N__27626\,
            lcout => \b2v_inst6.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36835\,
            ce => \N__27546\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_0_0_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33551\,
            lcout => \b2v_inst6.N_394\,
            ltout => \b2v_inst6.N_394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__27465\,
            in1 => \_gnd_net_\,
            in2 => \N__27483\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst6.m6_i_a3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIS68V1_1_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__27480\,
            in1 => \N__33611\,
            in2 => \N__27471\,
            in3 => \N__28382\,
            lcout => \b2v_inst6.curr_stateZ0Z_1\,
            ltout => \b2v_inst6.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__27627\,
            in1 => \N__29779\,
            in2 => \N__27444\,
            in3 => \N__27876\,
            lcout => OPEN,
            ltout => \b2v_inst6.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIR58V1_0_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27801\,
            in2 => \N__27795\,
            in3 => \N__28383\,
            lcout => \b2v_inst6.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNICV5H1_0_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__33552\,
            in1 => \N__33529\,
            in2 => \_gnd_net_\,
            in3 => \N__33101\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_RNICV5H1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNISGKB5_0_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33510\,
            in2 => \N__27792\,
            in3 => \N__33459\,
            lcout => \b2v_inst6.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIAQ3L3_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__27625\,
            in1 => \N__27899\,
            in2 => \N__27888\,
            in3 => \N__35832\,
            lcout => OPEN,
            ltout => \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU4NE4_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27789\,
            in3 => \N__29112\,
            lcout => \N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI_0_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27640\,
            lcout => \b2v_inst6.N_2992_i\,
            ltout => \b2v_inst6.N_2992_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIKIRD1_0_0_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27841\,
            in2 => \N__27738\,
            in3 => \N__27858\,
            lcout => \b2v_inst6.N_276_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst31.un6_output_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27730\,
            in1 => \N__27705\,
            in2 => \N__29118\,
            in3 => \N__27693\,
            lcout => vccinaux_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIKIRD1_0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__27641\,
            in1 => \N__27842\,
            in2 => \_gnd_net_\,
            in3 => \N__27859\,
            lcout => \b2v_inst6.curr_state_RNIKIRD1Z0Z_0\,
            ltout => \b2v_inst6.curr_state_RNIKIRD1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__27887\,
            in1 => \N__27900\,
            in2 => \N__27891\,
            in3 => \N__35833\,
            lcout => \b2v_inst6.delayed_vccin_vccinaux_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNICV5H1_0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27874\,
            in1 => \N__27860\,
            in2 => \N__28410\,
            in3 => \N__27843\,
            lcout => \b2v_inst6.curr_state_RNICV5H1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30083\,
            in2 => \_gnd_net_\,
            in3 => \N__30283\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI1LVK5_0_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27816\,
            in2 => \N__27828\,
            in3 => \N__33803\,
            lcout => \b2v_inst11.count_clkZ0Z_0\,
            ltout => \b2v_inst11.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_1_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30113\,
            in2 => \N__27825\,
            in3 => \N__30284\,
            lcout => \b2v_inst11.count_clk_RNIZ0Z_1\,
            ltout => \b2v_inst11.count_clk_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI2MVK5_1_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27809\,
            in2 => \N__27822\,
            in3 => \N__33802\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_1\,
            ltout => \b2v_inst11.un1_count_clk_2_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_1_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30084\,
            in2 => \N__27819\,
            in3 => \N__30286\,
            lcout => \b2v_inst11.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36840\,
            ce => \N__33808\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_0_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__30285\,
            in1 => \_gnd_net_\,
            in2 => \N__30094\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36840\,
            ce => \N__33808\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI2MVK5_0_1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27810\,
            in1 => \_gnd_net_\,
            in2 => \N__33830\,
            in3 => \N__27966\,
            lcout => \b2v_inst11.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVE6Q5_11_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30174\,
            in1 => \N__30201\,
            in2 => \_gnd_net_\,
            in3 => \N__33807\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI0TCLB_0_2_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__33639\,
            in1 => \N__27918\,
            in2 => \N__32883\,
            in3 => \N__32811\,
            lcout => \b2v_inst11.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI10NQ5_3_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__27909\,
            in1 => \N__30044\,
            in2 => \N__33831\,
            in3 => \N__30253\,
            lcout => \b2v_inst11.count_clkZ0Z_3\,
            ltout => \b2v_inst11.count_clkZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI0TCLB_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__32879\,
            in1 => \N__32810\,
            in2 => \N__27936\,
            in3 => \N__30521\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIG510T_7_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__33638\,
            in1 => \N__27933\,
            in2 => \N__27927\,
            in3 => \N__30150\,
            lcout => \b2v_inst11.count_clk_RNIG510TZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI10NQ5_2_3_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30522\,
            lcout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30252\,
            in2 => \_gnd_net_\,
            in3 => \N__30043\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI10NQ5_0_3_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27908\,
            in2 => \N__27912\,
            in3 => \N__33812\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30045\,
            in2 => \_gnd_net_\,
            in3 => \N__30254\,
            lcout => \b2v_inst11.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36862\,
            ce => \N__33836\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNILIMRT_7_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__39086\,
            in1 => \N__30644\,
            in2 => \N__38416\,
            in3 => \N__28047\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIJ9H9T_5_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39272\,
            in1 => \N__28580\,
            in2 => \N__30768\,
            in3 => \N__29304\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIOM65U_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__38409\,
            in1 => \N__39091\,
            in2 => \N__28041\,
            in3 => \N__38848\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIIGCET1_1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30370\,
            in1 => \N__28028\,
            in2 => \N__28038\,
            in3 => \N__28035\,
            lcout => \b2v_inst11.func_state_RNIIGCET1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30753\,
            lcout => \b2v_inst11.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIAK492_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111111"
        )
    port map (
            in0 => \N__30645\,
            in1 => \N__38408\,
            in2 => \N__39159\,
            in3 => \N__28029\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m2_am_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINCPR4_0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__28705\,
            in1 => \N__28004\,
            in2 => \N__28020\,
            in3 => \N__30754\,
            lcout => \b2v_inst11.func_state_RNINCPR4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8BVM1_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__28005\,
            in1 => \_gnd_net_\,
            in2 => \N__30769\,
            in3 => \N__28593\,
            lcout => \b2v_inst11.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.VCCST_EN_i_0_i_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__28113\,
            in1 => \N__28387\,
            in2 => \N__28815\,
            in3 => \N__38515\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39054\,
            in2 => \_gnd_net_\,
            in3 => \N__30634\,
            lcout => \b2v_inst11.func_state_RNI_0Z0Z_0\,
            ltout => \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28587\,
            in2 => \N__28563\,
            in3 => \N__28157\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_en_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__28560\,
            in1 => \N__35782\,
            in2 => \N__28554\,
            in3 => \N__28608\,
            lcout => \b2v_inst11.count_off_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__38704\,
            in1 => \N__38516\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__28144\,
            in1 => \N__28112\,
            in2 => \N__28413\,
            in3 => \N__28810\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__39273\,
            in1 => \N__38517\,
            in2 => \N__38723\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\,
            ltout => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_0_6_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__28388\,
            in1 => \N__28114\,
            in2 => \N__28161\,
            in3 => \N__28814\,
            lcout => \b2v_inst11.N_382_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIG2BA2_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__28740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37641\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_4_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIOFQO2_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111011"
        )
    port map (
            in0 => \N__28143\,
            in1 => \N__28111\,
            in2 => \N__28050\,
            in3 => \N__28808\,
            lcout => \b2v_inst11.N_140_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_0_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110010001"
        )
    port map (
            in0 => \N__38679\,
            in1 => \N__38553\,
            in2 => \N__30643\,
            in3 => \N__39287\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_7_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__38036\,
            in1 => \N__39127\,
            in2 => \_gnd_net_\,
            in3 => \N__32248\,
            lcout => \b2v_inst11.dutycycle_RNI_9Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_ss0_i_0_x2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__38677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38552\,
            lcout => \b2v_inst11.N_160_i\,
            ltout => \b2v_inst11.N_160_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI5DLR_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28631\,
            in1 => \N__28671\,
            in2 => \N__28722\,
            in3 => \N__30629\,
            lcout => \b2v_inst11.func_state_RNI5DLRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI2MQD_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__38678\,
            in1 => \N__30633\,
            in2 => \N__28679\,
            in3 => \N__28632\,
            lcout => \b2v_inst11.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__34058\,
            in1 => \N__30430\,
            in2 => \N__28680\,
            in3 => \N__28628\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_313_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIL4TIA_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__28934\,
            in1 => \N__35790\,
            in2 => \N__29169\,
            in3 => \N__28599\,
            lcout => \b2v_inst11.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2B_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31320\,
            in1 => \N__30561\,
            in2 => \_gnd_net_\,
            in3 => \N__35919\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIP2BZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNI6TFA1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101011"
        )
    port map (
            in0 => \N__30436\,
            in1 => \N__39117\,
            in2 => \N__28602\,
            in3 => \N__30627\,
            lcout => \b2v_inst11.dutycycle_1_0_1\,
            ltout => \b2v_inst11.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__29162\,
            in1 => \N__35798\,
            in2 => \N__28938\,
            in3 => \N__28935\,
            lcout => \b2v_inst11.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36973\,
            ce => 'H',
            sr => \N__36324\
        );

    \b2v_inst11.dutycycle_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__28923\,
            in1 => \N__29028\,
            in2 => \N__28917\,
            in3 => \N__35792\,
            lcout => \b2v_inst11.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36973\,
            ce => 'H',
            sr => \N__36324\
        );

    \b2v_inst11.func_state_RNIDQ4A1_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__30628\,
            in1 => \N__30437\,
            in2 => \N__31556\,
            in3 => \N__39128\,
            lcout => \b2v_inst11.dutycycle_1_0_0\,
            ltout => \b2v_inst11.dutycycle_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIR0IIA_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__28913\,
            in1 => \N__29027\,
            in2 => \N__28905\,
            in3 => \N__35791\,
            lcout => \b2v_inst11.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_0_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__31527\,
            in1 => \N__35920\,
            in2 => \N__31455\,
            in3 => \N__38274\,
            lcout => \b2v_inst11.dutycycle_RNI_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_1_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__32285\,
            in1 => \N__36174\,
            in2 => \N__28872\,
            in3 => \N__28885\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_RNIDQ4A1_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIQK9K2_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110001"
        )
    port map (
            in0 => \N__34050\,
            in1 => \N__28871\,
            in2 => \N__28830\,
            in3 => \N__28827\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIH3DN3_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__39295\,
            in1 => \_gnd_net_\,
            in2 => \N__28821\,
            in3 => \N__29088\,
            lcout => \b2v_inst11.N_186_i\,
            ltout => \b2v_inst11.N_186_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIH6AK7_2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__37340\,
            in1 => \N__29149\,
            in2 => \N__28818\,
            in3 => \N__29190\,
            lcout => \b2v_inst11.dutycycle_eena_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__31394\,
            in1 => \N__34051\,
            in2 => \N__31557\,
            in3 => \N__38846\,
            lcout => \b2v_inst11.un1_dutycycle_96_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5HTD8_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111111"
        )
    port map (
            in0 => \N__29124\,
            in1 => \N__31393\,
            in2 => \N__29107\,
            in3 => \N__37342\,
            lcout => \b2v_inst11.dutycycle_eena_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNII85R5_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__29150\,
            in1 => \N__29297\,
            in2 => \N__29108\,
            in3 => \N__29130\,
            lcout => \b2v_inst11.N_117_f0_1\,
            ltout => \b2v_inst11.N_117_f0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5HTD8_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__29089\,
            in1 => \N__31528\,
            in2 => \N__29031\,
            in3 => \N__37341\,
            lcout => \b2v_inst11.dutycycle_eena\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_9_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__35361\,
            in1 => \N__35345\,
            in2 => \N__35852\,
            in3 => \N__35325\,
            lcout => \b2v_inst11.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37068\,
            ce => 'H',
            sr => \N__36325\
        );

    \b2v_inst11.dutycycle_2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__29019\,
            in1 => \N__29009\,
            in2 => \N__35856\,
            in3 => \N__28989\,
            lcout => \b2v_inst11.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37068\,
            ce => 'H',
            sr => \N__36325\
        );

    \b2v_inst11.dutycycle_RNITBE6C_2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__29018\,
            in1 => \N__35817\,
            in2 => \N__29010\,
            in3 => \N__28988\,
            lcout => \b2v_inst11.dutycycleZ0Z_1\,
            ltout => \b2v_inst11.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__34165\,
            in1 => \N__28980\,
            in2 => \N__28968\,
            in3 => \N__28965\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__32268\,
            in1 => \_gnd_net_\,
            in2 => \N__39160\,
            in3 => \N__31257\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_2_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__31258\,
            in1 => \N__39095\,
            in2 => \_gnd_net_\,
            in3 => \N__32267\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__32269\,
            in1 => \_gnd_net_\,
            in2 => \N__39161\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.func_state_RNI_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICO933_12_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011111"
        )
    port map (
            in0 => \N__37344\,
            in1 => \N__37704\,
            in2 => \N__29247\,
            in3 => \N__29199\,
            lcout => \b2v_inst11.dutycycle_eena_9\,
            ltout => \b2v_inst11.dutycycle_eena_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNII1EI5_12_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__35779\,
            in1 => \N__31088\,
            in2 => \N__29286\,
            in3 => \N__29363\,
            lcout => \b2v_inst11.dutycycleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNICO933_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__29243\,
            in1 => \N__37343\,
            in2 => \N__29280\,
            in3 => \N__29198\,
            lcout => \b2v_inst11.dutycycle_eena_7\,
            ltout => \b2v_inst11.dutycycle_eena_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_11_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__29355\,
            in1 => \N__31598\,
            in2 => \N__29283\,
            in3 => \N__35781\,
            lcout => \b2v_inst11.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37126\,
            ce => 'H',
            sr => \N__36326\
        );

    \b2v_inst11.dutycycle_RNI_2_12_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__29275\,
            in1 => \N__37705\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5AV24_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__29242\,
            in1 => \N__37500\,
            in2 => \N__29208\,
            in3 => \N__29205\,
            lcout => \b2v_inst11.N_234_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_12_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__29364\,
            in1 => \N__35780\,
            in2 => \N__29373\,
            in3 => \N__31089\,
            lcout => \b2v_inst11.dutycycleZ1Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37126\,
            ce => 'H',
            sr => \N__36326\
        );

    \b2v_inst11.dutycycle_RNIFMPT5_11_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__29354\,
            in1 => \N__31599\,
            in2 => \N__35831\,
            in3 => \N__29346\,
            lcout => \b2v_inst11.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_9_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__38160\,
            in1 => \N__35545\,
            in2 => \N__38351\,
            in3 => \N__34953\,
            lcout => \b2v_inst11.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_8_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__34955\,
            in1 => \N__38336\,
            in2 => \N__37934\,
            in3 => \N__35070\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__29340\,
            in1 => \N__35370\,
            in2 => \N__29334\,
            in3 => \N__31948\,
            lcout => \b2v_inst11.un1_dutycycle_53_55_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__35544\,
            in1 => \_gnd_net_\,
            in2 => \N__34993\,
            in3 => \N__34355\,
            lcout => \b2v_inst11.N_355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_9_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__38161\,
            in1 => \N__34954\,
            in2 => \_gnd_net_\,
            in3 => \N__38329\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_6_a5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_7_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010111"
        )
    port map (
            in0 => \N__38023\,
            in1 => \N__29310\,
            in2 => \N__29313\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__34356\,
            in1 => \N__37923\,
            in2 => \_gnd_net_\,
            in3 => \N__38328\,
            lcout => \b2v_inst11.g0_6_a5_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_15_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__39175\,
            in1 => \N__37593\,
            in2 => \_gnd_net_\,
            in3 => \N__32309\,
            lcout => \b2v_inst11.un1_dutycycle_94_axb_15_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_7_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34982\,
            in1 => \N__38034\,
            in2 => \_gnd_net_\,
            in3 => \N__34382\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_11_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39171\,
            in1 => \N__31970\,
            in2 => \_gnd_net_\,
            in3 => \N__32308\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_7_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010011010"
        )
    port map (
            in0 => \N__37916\,
            in1 => \N__38035\,
            in2 => \N__35010\,
            in3 => \N__34383\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001100"
        )
    port map (
            in0 => \N__34962\,
            in1 => \N__37915\,
            in2 => \N__35554\,
            in3 => \N__38136\,
            lcout => \b2v_inst11.un1_dutycycle_53_44_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_6_i_l_fx_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111111110"
        )
    port map (
            in0 => \N__29442\,
            in1 => \N__29413\,
            in2 => \N__29481\,
            in3 => \N__29508\,
            lcout => \b2v_inst11.mult1_un54_sum_axb_6_i_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_axb_5_i_l_ofx_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29441\,
            in2 => \N__29415\,
            in3 => \N__29477\,
            lcout => \b2v_inst11.mult1_un54_sum_axb_5_i_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_1_axbxc3_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29447\,
            in3 => \N__29409\,
            lcout => \b2v_inst11.mult1_un47_sum1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_11_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011100011000"
        )
    port map (
            in0 => \N__35466\,
            in1 => \N__29601\,
            in2 => \N__31984\,
            in3 => \N__31818\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_15_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29382\,
            in3 => \N__37583\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__38337\,
            in1 => \N__34875\,
            in2 => \N__35490\,
            in3 => \N__29568\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_6\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_11_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__35199\,
            in1 => \N__35467\,
            in2 => \N__29595\,
            in3 => \N__31965\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_15_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__37584\,
            in1 => \_gnd_net_\,
            in2 => \N__29628\,
            in3 => \N__35195\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_14_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35209\,
            in3 => \N__29627\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_11_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111111"
        )
    port map (
            in0 => \N__29567\,
            in1 => \N__35486\,
            in2 => \N__35083\,
            in3 => \N__31961\,
            lcout => \b2v_inst11.un1_dutycycle_53_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_8_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111011"
        )
    port map (
            in0 => \N__35555\,
            in1 => \N__37927\,
            in2 => \N__29616\,
            in3 => \N__38162\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_9_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__38331\,
            in1 => \N__35556\,
            in2 => \N__38169\,
            in3 => \N__35007\,
            lcout => \b2v_inst11.N_35_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_10_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35464\,
            in2 => \_gnd_net_\,
            in3 => \N__34598\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_9_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110100101"
        )
    port map (
            in0 => \N__38167\,
            in1 => \N__29559\,
            in2 => \N__29553\,
            in3 => \N__29550\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_9_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110011"
        )
    port map (
            in0 => \N__35008\,
            in1 => \N__38166\,
            in2 => \N__35085\,
            in3 => \N__38332\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_10_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110101"
        )
    port map (
            in0 => \N__35465\,
            in1 => \N__37928\,
            in2 => \N__29640\,
            in3 => \N__29637\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_11_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__31985\,
            in1 => \N__34599\,
            in2 => \N__29631\,
            in3 => \N__37756\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38330\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35006\,
            lcout => \b2v_inst11.g0_6_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_c_RNI8C4L1_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__29815\,
            in1 => \N__29958\,
            in2 => \N__33230\,
            in3 => \N__29945\,
            lcout => \b2v_inst6.count_rst_7\,
            ltout => \b2v_inst6.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIV4JF5_7_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32447\,
            in2 => \N__29607\,
            in3 => \N__33408\,
            lcout => \b2v_inst6.un2_count_1_axb_7\,
            ltout => \b2v_inst6.un2_count_1_axb_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_7_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__29818\,
            in1 => \N__33198\,
            in2 => \N__29604\,
            in3 => \N__29946\,
            lcout => \b2v_inst6.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36861\,
            ce => \N__33418\,
            sr => \N__33196\
        );

    \b2v_inst6.count_5_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__29655\,
            in1 => \N__29819\,
            in2 => \N__32330\,
            in3 => \N__33195\,
            lcout => \b2v_inst6.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36861\,
            ce => \N__33418\,
            sr => \N__33196\
        );

    \b2v_inst6.un2_count_1_cry_10_c_RNIJOFS1_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__29816\,
            in1 => \N__32404\,
            in2 => \N__33231\,
            in3 => \N__29855\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNILTEO5_11_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29826\,
            in2 => \N__29832\,
            in3 => \N__33409\,
            lcout => \b2v_inst6.countZ0Z_11\,
            ltout => \b2v_inst6.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_11_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__29817\,
            in1 => \N__33197\,
            in2 => \N__29829\,
            in3 => \N__29856\,
            lcout => \b2v_inst6.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36861\,
            ce => \N__33418\,
            sr => \N__33196\
        );

    \b2v_inst6.un2_count_1_cry_4_c_RNI682L1_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__29654\,
            in1 => \N__33188\,
            in2 => \N__32331\,
            in3 => \N__29814\,
            lcout => \b2v_inst6.count_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32429\,
            in2 => \N__33590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_RNIN2P3_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32460\,
            in2 => \_gnd_net_\,
            in3 => \N__29742\,
            lcout => \b2v_inst6.un2_count_1_cry_1_c_RNIN2PZ0Z3\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_1\,
            carryout => \b2v_inst6.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29739\,
            in2 => \_gnd_net_\,
            in3 => \N__29703\,
            lcout => \b2v_inst6.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_2\,
            carryout => \b2v_inst6.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29700\,
            in2 => \_gnd_net_\,
            in3 => \N__29658\,
            lcout => \b2v_inst6.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_3\,
            carryout => \b2v_inst6.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32323\,
            in2 => \_gnd_net_\,
            in3 => \N__29646\,
            lcout => \b2v_inst6.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_4\,
            carryout => \b2v_inst6.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_5_c_RNIRAT3_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32598\,
            in3 => \N__29643\,
            lcout => \b2v_inst6.un2_count_1_cry_5_c_RNIRATZ0Z3\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_5\,
            carryout => \b2v_inst6.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29957\,
            in2 => \_gnd_net_\,
            in3 => \N__29937\,
            lcout => \b2v_inst6.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_6\,
            carryout => \b2v_inst6.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29934\,
            in2 => \_gnd_net_\,
            in3 => \N__29898\,
            lcout => \b2v_inst6.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_7\,
            carryout => \b2v_inst6.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29895\,
            in2 => \_gnd_net_\,
            in3 => \N__29862\,
            lcout => \b2v_inst6.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_9_c_RNIVI14_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32553\,
            in2 => \_gnd_net_\,
            in3 => \N__29859\,
            lcout => \b2v_inst6.un2_count_1_cry_9_c_RNIVIZ0Z14\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_9\,
            carryout => \b2v_inst6.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32408\,
            in2 => \_gnd_net_\,
            in3 => \N__29844\,
            lcout => \b2v_inst6.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_10\,
            carryout => \b2v_inst6.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_11_c_RNI8RAB_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32559\,
            in2 => \_gnd_net_\,
            in3 => \N__29841\,
            lcout => \b2v_inst6.un2_count_1_cry_11_c_RNI8RABZ0\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_11\,
            carryout => \b2v_inst6.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_12_c_RNI9TBB_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30009\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => \b2v_inst6.un2_count_1_cry_12_c_RNI9TBBZ0\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_12\,
            carryout => \b2v_inst6.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_13_c_RNIR6IO5_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32514\,
            in3 => \N__29835\,
            lcout => \b2v_inst6.un2_count_1_cry_13_c_RNIR6IOZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_13\,
            carryout => \b2v_inst6.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_14_c_RNIN0KS1_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__33163\,
            in1 => \_gnd_net_\,
            in2 => \N__32775\,
            in3 => \N__30012\,
            lcout => \b2v_inst6.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIP3HO5_13_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__32734\,
            in1 => \N__33162\,
            in2 => \N__32766\,
            in3 => \N__33410\,
            lcout => \b2v_inst6.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI1I7Q5_0_12_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__30682\,
            in1 => \N__32688\,
            in2 => \N__32709\,
            in3 => \N__30792\,
            lcout => \b2v_inst11.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIM2RL5_0_10_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__30126\,
            in1 => \N__30339\,
            in2 => \N__30801\,
            in3 => \N__30683\,
            lcout => \b2v_inst11.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVE6Q5_0_11_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__30173\,
            in1 => \N__30200\,
            in2 => \N__30687\,
            in3 => \N__30799\,
            lcout => \b2v_inst11.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI3L8Q5_0_13_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__32670\,
            in1 => \N__32651\,
            in2 => \N__30800\,
            in3 => \N__30681\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clkZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIPOH4N_10_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30003\,
            in1 => \N__29997\,
            in2 => \N__29991\,
            in3 => \N__29988\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_o2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIPOH4N_0_10_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33909\,
            in1 => \N__30095\,
            in2 => \N__29982\,
            in3 => \N__30846\,
            lcout => \b2v_inst11.N_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_10_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37087\,
            ce => \N__33797\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIM2RL5_10_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30125\,
            in1 => \N__30337\,
            in2 => \_gnd_net_\,
            in3 => \N__33796\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30117\,
            in2 => \N__30099\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__30289\,
            in1 => \_gnd_net_\,
            in2 => \N__32841\,
            in3 => \N__30060\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_1\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30057\,
            in3 => \N__30030\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_2\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__30287\,
            in1 => \_gnd_net_\,
            in2 => \N__32873\,
            in3 => \N__30027\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_3\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30296\,
            in1 => \N__32973\,
            in2 => \_gnd_net_\,
            in3 => \N__30024\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_4\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__30290\,
            in1 => \_gnd_net_\,
            in2 => \N__33631\,
            in3 => \N__30021\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_5\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__30297\,
            in1 => \_gnd_net_\,
            in2 => \N__32892\,
            in3 => \N__30018\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_6\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30288\,
            in1 => \N__30520\,
            in2 => \_gnd_net_\,
            in3 => \N__30015\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30264\,
            in1 => \N__30470\,
            in2 => \_gnd_net_\,
            in3 => \N__30351\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30279\,
            in1 => \N__30348\,
            in2 => \_gnd_net_\,
            in3 => \N__30324\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30265\,
            in1 => \N__30321\,
            in2 => \_gnd_net_\,
            in3 => \N__30309\,
            lcout => \b2v_inst11.count_clk_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30280\,
            in1 => \N__32715\,
            in2 => \_gnd_net_\,
            in3 => \N__30306\,
            lcout => \b2v_inst11.count_clk_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_11\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30266\,
            in1 => \N__32676\,
            in2 => \_gnd_net_\,
            in3 => \N__30303\,
            lcout => \b2v_inst11.count_clk_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_12\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30281\,
            in1 => \N__30845\,
            in2 => \_gnd_net_\,
            in3 => \N__30300\,
            lcout => \b2v_inst11.count_clk_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_13\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__33905\,
            in1 => \N__30282\,
            in2 => \_gnd_net_\,
            in3 => \N__30204\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_11_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30199\,
            lcout => \b2v_inst11.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37034\,
            ce => \N__33756\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI9CRQ5_0_7_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32924\,
            in1 => \N__33731\,
            in2 => \_gnd_net_\,
            in3 => \N__32909\,
            lcout => \b2v_inst11.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_7_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36967\,
            ce => \N__33835\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIBFSQ5_8_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30486\,
            in1 => \N__33730\,
            in2 => \_gnd_net_\,
            in3 => \N__30497\,
            lcout => \b2v_inst11.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_8_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36967\,
            ce => \N__33835\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIDITQ5_9_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30447\,
            in1 => \N__33732\,
            in2 => \_gnd_net_\,
            in3 => \N__30455\,
            lcout => \b2v_inst11.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_9_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30456\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36967\,
            ce => \N__33835\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_4_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__32147\,
            in1 => \N__39132\,
            in2 => \_gnd_net_\,
            in3 => \N__35027\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_4_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \N__35028\,
            in1 => \_gnd_net_\,
            in2 => \N__39176\,
            in3 => \N__32146\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_2_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30439\,
            in2 => \_gnd_net_\,
            in3 => \N__32163\,
            lcout => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0\,
            ltout => \b2v_inst11.func_state_RNIDQ4A1_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI0O4B5_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__30699\,
            in1 => \N__30782\,
            in2 => \N__30381\,
            in3 => \N__30378\,
            lcout => \b2v_inst11.count_clk_en\,
            ltout => \b2v_inst11.count_clk_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI5O9Q5_14_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30651\,
            in2 => \N__30849\,
            in3 => \N__30662\,
            lcout => \b2v_inst11.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNID7Q51_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000010000"
        )
    port map (
            in0 => \N__30636\,
            in1 => \N__39158\,
            in2 => \N__30828\,
            in3 => \N__30770\,
            lcout => \b2v_inst11.func_state_RNID7Q51Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIJGA54_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__30771\,
            in1 => \N__30705\,
            in2 => \N__39184\,
            in3 => \N__30698\,
            lcout => \b2v_inst11.func_state_RNIJGA54Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37099\,
            ce => \N__33801\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30635\,
            lcout => \b2v_inst11.N_2904_i\,
            ltout => \b2v_inst11.N_2904_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \N__31456\,
            in1 => \_gnd_net_\,
            in2 => \N__30579\,
            in3 => \N__39154\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31558\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_s1_c_RNID26_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30576\,
            in2 => \N__31440\,
            in3 => \N__30552\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_0_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_s1_c_RNIE7GA_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31298\,
            in2 => \N__30549\,
            in3 => \N__30987\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_1_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_s1_c_RNIFCQ4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31110\,
            in2 => \N__34323\,
            in3 => \N__30984\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_2_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_3_s1_c_RNIGH4F_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35025\,
            in2 => \N__30981\,
            in3 => \N__30954\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_3_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_s1_c_RNIHME9_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30951\,
            in2 => \N__32985\,
            in3 => \N__30903\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_4_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_s1_c_RNIIRO3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38227\,
            in2 => \N__31029\,
            in3 => \N__30900\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_5_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_s1_c_RNIJ03E_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38032\,
            in2 => \N__30897\,
            in3 => \N__30882\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_6_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_7_s1_c_RNIK5D8_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37911\,
            in2 => \N__30996\,
            in3 => \N__30879\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_8\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_8_s1_c_RNILAN2_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38158\,
            in2 => \N__30876\,
            in3 => \N__30864\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_9\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_8_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_9_s1_c_RNIMF1D_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30861\,
            in2 => \N__35462\,
            in3 => \N__30852\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_9_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_10_s1_c_RNIU1R8_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31983\,
            in2 => \N__31017\,
            in3 => \N__31074\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_10_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_11_s1_c_RNIV653_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37767\,
            in2 => \N__32055\,
            in3 => \N__31071\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_11_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_12_s1_c_RNI0CFD_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34606\,
            in2 => \N__31068\,
            in3 => \N__31053\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_12_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_13_s1_c_RNI1HP7_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35204\,
            in2 => \N__31050\,
            in3 => \N__31035\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_13_s1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_14_s1_c_RNI2M32_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__39084\,
            in1 => \N__37596\,
            in2 => \N__32278\,
            in3 => \N__31032\,
            lcout => \b2v_inst11.un1_dutycycle_94_s1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_6_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \N__38257\,
            in1 => \_gnd_net_\,
            in2 => \N__32273\,
            in3 => \N__39168\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_11_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39170\,
            in1 => \N__31986\,
            in2 => \_gnd_net_\,
            in3 => \N__32204\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJ9_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31005\,
            in1 => \N__31152\,
            in2 => \_gnd_net_\,
            in3 => \N__36009\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNITMJZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_8_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39169\,
            in1 => \_gnd_net_\,
            in2 => \N__37929\,
            in3 => \N__32203\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_12_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__32199\,
            in1 => \N__37768\,
            in2 => \_gnd_net_\,
            in3 => \N__39167\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_6_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38258\,
            in2 => \N__39185\,
            in3 => \N__32196\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_9_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__32198\,
            in1 => \N__38154\,
            in2 => \_gnd_net_\,
            in3 => \N__39166\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39165\,
            in1 => \_gnd_net_\,
            in2 => \N__34379\,
            in3 => \N__32197\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_7_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__32182\,
            in1 => \_gnd_net_\,
            in2 => \N__38033\,
            in3 => \N__39139\,
            lcout => \b2v_inst11.dutycycle_RNI_10Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_3_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34354\,
            in2 => \N__39178\,
            in3 => \N__32181\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_14_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__32185\,
            in1 => \N__39146\,
            in2 => \_gnd_net_\,
            in3 => \N__35189\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_10_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \N__35434\,
            in1 => \_gnd_net_\,
            in2 => \N__39179\,
            in3 => \N__32183\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EG1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__36211\,
            in1 => \N__36004\,
            in2 => \N__31101\,
            in3 => \N__31638\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIA6EGZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_13_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \N__34563\,
            in1 => \_gnd_net_\,
            in2 => \N__39180\,
            in3 => \N__32184\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNI8SPR1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__36049\,
            in1 => \N__31608\,
            in2 => \N__36230\,
            in3 => \N__31659\,
            lcout => \b2v_inst11.dutycycle_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39177\,
            in3 => \N__32180\,
            lcout => \b2v_inst11.N_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31584\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_s0_c_RNIC05_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31464\,
            in2 => \N__31332\,
            in3 => \N__31305\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_1\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_0_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_s0_c_RNID5FA_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31300\,
            in2 => \N__31194\,
            in3 => \N__31164\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_1_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_s0_c_RNIEAP4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34378\,
            in2 => \N__31161\,
            in3 => \N__31143\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_2_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_3_s0_c_RNIFF3F_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35011\,
            in2 => \N__31140\,
            in3 => \N__31116\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_3_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIGKD9_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34209\,
            in3 => \N__31113\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_4_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIHPN3_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38295\,
            in2 => \N__31734\,
            in3 => \N__31722\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_5_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNIIU1E_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31719\,
            in2 => \N__38022\,
            in3 => \N__31713\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_6_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIJ3C8_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31710\,
            in2 => \N__37875\,
            in3 => \N__31698\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_8\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIK8M2_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31695\,
            in2 => \N__38135\,
            in3 => \N__31686\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_9\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_8_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNILD0D_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31683\,
            in2 => \N__35435\,
            in3 => \N__31674\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_9_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_10_s0_c_RNITVP8_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31671\,
            in2 => \N__31989\,
            in3 => \N__31650\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_10_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_11_s0_c_RNIU443_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31647\,
            in2 => \N__37769\,
            in3 => \N__31629\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_11_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIV9ED_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34567\,
            in2 => \N__31626\,
            in3 => \N__31611\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_12_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI0FO7_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35188\,
            in2 => \N__31857\,
            in3 => \N__31845\,
            lcout => \b2v_inst11.un1_dutycycle_94_s0_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_13_s0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3A64_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__31842\,
            in1 => \N__31830\,
            in2 => \N__36068\,
            in3 => \N__31821\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_14_s0_c_RNI3AZ0Z64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_15_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37540\,
            in2 => \_gnd_net_\,
            in3 => \N__37762\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_6_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__38342\,
            in1 => \N__34874\,
            in2 => \N__31809\,
            in3 => \N__35069\,
            lcout => \b2v_inst11.un1_dutycycle_53_31\,
            ltout => \b2v_inst11.un1_dutycycle_53_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_13_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110000"
        )
    port map (
            in0 => \N__34569\,
            in1 => \N__31779\,
            in2 => \N__31797\,
            in3 => \N__37764\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_13_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35194\,
            in3 => \N__34568\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_14_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_12_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011110000"
        )
    port map (
            in0 => \N__31785\,
            in1 => \N__31778\,
            in2 => \N__31764\,
            in3 => \N__37763\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_14_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__35169\,
            in1 => \_gnd_net_\,
            in2 => \N__31761\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_9_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38309\,
            in1 => \N__38123\,
            in2 => \N__36069\,
            in3 => \N__32040\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_12_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__37765\,
            in1 => \N__39186\,
            in2 => \_gnd_net_\,
            in3 => \N__32306\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100000"
        )
    port map (
            in0 => \N__34368\,
            in1 => \N__38027\,
            in2 => \N__35026\,
            in3 => \N__37871\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_7\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__38340\,
            in1 => \_gnd_net_\,
            in2 => \N__32034\,
            in3 => \N__38131\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_10_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__35463\,
            in1 => \_gnd_net_\,
            in2 => \N__32031\,
            in3 => \N__31883\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIF1_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__36224\,
            in1 => \N__32013\,
            in2 => \N__36059\,
            in3 => \N__32001\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_8_s0_c_RNIMDIFZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_7_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38028\,
            in2 => \_gnd_net_\,
            in3 => \N__38338\,
            lcout => \b2v_inst11.un1_i2_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_7_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000111000"
        )
    port map (
            in0 => \N__37870\,
            in1 => \N__35016\,
            in2 => \N__38037\,
            in3 => \N__34369\,
            lcout => OPEN,
            ltout => \b2v_inst11.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_7_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011100100"
        )
    port map (
            in0 => \N__38130\,
            in1 => \N__38029\,
            in2 => \N__31992\,
            in3 => \N__38339\,
            lcout => \b2v_inst11.un1_N_5\,
            ltout => \b2v_inst11.un1_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_11_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__37872\,
            in1 => \N__31988\,
            in2 => \N__31887\,
            in3 => \N__31884\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRUGF5_0_5_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32340\,
            in1 => \_gnd_net_\,
            in2 => \N__33443\,
            in3 => \N__32349\,
            lcout => OPEN,
            ltout => \b2v_inst6.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIQ34VA_7_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__32454\,
            in1 => \N__32448\,
            in2 => \N__32436\,
            in3 => \N__33379\,
            lcout => \b2v_inst6.count_1_i_a3_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNICV5H1_1_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33186\,
            in1 => \N__32430\,
            in2 => \_gnd_net_\,
            in3 => \N__33588\,
            lcout => \b2v_inst6.count_RNICV5H1Z0Z_1\,
            ltout => \b2v_inst6.count_RNICV5H1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNITHKB5_1_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32384\,
            in2 => \N__32433\,
            in3 => \N__33377\,
            lcout => \b2v_inst6.un2_count_1_axb_1\,
            ltout => \b2v_inst6.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_1_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__33187\,
            in1 => \_gnd_net_\,
            in2 => \N__32418\,
            in3 => \N__33589\,
            lcout => \b2v_inst6.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36968\,
            ce => \N__33417\,
            sr => \N__33240\
        );

    \b2v_inst6.count_RNITHKB5_0_1_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__32415\,
            in1 => \N__33383\,
            in2 => \N__32409\,
            in3 => \N__32385\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIBT0961_1_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32376\,
            in1 => \N__32367\,
            in2 => \N__32358\,
            in3 => \N__32355\,
            lcout => \b2v_inst6.count_1_i_a3_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRUGF5_5_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32348\,
            in1 => \N__32339\,
            in2 => \_gnd_net_\,
            in3 => \N__33378\,
            lcout => \b2v_inst6.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_2_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__33204\,
            in1 => \N__32470\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36899\,
            ce => \N__33385\,
            sr => \N__33222\
        );

    \b2v_inst6.count_RNIH75D5_0_14_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__32535\,
            in1 => \N__32526\,
            in2 => \N__33455\,
            in3 => \N__33223\,
            lcout => \b2v_inst6.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_14_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__32525\,
            in1 => \_gnd_net_\,
            in2 => \N__33235\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36899\,
            ce => \N__33385\,
            sr => \N__33222\
        );

    \b2v_inst6.count_RNIH75D5_14_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__32534\,
            in1 => \N__32524\,
            in2 => \N__33454\,
            in3 => \N__33203\,
            lcout => \b2v_inst6.un2_count_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_RNI32VK1_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__33208\,
            in1 => \N__32474\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI6TISA_2_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010001"
        )
    port map (
            in0 => \N__32484\,
            in1 => \N__32505\,
            in2 => \N__32499\,
            in3 => \N__33386\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIANDN72_2_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32634\,
            in1 => \N__32496\,
            in2 => \N__32487\,
            in3 => \N__32748\,
            lcout => \b2v_inst6.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNILLDF5_2_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__32483\,
            in1 => \N__33202\,
            in2 => \N__32475\,
            in3 => \N__33384\,
            lcout => \b2v_inst6.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIT1IF5_0_6_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__32628\,
            in1 => \N__32619\,
            in2 => \N__33465\,
            in3 => \N__33157\,
            lcout => OPEN,
            ltout => \b2v_inst6.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI9OO0B_10_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__32547\,
            in1 => \N__32781\,
            in2 => \N__32640\,
            in3 => \N__33446\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI0P8PG_12_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__33445\,
            in1 => \N__32589\,
            in2 => \N__32637\,
            in3 => \N__32582\,
            lcout => \b2v_inst6.count_1_i_a3_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_6_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32611\,
            in2 => \_gnd_net_\,
            in3 => \N__33159\,
            lcout => \b2v_inst6.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36830\,
            ce => \N__33444\,
            sr => \N__33160\
        );

    \b2v_inst6.count_RNIT1IF5_6_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__32627\,
            in1 => \N__33155\,
            in2 => \N__32618\,
            in3 => \N__33387\,
            lcout => \b2v_inst6.un2_count_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_11_c_RNIKQGS1_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33161\,
            in2 => \_gnd_net_\,
            in3 => \N__32571\,
            lcout => \b2v_inst6.count_rst_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_12_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32570\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33156\,
            lcout => \b2v_inst6.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36830\,
            ce => \N__33444\,
            sr => \N__33160\
        );

    \b2v_inst6.count_RNIN0GO5_12_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33388\,
            in1 => \N__33158\,
            in2 => \N__32583\,
            in3 => \N__32569\,
            lcout => \b2v_inst6.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNICM6H5_10_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__33341\,
            in1 => \N__32546\,
            in2 => \N__32796\,
            in3 => \N__33217\,
            lcout => \b2v_inst6.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_10_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33218\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32791\,
            lcout => \b2v_inst6.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36890\,
            ce => \N__33457\,
            sr => \N__33216\
        );

    \b2v_inst6.un2_count_1_cry_9_c_RNIBI7L1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33221\,
            lcout => \b2v_inst6.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_13_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__33219\,
            in1 => \_gnd_net_\,
            in2 => \N__32739\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36890\,
            ce => \N__33457\,
            sr => \N__33216\
        );

    \b2v_inst6.count_RNIT9JO5_15_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33458\,
            in1 => \N__33474\,
            in2 => \_gnd_net_\,
            in3 => \N__33488\,
            lcout => \b2v_inst6.countZ0Z_15\,
            ltout => \b2v_inst6.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIP3HO5_0_13_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__32721\,
            in1 => \N__32762\,
            in2 => \N__32751\,
            in3 => \N__33340\,
            lcout => \b2v_inst6.count_1_i_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_12_c_RNILSHS1_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32738\,
            in2 => \_gnd_net_\,
            in3 => \N__33220\,
            lcout => \b2v_inst6.count_rst_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI1I7Q5_12_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__32687\,
            in1 => \N__32701\,
            in2 => \N__33825\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_12_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37067\,
            ce => \N__33822\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI3L8Q5_13_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__32665\,
            in1 => \N__32652\,
            in2 => \N__33826\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_13_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32666\,
            lcout => \b2v_inst11.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37067\,
            ce => \N__33822\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI56PQ5_5_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32966\,
            in2 => \N__33823\,
            in3 => \N__32956\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37067\,
            ce => \N__33822\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI56PQ5_0_5_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32967\,
            in2 => \N__33824\,
            in3 => \N__32957\,
            lcout => \b2v_inst11.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI9CRQ5_7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32928\,
            in1 => \N__33786\,
            in2 => \_gnd_net_\,
            in3 => \N__32903\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI33OQ5_4_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32847\,
            in1 => \_gnd_net_\,
            in2 => \N__33810\,
            in3 => \N__32855\,
            lcout => \b2v_inst11.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_4_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37006\,
            ce => \N__33767\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVSLQ5_2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__32831\,
            in1 => \N__32823\,
            in2 => \N__33809\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_count_clk_2_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_2_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32822\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37006\,
            ce => \N__33767\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVSLQ5_0_2_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__32832\,
            in1 => \N__32821\,
            in2 => \N__33811\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI7RAQ5_15_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33894\,
            in1 => \N__33885\,
            in2 => \_gnd_net_\,
            in3 => \N__33768\,
            lcout => \b2v_inst11.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_15_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33893\,
            lcout => \b2v_inst11.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37006\,
            ce => \N__33767\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI79QQ5_6_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33869\,
            in1 => \N__33855\,
            in2 => \_gnd_net_\,
            in3 => \N__33763\,
            lcout => \b2v_inst11.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIK0DK3_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__33239\,
            in1 => \N__33612\,
            in2 => \_gnd_net_\,
            in3 => \N__35864\,
            lcout => \b2v_inst6.count_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33591\,
            lcout => \b2v_inst6.N_2994_i\,
            ltout => \b2v_inst6.N_2994_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33229\,
            in2 => \N__33534\,
            in3 => \N__33531\,
            lcout => \b2v_inst6.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37100\,
            ce => \N__33407\,
            sr => \N__33238\
        );

    \b2v_inst6.count_15_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33492\,
            lcout => \b2v_inst6.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37100\,
            ce => \N__33407\,
            sr => \N__33238\
        );

    \b2v_inst11.func_state_RNI_4_1_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.func_state_RNI_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_5_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34025\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_5_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_7_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34166\,
            lcout => \b2v_inst11.N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITSFK3_6_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001001110"
        )
    port map (
            in0 => \N__38228\,
            in1 => \N__37178\,
            in2 => \N__34837\,
            in3 => \N__34065\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_231_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIJS2L6_6_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__34131\,
            in1 => \N__34119\,
            in2 => \N__34110\,
            in3 => \N__37278\,
            lcout => \b2v_inst11.dutycycle_eena_13\,
            ltout => \b2v_inst11.dutycycle_eena_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_6_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__34098\,
            in1 => \N__34104\,
            in2 => \N__34107\,
            in3 => \N__35859\,
            lcout => \b2v_inst11.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37085\,
            ce => 'H',
            sr => \N__36362\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVB4_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110111"
        )
    port map (
            in0 => \N__33941\,
            in1 => \N__37277\,
            in2 => \N__34048\,
            in3 => \N__35244\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4\,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNI3QVBZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5IIRB_6_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__34097\,
            in1 => \N__35857\,
            in2 => \N__34089\,
            in3 => \N__34086\,
            lcout => \b2v_inst11.dutycycleZ1Z_6\,
            ltout => \b2v_inst11.dutycycleZ1Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNILF063_6_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110100"
        )
    port map (
            in0 => \N__34030\,
            in1 => \N__34080\,
            in2 => \N__34068\,
            in3 => \N__37617\,
            lcout => \b2v_inst11.dutycycle_RNILF063Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNI1GBN4_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011111"
        )
    port map (
            in0 => \N__34031\,
            in1 => \N__33942\,
            in2 => \N__37316\,
            in3 => \N__35271\,
            lcout => \b2v_inst11.dutycycle_set_1\,
            ltout => \b2v_inst11.dutycycle_set_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_5_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35858\,
            in1 => \N__34451\,
            in2 => \N__34479\,
            in3 => \N__34476\,
            lcout => \b2v_inst11.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37085\,
            ce => 'H',
            sr => \N__36362\
        );

    \b2v_inst11.dutycycle_RNIOFQO2_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__37507\,
            in1 => \N__34322\,
            in2 => \N__37179\,
            in3 => \N__37426\,
            lcout => \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3\,
            ltout => \b2v_inst11.dutycycle_RNIOFQO2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__34412\,
            in1 => \N__34422\,
            in2 => \N__34437\,
            in3 => \N__37283\,
            lcout => \b2v_inst11.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37070\,
            ce => 'H',
            sr => \N__36368\
        );

    \b2v_inst11.dutycycle_RNIM98E2_3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__35835\,
            in1 => \N__34434\,
            in2 => \N__34416\,
            in3 => \N__36220\,
            lcout => \b2v_inst11.dutycycle_RNIM98E2Z0Z_3\,
            ltout => \b2v_inst11.dutycycle_RNIM98E2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI51C57_3_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__34411\,
            in1 => \N__37282\,
            in2 => \N__34398\,
            in3 => \N__34395\,
            lcout => \b2v_inst11.dutycycleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__39280\,
            in1 => \N__34266\,
            in2 => \N__38391\,
            in3 => \N__34819\,
            lcout => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\,
            ltout => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIOMFH6_13_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000000"
        )
    port map (
            in0 => \N__37427\,
            in1 => \N__34497\,
            in2 => \N__34212\,
            in3 => \N__35834\,
            lcout => \b2v_inst11.dutycycle_en_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDQ4A1_4_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36215\,
            in1 => \N__38813\,
            in2 => \_gnd_net_\,
            in3 => \N__37431\,
            lcout => \b2v_inst11.un1_clk_100khz_32_and_i_0_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_8_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__37433\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37876\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_32_and_i_0_c_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI484S5_8_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__34509\,
            in1 => \N__37290\,
            in2 => \N__34512\,
            in3 => \N__37502\,
            lcout => \b2v_inst11.dutycycle_eena_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_10_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__37432\,
            in1 => \_gnd_net_\,
            in2 => \N__35461\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_33_and_i_0_c_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI484S5_10_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__34508\,
            in1 => \N__37289\,
            in2 => \N__34500\,
            in3 => \N__37501\,
            lcout => \b2v_inst11.dutycycle_eena_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5AV24_13_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__38814\,
            in1 => \N__34607\,
            in2 => \N__37512\,
            in3 => \N__36216\,
            lcout => \b2v_inst11.N_153_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5AV24_14_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__35205\,
            in1 => \N__37506\,
            in2 => \N__36231\,
            in3 => \N__38815\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_155_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIOMFH6_14_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__37434\,
            in1 => \N__35788\,
            in2 => \N__34491\,
            in3 => \N__37291\,
            lcout => \b2v_inst11.dutycycle_en_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIG6AA9_7_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__34485\,
            in1 => \N__35845\,
            in2 => \N__37323\,
            in3 => \N__34716\,
            lcout => \b2v_inst11.g0_0_1_0\,
            ltout => \b2v_inst11.g0_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_7_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__34686\,
            in1 => \N__34674\,
            in2 => \N__34488\,
            in3 => \N__36210\,
            lcout => \b2v_inst11.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37144\,
            ce => 'H',
            sr => \N__36348\
        );

    \b2v_inst11.dutycycle_RNI5AV24_7_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__36209\,
            in1 => \N__37981\,
            in2 => \_gnd_net_\,
            in3 => \N__37509\,
            lcout => \b2v_inst11.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIG2BA2_0_0_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__35530\,
            in1 => \N__34854\,
            in2 => \N__38742\,
            in3 => \N__38812\,
            lcout => \b2v_inst11.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_7_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37980\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_7\,
            ltout => \b2v_inst11.dutycycle_RNI_7Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIOFQO2_7_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__37428\,
            in1 => \N__34838\,
            in2 => \N__34725\,
            in3 => \N__34722\,
            lcout => \b2v_inst11.un1_clk_100khz_36_and_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_s0_c_RNI5V4S_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34710\,
            in1 => \N__34698\,
            in2 => \_gnd_net_\,
            in3 => \N__36050\,
            lcout => \b2v_inst11.un1_dutycycle_94_0_7\,
            ltout => \b2v_inst11.un1_dutycycle_94_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIUDOLB_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__34680\,
            in1 => \N__34673\,
            in2 => \N__34665\,
            in3 => \N__36208\,
            lcout => \b2v_inst11.dutycycleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_13_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__34641\,
            in1 => \N__34622\,
            in2 => \N__34635\,
            in3 => \N__36207\,
            lcout => \b2v_inst11.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37086\,
            ce => 'H',
            sr => \N__36361\
        );

    \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQ_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36005\,
            in1 => \N__34662\,
            in2 => \_gnd_net_\,
            in3 => \N__34650\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0\,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_12_s0_c_RNIVLTQZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDSSV8_13_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__34631\,
            in1 => \N__34623\,
            in2 => \N__34611\,
            in3 => \N__36204\,
            lcout => \b2v_inst11.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_s0_c_RNIE51T1_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__36203\,
            in1 => \N__36057\,
            in2 => \N__35289\,
            in3 => \N__35280\,
            lcout => \b2v_inst11.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_s0_c_RNIGFLH1_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__36058\,
            in1 => \N__35262\,
            in2 => \N__36221\,
            in3 => \N__35250\,
            lcout => \b2v_inst11.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IF_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35232\,
            in1 => \_gnd_net_\,
            in2 => \N__36042\,
            in3 => \N__35223\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0\,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_13_s0_c_RNI10IFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIG7HK8_14_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35109\,
            in1 => \N__35093\,
            in2 => \N__35214\,
            in3 => \N__36205\,
            lcout => \b2v_inst11.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_14_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__36206\,
            in1 => \N__35115\,
            in2 => \N__35097\,
            in3 => \N__35108\,
            lcout => \b2v_inst11.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37086\,
            ce => 'H',
            sr => \N__36361\
        );

    \b2v_inst11.dutycycle_RNI_2_10_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35422\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_10\,
            ltout => \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_4_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35031\,
            in3 => \N__35015\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_44_0_3_tz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_8_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__35537\,
            in1 => \N__38108\,
            in2 => \N__34878\,
            in3 => \N__37881\,
            lcout => \b2v_inst11.un1_dutycycle_53_44_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_10_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__35589\,
            in1 => \N__35571\,
            in2 => \N__35583\,
            in3 => \N__35837\,
            lcout => \b2v_inst11.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37142\,
            ce => 'H',
            sr => \N__36366\
        );

    \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNION642_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__36229\,
            in2 => \N__36041\,
            in3 => \N__35595\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642\,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_9_s0_c_RNIONZ0Z642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIM01V8_10_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35579\,
            in1 => \N__35570\,
            in2 => \N__35559\,
            in3 => \N__35836\,
            lcout => \b2v_inst11.dutycycleZ0Z_3\,
            ltout => \b2v_inst11.dutycycleZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__35536\,
            in1 => \N__38106\,
            in2 => \N__35493\,
            in3 => \N__37877\,
            lcout => \b2v_inst11.un1_dutycycle_53_44_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_10_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111111111"
        )
    port map (
            in0 => \N__38107\,
            in1 => \_gnd_net_\,
            in2 => \N__37910\,
            in3 => \N__35423\,
            lcout => \b2v_inst11.g1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI484S5_9_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__37293\,
            in1 => \N__37511\,
            in2 => \N__35298\,
            in3 => \N__37168\,
            lcout => \b2v_inst11.dutycycle_eena_2\,
            ltout => \b2v_inst11.dutycycle_eena_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICK668_9_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__35349\,
            in1 => \N__35830\,
            in2 => \N__35328\,
            in3 => \N__35318\,
            lcout => \b2v_inst11.dutycycleZ0Z_0\,
            ltout => \b2v_inst11.dutycycleZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIDQ4A1_9_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__38802\,
            in1 => \N__36225\,
            in2 => \N__35301\,
            in3 => \N__37429\,
            lcout => \b2v_inst11.un1_clk_100khz_30_and_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIJI598_15_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__36228\,
            in1 => \N__37203\,
            in2 => \N__37191\,
            in3 => \N__37209\,
            lcout => \b2v_inst11.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5AV24_15_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__38803\,
            in1 => \N__36227\,
            in2 => \N__37582\,
            in3 => \N__37510\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_158_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIOMFH6_15_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__37430\,
            in1 => \N__35829\,
            in2 => \N__37365\,
            in3 => \N__37292\,
            lcout => \b2v_inst11.dutycycle_en_12\,
            ltout => \b2v_inst11.dutycycle_en_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_15_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__37202\,
            in1 => \N__37190\,
            in2 => \N__37194\,
            in3 => \N__36226\,
            lcout => \b2v_inst11.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37127\,
            ce => 'H',
            sr => \N__36369\
        );

    \b2v_inst11.func_state_RNIDQ4A1_3_1_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36222\,
            in2 => \_gnd_net_\,
            in3 => \N__38801\,
            lcout => \b2v_inst11.N_326_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_8_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__35889\,
            in1 => \N__35880\,
            in2 => \N__35865\,
            in3 => \N__35895\,
            lcout => \b2v_inst11.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37149\,
            ce => 'H',
            sr => \N__36367\
        );

    \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQ1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__36246\,
            in1 => \N__36223\,
            in2 => \N__36078\,
            in3 => \N__36037\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1\,
            ltout => \b2v_inst11.un1_dutycycle_94_cry_7_s0_c_RNIK3UQZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI99IH8_8_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35888\,
            in1 => \N__35879\,
            in2 => \N__35868\,
            in3 => \N__35860\,
            lcout => \b2v_inst11.dutycycleZ0Z_4\,
            ltout => \b2v_inst11.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_7_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35610\,
            in3 => \N__38030\,
            lcout => \b2v_inst11.un1_i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_12_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37873\,
            in1 => \N__38121\,
            in2 => \N__38341\,
            in3 => \N__37757\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_7_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38122\,
            in1 => \N__38031\,
            in2 => \N__37770\,
            in3 => \N__37874\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_12_7_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__37791\,
            in1 => \N__37785\,
            in2 => \N__37779\,
            in3 => \N__37776\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_s_9_sf_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_12_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__37761\,
            in1 => \_gnd_net_\,
            in2 => \N__37656\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_0_1_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__37602\,
            in1 => \N__38587\,
            in2 => \N__38849\,
            in3 => \N__39182\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_clk_100khz_42_and_i_a2_5_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39283\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38526\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_1_1_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__38590\,
            in1 => \N__39183\,
            in2 => \N__37623\,
            in3 => \N__38832\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDUQ02_1_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__38588\,
            in1 => \_gnd_net_\,
            in2 => \N__37620\,
            in3 => \N__38523\,
            lcout => \b2v_inst11.func_state_RNIDUQ02Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.g2_0_0_0_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__38524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39281\,
            lcout => \b2v_inst11.g2_0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.g2_3_0_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38525\,
            lcout => OPEN,
            ltout => \b2v_inst11.g2_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8H551_1_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__38591\,
            in1 => \N__39181\,
            in2 => \N__38862\,
            in3 => \N__38831\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__38589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38527\,
            lcout => \b2v_inst11.N_161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
